magic
tech sky130A
magscale 1 2
timestamp 1711752077
<< viali >>
rect 10425 18785 10459 18819
rect 11069 18785 11103 18819
rect 12357 18785 12391 18819
rect 13001 18785 13035 18819
rect 16221 18785 16255 18819
rect 18153 18785 18187 18819
rect 18797 18785 18831 18819
rect 19441 18785 19475 18819
rect 20085 18785 20119 18819
rect 20729 18785 20763 18819
rect 21373 18785 21407 18819
rect 22017 18785 22051 18819
rect 31033 18581 31067 18615
rect 18245 16745 18279 16779
rect 9045 16609 9079 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 11345 16609 11379 16643
rect 18061 16609 18095 16643
rect 21465 16609 21499 16643
rect 11621 16541 11655 16575
rect 9137 16405 9171 16439
rect 9781 16405 9815 16439
rect 13093 16405 13127 16439
rect 21557 16405 21591 16439
rect 10425 16201 10459 16235
rect 11345 16201 11379 16235
rect 12541 16201 12575 16235
rect 15393 16201 15427 16235
rect 16129 16201 16163 16235
rect 16570 16201 16604 16235
rect 9873 16065 9907 16099
rect 10149 16065 10183 16099
rect 11069 16065 11103 16099
rect 12909 16065 12943 16099
rect 13369 16065 13403 16099
rect 13921 16065 13955 16099
rect 15761 16065 15795 16099
rect 16313 16065 16347 16099
rect 18705 16065 18739 16099
rect 20637 16065 20671 16099
rect 10241 15997 10275 16031
rect 10425 15997 10459 16031
rect 10977 15997 11011 16031
rect 12633 15997 12667 16031
rect 13001 15997 13035 16031
rect 13645 15997 13679 16031
rect 15853 15997 15887 16031
rect 18337 15997 18371 16031
rect 22753 15997 22787 16031
rect 18245 15929 18279 15963
rect 18981 15929 19015 15963
rect 20913 15929 20947 15963
rect 8401 15861 8435 15895
rect 18061 15861 18095 15895
rect 20453 15861 20487 15895
rect 22385 15861 22419 15895
rect 22845 15861 22879 15895
rect 8401 15657 8435 15691
rect 10701 15657 10735 15691
rect 11437 15657 11471 15691
rect 14749 15657 14783 15691
rect 15761 15657 15795 15691
rect 18245 15657 18279 15691
rect 19165 15657 19199 15691
rect 21373 15657 21407 15691
rect 9673 15589 9707 15623
rect 9873 15589 9907 15623
rect 20453 15589 20487 15623
rect 22109 15589 22143 15623
rect 8677 15521 8711 15555
rect 8953 15521 8987 15555
rect 9137 15521 9171 15555
rect 10517 15521 10551 15555
rect 11345 15521 11379 15555
rect 11621 15521 11655 15555
rect 11713 15521 11747 15555
rect 11897 15521 11931 15555
rect 14657 15521 14691 15555
rect 15669 15521 15703 15555
rect 15853 15521 15887 15555
rect 18337 15521 18371 15555
rect 19073 15521 19107 15555
rect 19901 15521 19935 15555
rect 20637 15521 20671 15555
rect 20821 15521 20855 15555
rect 21005 15521 21039 15555
rect 21281 15521 21315 15555
rect 21465 15521 21499 15555
rect 23673 15521 23707 15555
rect 6653 15453 6687 15487
rect 6929 15453 6963 15487
rect 8493 15453 8527 15487
rect 10333 15453 10367 15487
rect 19993 15453 20027 15487
rect 21833 15453 21867 15487
rect 11621 15385 11655 15419
rect 20269 15385 20303 15419
rect 21005 15385 21039 15419
rect 23857 15385 23891 15419
rect 9505 15317 9539 15351
rect 9689 15317 9723 15351
rect 11897 15317 11931 15351
rect 23581 15317 23615 15351
rect 7941 15113 7975 15147
rect 10425 15113 10459 15147
rect 11161 15113 11195 15147
rect 15301 15113 15335 15147
rect 20637 15113 20671 15147
rect 20913 15113 20947 15147
rect 21097 15113 21131 15147
rect 15485 15045 15519 15079
rect 19993 15045 20027 15079
rect 20085 15045 20119 15079
rect 6193 14977 6227 15011
rect 14933 14977 14967 15011
rect 16129 14977 16163 15011
rect 16681 14977 16715 15011
rect 17141 14977 17175 15011
rect 21649 14977 21683 15011
rect 3801 14909 3835 14943
rect 6285 14909 6319 14943
rect 6469 14909 6503 14943
rect 8033 14909 8067 14943
rect 9137 14909 9171 14943
rect 9321 14909 9355 14943
rect 9965 14909 9999 14943
rect 10977 14909 11011 14943
rect 11345 14909 11379 14943
rect 11437 14909 11471 14943
rect 11621 14909 11655 14943
rect 13737 14909 13771 14943
rect 14841 14909 14875 14943
rect 15025 14909 15059 14943
rect 16773 14909 16807 14943
rect 17417 14909 17451 14943
rect 18521 14909 18555 14943
rect 18705 14909 18739 14943
rect 19257 14909 19291 14943
rect 19717 14909 19751 14943
rect 19809 14909 19843 14943
rect 21189 14909 21223 14943
rect 21373 14909 21407 14943
rect 23857 14909 23891 14943
rect 24124 14909 24158 14943
rect 4077 14841 4111 14875
rect 9505 14841 9539 14875
rect 9873 14841 9907 14875
rect 10149 14841 10183 14875
rect 10241 14841 10275 14875
rect 10793 14841 10827 14875
rect 11897 14841 11931 14875
rect 13645 14841 13679 14875
rect 15117 14841 15151 14875
rect 15761 14841 15795 14875
rect 15853 14841 15887 14875
rect 18981 14841 19015 14875
rect 19993 14841 20027 14875
rect 20361 14841 20395 14875
rect 20729 14841 20763 14875
rect 21281 14841 21315 14875
rect 21925 14841 21959 14875
rect 5549 14773 5583 14807
rect 6653 14773 6687 14807
rect 9597 14773 9631 14807
rect 9781 14773 9815 14807
rect 10441 14773 10475 14807
rect 10609 14773 10643 14807
rect 13369 14773 13403 14807
rect 15317 14773 15351 14807
rect 15577 14773 15611 14807
rect 15945 14773 15979 14807
rect 17325 14773 17359 14807
rect 18429 14773 18463 14807
rect 19441 14773 19475 14807
rect 20269 14773 20303 14807
rect 20453 14773 20487 14807
rect 20939 14773 20973 14807
rect 23397 14773 23431 14807
rect 25237 14773 25271 14807
rect 4905 14569 4939 14603
rect 6193 14569 6227 14603
rect 15025 14569 15059 14603
rect 16681 14569 16715 14603
rect 22661 14569 22695 14603
rect 6561 14501 6595 14535
rect 8484 14501 8518 14535
rect 11590 14501 11624 14535
rect 13522 14501 13556 14535
rect 16313 14501 16347 14535
rect 16405 14501 16439 14535
rect 17693 14501 17727 14535
rect 25114 14501 25148 14535
rect 857 14433 891 14467
rect 2605 14433 2639 14467
rect 2789 14433 2823 14467
rect 3157 14433 3191 14467
rect 3617 14433 3651 14467
rect 4813 14433 4847 14467
rect 6009 14433 6043 14467
rect 6193 14433 6227 14467
rect 6285 14433 6319 14467
rect 10149 14433 10183 14467
rect 15117 14433 15151 14467
rect 15485 14433 15519 14467
rect 16129 14433 16163 14467
rect 16497 14433 16531 14467
rect 17325 14433 17359 14467
rect 22569 14433 22603 14467
rect 23305 14433 23339 14467
rect 23397 14433 23431 14467
rect 23653 14433 23687 14467
rect 24869 14433 24903 14467
rect 3709 14365 3743 14399
rect 3985 14365 4019 14399
rect 8217 14365 8251 14399
rect 11345 14365 11379 14399
rect 13277 14365 13311 14399
rect 15669 14365 15703 14399
rect 15761 14365 15795 14399
rect 17417 14365 17451 14399
rect 19165 14365 19199 14399
rect 2973 14297 3007 14331
rect 1041 14229 1075 14263
rect 8033 14229 8067 14263
rect 9597 14229 9631 14263
rect 9965 14229 9999 14263
rect 12725 14229 12759 14263
rect 14657 14229 14691 14263
rect 15301 14229 15335 14263
rect 17141 14229 17175 14263
rect 23121 14229 23155 14263
rect 24777 14229 24811 14263
rect 26249 14229 26283 14263
rect 3433 14025 3467 14059
rect 7481 14025 7515 14059
rect 2513 13957 2547 13991
rect 4721 13957 4755 13991
rect 6377 13957 6411 13991
rect 14933 13957 14967 13991
rect 23029 13957 23063 13991
rect 3893 13889 3927 13923
rect 6469 13889 6503 13923
rect 13553 13889 13587 13923
rect 15301 13889 15335 13923
rect 16773 13889 16807 13923
rect 21557 13889 21591 13923
rect 21649 13889 21683 13923
rect 2329 13821 2363 13855
rect 2605 13821 2639 13855
rect 2881 13821 2915 13855
rect 3249 13821 3283 13855
rect 3709 13821 3743 13855
rect 4077 13821 4111 13855
rect 4537 13821 4571 13855
rect 4997 13821 5031 13855
rect 6653 13821 6687 13855
rect 6929 13821 6963 13855
rect 7389 13821 7423 13855
rect 9873 13821 9907 13855
rect 10129 13821 10163 13855
rect 13820 13821 13854 13855
rect 15025 13821 15059 13855
rect 18429 13821 18463 13855
rect 18705 13821 18739 13855
rect 21905 13821 21939 13855
rect 24685 13821 24719 13855
rect 24778 13821 24812 13855
rect 25053 13821 25087 13855
rect 25150 13821 25184 13855
rect 3801 13753 3835 13787
rect 4353 13753 4387 13787
rect 4445 13753 4479 13787
rect 5242 13753 5276 13787
rect 18162 13753 18196 13787
rect 18950 13753 18984 13787
rect 21290 13753 21324 13787
rect 24961 13753 24995 13787
rect 2789 13685 2823 13719
rect 3065 13685 3099 13719
rect 3985 13685 4019 13719
rect 4169 13685 4203 13719
rect 6837 13685 6871 13719
rect 11253 13685 11287 13719
rect 17049 13685 17083 13719
rect 20085 13685 20119 13719
rect 20177 13685 20211 13719
rect 25329 13685 25363 13719
rect 2973 13481 3007 13515
rect 3341 13481 3375 13515
rect 10057 13481 10091 13515
rect 14933 13481 14967 13515
rect 3893 13413 3927 13447
rect 7472 13413 7506 13447
rect 10333 13413 10367 13447
rect 12725 13413 12759 13447
rect 15301 13413 15335 13447
rect 20453 13413 20487 13447
rect 26709 13413 26743 13447
rect 2789 13345 2823 13379
rect 3157 13345 3191 13379
rect 3709 13345 3743 13379
rect 4169 13345 4203 13379
rect 4353 13345 4387 13379
rect 8933 13345 8967 13379
rect 10149 13345 10183 13379
rect 10425 13345 10459 13379
rect 10517 13345 10551 13379
rect 11244 13345 11278 13379
rect 12449 13345 12483 13379
rect 12633 13345 12667 13379
rect 12817 13345 12851 13379
rect 13553 13345 13587 13379
rect 13820 13345 13854 13379
rect 15025 13345 15059 13379
rect 15209 13345 15243 13379
rect 15393 13345 15427 13379
rect 16313 13345 16347 13379
rect 16661 13345 16695 13379
rect 18797 13345 18831 13379
rect 18981 13345 19015 13379
rect 19073 13345 19107 13379
rect 19165 13345 19199 13379
rect 20177 13345 20211 13379
rect 20270 13345 20304 13379
rect 20545 13345 20579 13379
rect 20642 13345 20676 13379
rect 22008 13345 22042 13379
rect 23480 13345 23514 13379
rect 24869 13345 24903 13379
rect 25125 13345 25159 13379
rect 26433 13345 26467 13379
rect 26617 13345 26651 13379
rect 26801 13345 26835 13379
rect 7205 13277 7239 13311
rect 8677 13277 8711 13311
rect 10977 13277 11011 13311
rect 16405 13277 16439 13311
rect 21741 13277 21775 13311
rect 23213 13277 23247 13311
rect 4077 13209 4111 13243
rect 16221 13209 16255 13243
rect 17785 13209 17819 13243
rect 26249 13209 26283 13243
rect 3525 13141 3559 13175
rect 4169 13141 4203 13175
rect 5273 13141 5307 13175
rect 5825 13141 5859 13175
rect 6653 13141 6687 13175
rect 8585 13141 8619 13175
rect 10701 13141 10735 13175
rect 12357 13141 12391 13175
rect 13001 13141 13035 13175
rect 13093 13141 13127 13175
rect 15577 13141 15611 13175
rect 19349 13141 19383 13175
rect 20821 13141 20855 13175
rect 23121 13141 23155 13175
rect 24593 13141 24627 13175
rect 26985 13141 27019 13175
rect 4997 12937 5031 12971
rect 8769 12937 8803 12971
rect 14105 12937 14139 12971
rect 15669 12937 15703 12971
rect 18521 12937 18555 12971
rect 21925 12937 21959 12971
rect 23489 12937 23523 12971
rect 24501 12937 24535 12971
rect 24961 12937 24995 12971
rect 7573 12869 7607 12903
rect 12449 12869 12483 12903
rect 15945 12869 15979 12903
rect 21005 12869 21039 12903
rect 23213 12869 23247 12903
rect 3525 12801 3559 12835
rect 5825 12801 5859 12835
rect 16221 12801 16255 12835
rect 3065 12733 3099 12767
rect 3249 12733 3283 12767
rect 5273 12733 5307 12767
rect 5549 12733 5583 12767
rect 5733 12733 5767 12767
rect 6193 12733 6227 12767
rect 6460 12733 6494 12767
rect 7665 12733 7699 12767
rect 8585 12733 8619 12767
rect 9781 12733 9815 12767
rect 11437 12733 11471 12767
rect 11530 12733 11564 12767
rect 11713 12733 11747 12767
rect 11805 12733 11839 12767
rect 11943 12733 11977 12767
rect 12449 12733 12483 12767
rect 12541 12733 12575 12767
rect 12817 12733 12851 12767
rect 13001 12733 13035 12767
rect 13093 12733 13127 12767
rect 13277 12733 13311 12767
rect 14565 12733 14599 12767
rect 14841 12733 14875 12767
rect 15485 12733 15519 12767
rect 16313 12733 16347 12767
rect 17141 12733 17175 12767
rect 19349 12733 19383 12767
rect 19625 12733 19659 12767
rect 21097 12733 21131 12767
rect 21189 12733 21223 12767
rect 21373 12733 21407 12767
rect 21465 12733 21499 12767
rect 21741 12733 21775 12767
rect 22293 12733 22327 12767
rect 22477 12733 22511 12767
rect 23305 12733 23339 12767
rect 23949 12733 23983 12767
rect 24225 12733 24259 12767
rect 24317 12733 24351 12767
rect 24777 12733 24811 12767
rect 26893 12733 26927 12767
rect 27041 12733 27075 12767
rect 27358 12733 27392 12767
rect 12725 12665 12759 12699
rect 12909 12665 12943 12699
rect 13829 12665 13863 12699
rect 16037 12665 16071 12699
rect 16405 12665 16439 12699
rect 16773 12665 16807 12699
rect 17408 12665 17442 12699
rect 19870 12665 19904 12699
rect 21649 12665 21683 12699
rect 24133 12665 24167 12699
rect 27169 12665 27203 12699
rect 27261 12665 27295 12699
rect 5457 12597 5491 12631
rect 5641 12597 5675 12631
rect 9597 12597 9631 12631
rect 12081 12597 12115 12631
rect 13185 12597 13219 12631
rect 14381 12597 14415 12631
rect 14657 12597 14691 12631
rect 16313 12597 16347 12631
rect 19533 12597 19567 12631
rect 22385 12597 22419 12631
rect 27537 12597 27571 12631
rect 3985 12393 4019 12427
rect 4905 12393 4939 12427
rect 5273 12393 5307 12427
rect 7297 12393 7331 12427
rect 11161 12393 11195 12427
rect 12725 12393 12759 12427
rect 13277 12393 13311 12427
rect 13645 12393 13679 12427
rect 16221 12393 16255 12427
rect 17877 12393 17911 12427
rect 19441 12393 19475 12427
rect 23121 12393 23155 12427
rect 25237 12393 25271 12427
rect 26249 12393 26283 12427
rect 27905 12393 27939 12427
rect 3709 12325 3743 12359
rect 5549 12325 5583 12359
rect 7205 12325 7239 12359
rect 7757 12325 7791 12359
rect 9680 12325 9714 12359
rect 12633 12325 12667 12359
rect 13001 12325 13035 12359
rect 14372 12325 14406 12359
rect 18245 12325 18279 12359
rect 18889 12325 18923 12359
rect 22477 12325 22511 12359
rect 25605 12325 25639 12359
rect 25697 12325 25731 12359
rect 26678 12325 26712 12359
rect 3893 12257 3927 12291
rect 4635 12257 4669 12291
rect 4813 12257 4847 12291
rect 4905 12257 4939 12291
rect 4997 12257 5031 12291
rect 5273 12257 5307 12291
rect 5825 12247 5859 12281
rect 6377 12257 6411 12291
rect 6561 12257 6595 12291
rect 6653 12257 6687 12291
rect 6837 12257 6871 12291
rect 6929 12257 6963 12291
rect 7297 12257 7331 12291
rect 7665 12257 7699 12291
rect 7849 12257 7883 12291
rect 7941 12257 7975 12291
rect 8208 12257 8242 12291
rect 9413 12257 9447 12291
rect 10977 12257 11011 12291
rect 11621 12257 11655 12291
rect 11805 12257 11839 12291
rect 12725 12257 12759 12291
rect 12817 12257 12851 12291
rect 13277 12257 13311 12291
rect 13369 12257 13403 12291
rect 13645 12257 13679 12291
rect 13921 12257 13955 12291
rect 15945 12257 15979 12291
rect 16221 12257 16255 12291
rect 16313 12257 16347 12291
rect 16589 12257 16623 12291
rect 16773 12257 16807 12291
rect 16865 12257 16899 12291
rect 17049 12257 17083 12291
rect 17325 12257 17359 12291
rect 17509 12257 17543 12291
rect 18061 12257 18095 12291
rect 18153 12257 18187 12291
rect 18337 12257 18371 12291
rect 18797 12257 18831 12291
rect 19165 12257 19199 12291
rect 19257 12257 19291 12291
rect 19717 12257 19751 12291
rect 19809 12257 19843 12291
rect 20361 12257 20395 12291
rect 20545 12257 20579 12291
rect 20913 12257 20947 12291
rect 21097 12257 21131 12291
rect 21465 12257 21499 12291
rect 21557 12257 21591 12291
rect 21649 12257 21683 12291
rect 22017 12257 22051 12291
rect 22201 12257 22235 12291
rect 22661 12257 22695 12291
rect 22753 12257 22787 12291
rect 23121 12247 23155 12281
rect 23213 12257 23247 12291
rect 23397 12257 23431 12291
rect 23489 12257 23523 12291
rect 23673 12257 23707 12291
rect 24124 12257 24158 12291
rect 25329 12257 25363 12291
rect 25422 12257 25456 12291
rect 25794 12257 25828 12291
rect 26065 12257 26099 12291
rect 26433 12257 26467 12291
rect 29018 12257 29052 12291
rect 5181 12189 5215 12223
rect 6101 12189 6135 12223
rect 6469 12189 6503 12223
rect 6745 12189 6779 12223
rect 7573 12189 7607 12223
rect 12081 12189 12115 12223
rect 13553 12189 13587 12223
rect 14105 12189 14139 12223
rect 16497 12189 16531 12223
rect 16681 12189 16715 12223
rect 17601 12189 17635 12223
rect 18521 12189 18555 12223
rect 19993 12189 20027 12223
rect 21005 12189 21039 12223
rect 21281 12189 21315 12223
rect 21925 12189 21959 12223
rect 22845 12189 22879 12223
rect 23857 12189 23891 12223
rect 29285 12189 29319 12223
rect 4813 12121 4847 12155
rect 5365 12121 5399 12155
rect 5917 12121 5951 12155
rect 7021 12121 7055 12155
rect 7389 12121 7423 12155
rect 13737 12121 13771 12155
rect 15761 12121 15795 12155
rect 17325 12121 17359 12155
rect 18705 12121 18739 12155
rect 18797 12121 18831 12155
rect 19073 12121 19107 12155
rect 19165 12121 19199 12155
rect 20361 12121 20395 12155
rect 21557 12121 21591 12155
rect 21741 12121 21775 12155
rect 22017 12121 22051 12155
rect 22753 12121 22787 12155
rect 23029 12121 23063 12155
rect 3617 12053 3651 12087
rect 6009 12053 6043 12087
rect 7113 12053 7147 12087
rect 9321 12053 9355 12087
rect 10793 12053 10827 12087
rect 15485 12053 15519 12087
rect 17049 12053 17083 12087
rect 19717 12053 19751 12087
rect 20637 12053 20671 12087
rect 21833 12053 21867 12087
rect 23213 12053 23247 12087
rect 23489 12053 23523 12087
rect 25973 12053 26007 12087
rect 27813 12053 27847 12087
rect 7665 11849 7699 11883
rect 8677 11849 8711 11883
rect 11713 11849 11747 11883
rect 18337 11849 18371 11883
rect 19165 11849 19199 11883
rect 19717 11849 19751 11883
rect 21557 11849 21591 11883
rect 23305 11849 23339 11883
rect 24041 11849 24075 11883
rect 27721 11849 27755 11883
rect 7941 11781 7975 11815
rect 17509 11781 17543 11815
rect 17969 11781 18003 11815
rect 19625 11781 19659 11815
rect 22845 11781 22879 11815
rect 23213 11781 23247 11815
rect 3525 11713 3559 11747
rect 3801 11713 3835 11747
rect 8401 11713 8435 11747
rect 9781 11713 9815 11747
rect 13185 11713 13219 11747
rect 17693 11713 17727 11747
rect 23029 11713 23063 11747
rect 23397 11713 23431 11747
rect 3433 11645 3467 11679
rect 4077 11645 4111 11679
rect 4629 11621 4663 11655
rect 4905 11645 4939 11679
rect 6929 11645 6963 11679
rect 7481 11645 7515 11679
rect 7665 11645 7699 11679
rect 7757 11645 7791 11679
rect 7941 11645 7975 11679
rect 8033 11645 8067 11679
rect 8217 11645 8251 11679
rect 8861 11645 8895 11679
rect 9505 11645 9539 11679
rect 9689 11645 9723 11679
rect 11069 11645 11103 11679
rect 11162 11645 11196 11679
rect 11437 11645 11471 11679
rect 11575 11645 11609 11679
rect 11989 11645 12023 11679
rect 12081 11645 12115 11679
rect 12633 11645 12667 11679
rect 12817 11645 12851 11679
rect 12909 11645 12943 11679
rect 13645 11645 13679 11679
rect 13737 11645 13771 11679
rect 13921 11645 13955 11679
rect 15393 11645 15427 11679
rect 15577 11645 15611 11679
rect 15669 11645 15703 11679
rect 17601 11645 17635 11679
rect 17877 11645 17911 11679
rect 17969 11645 18003 11679
rect 18153 11645 18187 11679
rect 18337 11645 18371 11679
rect 18705 11645 18739 11679
rect 19165 11645 19199 11679
rect 19349 11645 19383 11679
rect 19533 11645 19567 11679
rect 19901 11645 19935 11679
rect 22385 11645 22419 11679
rect 22477 11645 22511 11679
rect 22661 11645 22695 11679
rect 22753 11645 22787 11679
rect 23121 11645 23155 11679
rect 23857 11645 23891 11679
rect 25973 11645 26007 11679
rect 26249 11645 26283 11679
rect 26433 11645 26467 11679
rect 26709 11645 26743 11679
rect 27261 11645 27295 11679
rect 27537 11645 27571 11679
rect 5150 11577 5184 11611
rect 8125 11577 8159 11611
rect 11345 11577 11379 11611
rect 11805 11577 11839 11611
rect 12725 11577 12759 11611
rect 17325 11577 17359 11611
rect 19809 11577 19843 11611
rect 20168 11577 20202 11611
rect 3985 11509 4019 11543
rect 4813 11509 4847 11543
rect 6285 11509 6319 11543
rect 6745 11509 6779 11543
rect 9597 11509 9631 11543
rect 12081 11509 12115 11543
rect 14105 11509 14139 11543
rect 15209 11509 15243 11543
rect 17601 11509 17635 11543
rect 21281 11509 21315 11543
rect 22569 11509 22603 11543
rect 22753 11509 22787 11543
rect 26157 11509 26191 11543
rect 2237 11305 2271 11339
rect 4997 11305 5031 11339
rect 7665 11305 7699 11339
rect 8677 11305 8711 11339
rect 9321 11305 9355 11339
rect 11253 11305 11287 11339
rect 11897 11305 11931 11339
rect 13645 11305 13679 11339
rect 16221 11305 16255 11339
rect 18337 11305 18371 11339
rect 20085 11305 20119 11339
rect 20361 11305 20395 11339
rect 22753 11305 22787 11339
rect 23949 11305 23983 11339
rect 25421 11305 25455 11339
rect 26433 11305 26467 11339
rect 3709 11237 3743 11271
rect 8861 11237 8895 11271
rect 9658 11237 9692 11271
rect 13982 11237 14016 11271
rect 15485 11237 15519 11271
rect 16497 11237 16531 11271
rect 18674 11237 18708 11271
rect 22477 11237 22511 11271
rect 24286 11237 24320 11271
rect 25789 11237 25823 11271
rect 25881 11237 25915 11271
rect 27546 11237 27580 11271
rect 5181 11169 5215 11203
rect 6009 11169 6043 11203
rect 7297 11169 7331 11203
rect 7573 11169 7607 11203
rect 7665 11169 7699 11203
rect 8033 11169 8067 11203
rect 8309 11169 8343 11203
rect 8677 11169 8711 11203
rect 8769 11169 8803 11203
rect 8953 11169 8987 11203
rect 9137 11169 9171 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 11805 11169 11839 11203
rect 11989 11169 12023 11203
rect 12541 11169 12575 11203
rect 12725 11169 12759 11203
rect 12817 11169 12851 11203
rect 13001 11169 13035 11203
rect 13461 11169 13495 11203
rect 15209 11169 15243 11203
rect 15393 11169 15427 11203
rect 15577 11169 15611 11203
rect 16221 11169 16255 11203
rect 16589 11169 16623 11203
rect 16681 11169 16715 11203
rect 16957 11169 16991 11203
rect 17141 11169 17175 11203
rect 17233 11169 17267 11203
rect 17417 11169 17451 11203
rect 17877 11169 17911 11203
rect 18153 11169 18187 11203
rect 19901 11169 19935 11203
rect 20269 11169 20303 11203
rect 20453 11169 20487 11203
rect 22109 11169 22143 11203
rect 22201 11169 22235 11203
rect 22661 11169 22695 11203
rect 22753 11169 22787 11203
rect 22845 11169 22879 11203
rect 23121 11169 23155 11203
rect 23305 11169 23339 11203
rect 23765 11169 23799 11203
rect 25513 11169 25547 11203
rect 25606 11169 25640 11203
rect 25978 11169 26012 11203
rect 3985 11101 4019 11135
rect 7389 11101 7423 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 8401 11101 8435 11135
rect 9413 11101 9447 11135
rect 11529 11101 11563 11135
rect 12633 11101 12667 11135
rect 13737 11101 13771 11135
rect 16313 11101 16347 11135
rect 16865 11101 16899 11135
rect 17049 11101 17083 11135
rect 18429 11101 18463 11135
rect 22385 11101 22419 11135
rect 24041 11101 24075 11135
rect 27813 11101 27847 11135
rect 7297 11033 7331 11067
rect 7757 11033 7791 11067
rect 8033 11033 8067 11067
rect 8585 11033 8619 11067
rect 13001 11033 13035 11067
rect 16589 11033 16623 11067
rect 17509 11033 17543 11067
rect 19809 11033 19843 11067
rect 22109 11033 22143 11067
rect 5825 10965 5859 10999
rect 10793 10965 10827 10999
rect 15117 10965 15151 10999
rect 15761 10965 15795 10999
rect 17233 10965 17267 10999
rect 18061 10965 18095 10999
rect 23029 10965 23063 10999
rect 23121 10965 23155 10999
rect 26157 10965 26191 10999
rect 1041 10761 1075 10795
rect 4813 10761 4847 10795
rect 11253 10761 11287 10795
rect 14197 10761 14231 10795
rect 15577 10761 15611 10795
rect 7021 10693 7055 10727
rect 10425 10693 10459 10727
rect 14105 10693 14139 10727
rect 3433 10625 3467 10659
rect 5641 10625 5675 10659
rect 10057 10625 10091 10659
rect 11713 10625 11747 10659
rect 14289 10625 14323 10659
rect 15485 10625 15519 10659
rect 25605 10625 25639 10659
rect 857 10557 891 10591
rect 3689 10557 3723 10591
rect 5181 10557 5215 10591
rect 5908 10557 5942 10591
rect 7757 10533 7791 10567
rect 10241 10557 10275 10591
rect 10701 10557 10735 10591
rect 10977 10557 11011 10591
rect 11069 10557 11103 10591
rect 11437 10557 11471 10591
rect 13553 10557 13587 10591
rect 13921 10557 13955 10591
rect 14197 10557 14231 10591
rect 15577 10557 15611 10591
rect 16221 10557 16255 10591
rect 18705 10557 18739 10591
rect 18961 10557 18995 10591
rect 20729 10557 20763 10591
rect 21557 10557 21591 10591
rect 21741 10557 21775 10591
rect 21925 10557 21959 10591
rect 23406 10557 23440 10591
rect 23673 10557 23707 10591
rect 25145 10557 25179 10591
rect 25329 10557 25363 10591
rect 25697 10557 25731 10591
rect 10885 10489 10919 10523
rect 11958 10489 11992 10523
rect 13737 10489 13771 10523
rect 13829 10489 13863 10523
rect 15853 10489 15887 10523
rect 21649 10489 21683 10523
rect 26341 10489 26375 10523
rect 4997 10421 5031 10455
rect 7941 10421 7975 10455
rect 11621 10421 11655 10455
rect 13093 10421 13127 10455
rect 14565 10421 14599 10455
rect 15209 10421 15243 10455
rect 15761 10421 15795 10455
rect 16405 10421 16439 10455
rect 20085 10421 20119 10455
rect 20913 10421 20947 10455
rect 21373 10421 21407 10455
rect 22293 10421 22327 10455
rect 14381 10217 14415 10251
rect 15209 10217 15243 10251
rect 17601 10217 17635 10251
rect 18061 10217 18095 10251
rect 19441 10217 19475 10251
rect 20361 10217 20395 10251
rect 22661 10217 22695 10251
rect 3249 10149 3283 10183
rect 4528 10149 4562 10183
rect 6460 10149 6494 10183
rect 9689 10149 9723 10183
rect 9781 10149 9815 10183
rect 12449 10149 12483 10183
rect 14105 10149 14139 10183
rect 19650 10149 19684 10183
rect 21526 10149 21560 10183
rect 4261 10081 4295 10115
rect 7665 10081 7699 10115
rect 7932 10081 7966 10115
rect 9413 10081 9447 10115
rect 9506 10081 9540 10115
rect 9878 10081 9912 10115
rect 10149 10081 10183 10115
rect 10333 10081 10367 10115
rect 10425 10081 10459 10115
rect 10517 10081 10551 10115
rect 10977 10081 11011 10115
rect 11069 10081 11103 10115
rect 12081 10081 12115 10115
rect 12633 10081 12667 10115
rect 14933 10081 14967 10115
rect 16221 10081 16255 10115
rect 16477 10081 16511 10115
rect 20729 10081 20763 10115
rect 20913 10081 20947 10115
rect 23121 10081 23155 10115
rect 23388 10081 23422 10115
rect 24685 10081 24719 10115
rect 24869 10081 24903 10115
rect 25421 10081 25455 10115
rect 25605 10081 25639 10115
rect 26617 10081 26651 10115
rect 26884 10081 26918 10115
rect 28345 10081 28379 10115
rect 6193 10013 6227 10047
rect 14841 10013 14875 10047
rect 15025 10013 15059 10047
rect 18153 10013 18187 10047
rect 18245 10013 18279 10047
rect 19165 10013 19199 10047
rect 19533 10013 19567 10047
rect 21281 10013 21315 10047
rect 28089 10013 28123 10047
rect 10057 9945 10091 9979
rect 11345 9945 11379 9979
rect 19809 9945 19843 9979
rect 3157 9877 3191 9911
rect 5641 9877 5675 9911
rect 7573 9877 7607 9911
rect 9045 9877 9079 9911
rect 10701 9877 10735 9911
rect 10977 9877 11011 9911
rect 12725 9877 12759 9911
rect 17693 9877 17727 9911
rect 20729 9877 20763 9911
rect 21097 9877 21131 9911
rect 24501 9877 24535 9911
rect 25881 9877 25915 9911
rect 27997 9877 28031 9911
rect 29469 9877 29503 9911
rect 18061 9673 18095 9707
rect 21465 9673 21499 9707
rect 23305 9673 23339 9707
rect 24869 9673 24903 9707
rect 26157 9673 26191 9707
rect 26341 9673 26375 9707
rect 26801 9673 26835 9707
rect 27261 9673 27295 9707
rect 27629 9673 27663 9707
rect 6469 9605 6503 9639
rect 9321 9605 9355 9639
rect 16221 9605 16255 9639
rect 20545 9605 20579 9639
rect 29009 9605 29043 9639
rect 4905 9537 4939 9571
rect 5917 9537 5951 9571
rect 10793 9537 10827 9571
rect 10977 9537 11011 9571
rect 14013 9537 14047 9571
rect 15761 9537 15795 9571
rect 20386 9537 20420 9571
rect 22293 9537 22327 9571
rect 22569 9537 22603 9571
rect 22753 9537 22787 9571
rect 3249 9469 3283 9503
rect 3505 9469 3539 9503
rect 6101 9469 6135 9503
rect 7113 9469 7147 9503
rect 9229 9469 9263 9503
rect 10057 9469 10091 9503
rect 10701 9469 10735 9503
rect 11069 9469 11103 9503
rect 11621 9469 11655 9503
rect 14197 9469 14231 9503
rect 14565 9469 14599 9503
rect 14657 9469 14691 9503
rect 15393 9469 15427 9503
rect 15485 9469 15519 9503
rect 15853 9469 15887 9503
rect 16681 9469 16715 9503
rect 19901 9469 19935 9503
rect 20269 9469 20303 9503
rect 21649 9469 21683 9503
rect 22017 9469 22051 9503
rect 22109 9469 22143 9503
rect 22385 9469 22419 9503
rect 22477 9469 22511 9503
rect 23121 9469 23155 9503
rect 24501 9469 24535 9503
rect 24593 9469 24627 9503
rect 24869 9469 24903 9503
rect 25973 9469 26007 9503
rect 26065 9469 26099 9503
rect 26985 9469 27019 9503
rect 27077 9469 27111 9503
rect 27261 9469 27295 9503
rect 27445 9469 27479 9503
rect 27905 9469 27939 9503
rect 29193 9469 29227 9503
rect 29285 9469 29319 9503
rect 29561 9469 29595 9503
rect 5089 9401 5123 9435
rect 9597 9401 9631 9435
rect 11888 9401 11922 9435
rect 16948 9401 16982 9435
rect 21743 9401 21777 9435
rect 21833 9401 21867 9435
rect 24685 9401 24719 9435
rect 29377 9401 29411 9435
rect 4629 9333 4663 9367
rect 4997 9333 5031 9367
rect 5457 9333 5491 9367
rect 6009 9333 6043 9367
rect 7297 9333 7331 9367
rect 9873 9333 9907 9367
rect 13001 9333 13035 9367
rect 13645 9333 13679 9367
rect 20177 9333 20211 9367
rect 24317 9333 24351 9367
rect 28089 9333 28123 9367
rect 5641 9129 5675 9163
rect 6929 9129 6963 9163
rect 8677 9129 8711 9163
rect 13921 9129 13955 9163
rect 14933 9129 14967 9163
rect 16497 9129 16531 9163
rect 16681 9129 16715 9163
rect 16957 9129 16991 9163
rect 17509 9129 17543 9163
rect 17693 9129 17727 9163
rect 19349 9129 19383 9163
rect 19901 9129 19935 9163
rect 22661 9129 22695 9163
rect 24041 9129 24075 9163
rect 25513 9129 25547 9163
rect 25973 9129 26007 9163
rect 29929 9129 29963 9163
rect 7542 9061 7576 9095
rect 10425 9061 10459 9095
rect 11069 9061 11103 9095
rect 11437 9061 11471 9095
rect 11897 9061 11931 9095
rect 13093 9061 13127 9095
rect 14197 9061 14231 9095
rect 24378 9061 24412 9095
rect 25605 9061 25639 9095
rect 26893 9061 26927 9095
rect 27261 9061 27295 9095
rect 28702 9061 28736 9095
rect 30297 9061 30331 9095
rect 3249 8993 3283 9027
rect 3617 8993 3651 9027
rect 4528 8993 4562 9027
rect 6745 8993 6779 9027
rect 7297 8993 7331 9027
rect 9597 8993 9631 9027
rect 10057 8993 10091 9027
rect 12265 8993 12299 9027
rect 12541 8993 12575 9027
rect 12817 8993 12851 9027
rect 13001 8993 13035 9027
rect 13231 8993 13265 9027
rect 13553 8993 13587 9027
rect 13737 8993 13771 9027
rect 14565 8993 14599 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 15485 8993 15519 9027
rect 16129 8993 16163 9027
rect 16865 8993 16899 9027
rect 17325 8993 17359 9027
rect 17877 8993 17911 9027
rect 18521 8993 18555 9027
rect 19441 8993 19475 9027
rect 20085 8993 20119 9027
rect 20361 8993 20395 9027
rect 21537 8993 21571 9027
rect 23029 8993 23063 9027
rect 23121 8993 23155 9027
rect 23857 8993 23891 9027
rect 26065 8993 26099 9027
rect 26525 8993 26559 9027
rect 26801 8993 26835 9027
rect 27169 8993 27203 9027
rect 27537 8993 27571 9027
rect 27629 8993 27663 9027
rect 30113 8993 30147 9027
rect 30205 8993 30239 9027
rect 30481 8993 30515 9027
rect 4261 8925 4295 8959
rect 18429 8925 18463 8959
rect 21281 8925 21315 8959
rect 22845 8925 22879 8959
rect 24133 8925 24167 8959
rect 25697 8925 25731 8959
rect 25789 8925 25823 8959
rect 27905 8925 27939 8959
rect 28457 8925 28491 8959
rect 12357 8857 12391 8891
rect 14013 8857 14047 8891
rect 23121 8857 23155 8891
rect 26709 8857 26743 8891
rect 26801 8857 26835 8891
rect 27077 8857 27111 8891
rect 27169 8857 27203 8891
rect 27445 8857 27479 8891
rect 27537 8857 27571 8891
rect 27721 8857 27755 8891
rect 29837 8857 29871 8891
rect 7205 8789 7239 8823
rect 9413 8789 9447 8823
rect 11805 8789 11839 8823
rect 13369 8789 13403 8823
rect 13553 8789 13587 8823
rect 14197 8789 14231 8823
rect 16488 8789 16522 8823
rect 19533 8789 19567 8823
rect 23765 8789 23799 8823
rect 27629 8789 27663 8823
rect 27997 8789 28031 8823
rect 4629 8585 4663 8619
rect 4997 8585 5031 8619
rect 5733 8585 5767 8619
rect 11805 8585 11839 8619
rect 13829 8585 13863 8619
rect 19993 8585 20027 8619
rect 21189 8585 21223 8619
rect 23121 8585 23155 8619
rect 25421 8585 25455 8619
rect 27905 8585 27939 8619
rect 30389 8585 30423 8619
rect 10885 8517 10919 8551
rect 12081 8517 12115 8551
rect 12173 8517 12207 8551
rect 14473 8517 14507 8551
rect 16773 8517 16807 8551
rect 23949 8517 23983 8551
rect 26617 8517 26651 8551
rect 6469 8449 6503 8483
rect 8861 8449 8895 8483
rect 11253 8449 11287 8483
rect 11897 8449 11931 8483
rect 17141 8449 17175 8483
rect 19625 8449 19659 8483
rect 23029 8449 23063 8483
rect 27997 8449 28031 8483
rect 3249 8381 3283 8415
rect 5181 8381 5215 8415
rect 5549 8381 5583 8415
rect 5917 8381 5951 8415
rect 6193 8381 6227 8415
rect 6285 8381 6319 8415
rect 6561 8381 6595 8415
rect 6837 8381 6871 8415
rect 7021 8381 7055 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 7481 8381 7515 8415
rect 9128 8381 9162 8415
rect 10701 8381 10735 8415
rect 10885 8381 10919 8415
rect 10977 8381 11011 8415
rect 11161 8381 11195 8415
rect 11713 8381 11747 8415
rect 11805 8381 11839 8415
rect 12173 8381 12207 8415
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 12725 8381 12759 8415
rect 14013 8381 14047 8415
rect 14105 8381 14139 8415
rect 14289 8381 14323 8415
rect 14473 8381 14507 8415
rect 15853 8381 15887 8415
rect 16313 8381 16347 8415
rect 16497 8381 16531 8415
rect 16589 8381 16623 8415
rect 18890 8375 18924 8409
rect 19073 8381 19107 8415
rect 19257 8381 19291 8415
rect 19349 8381 19383 8415
rect 19809 8381 19843 8415
rect 21005 8381 21039 8415
rect 22569 8381 22603 8415
rect 22753 8381 22787 8415
rect 23121 8381 23155 8415
rect 23397 8381 23431 8415
rect 23489 8381 23523 8415
rect 23857 8381 23891 8415
rect 24225 8381 24259 8415
rect 24409 8381 24443 8415
rect 25605 8381 25639 8415
rect 25697 8381 25731 8415
rect 25881 8381 25915 8415
rect 25973 8381 26007 8415
rect 26433 8381 26467 8415
rect 26617 8381 26651 8415
rect 26709 8381 26743 8415
rect 26893 8381 26927 8415
rect 26985 8381 27019 8415
rect 27353 8381 27387 8415
rect 27721 8381 27755 8415
rect 27905 8381 27939 8415
rect 28273 8381 28307 8415
rect 29009 8381 29043 8415
rect 3494 8313 3528 8347
rect 7389 8313 7423 8347
rect 11069 8313 11103 8347
rect 11529 8313 11563 8347
rect 17408 8313 17442 8347
rect 18981 8313 19015 8347
rect 22661 8313 22695 8347
rect 22845 8313 22879 8347
rect 23213 8313 23247 8347
rect 24133 8313 24167 8347
rect 24317 8313 24351 8347
rect 29254 8313 29288 8347
rect 10241 8245 10275 8279
rect 12357 8245 12391 8279
rect 12541 8245 12575 8279
rect 16313 8245 16347 8279
rect 18521 8245 18555 8279
rect 18705 8245 18739 8279
rect 23489 8245 23523 8279
rect 23857 8245 23891 8279
rect 26801 8245 26835 8279
rect 27169 8245 27203 8279
rect 27537 8245 27571 8279
rect 28457 8245 28491 8279
rect 5273 8041 5307 8075
rect 7297 8041 7331 8075
rect 9045 8041 9079 8075
rect 10149 8041 10183 8075
rect 10609 8041 10643 8075
rect 11161 8041 11195 8075
rect 13369 8041 13403 8075
rect 13461 8041 13495 8075
rect 15393 8041 15427 8075
rect 16957 8041 16991 8075
rect 17693 8041 17727 8075
rect 18705 8041 18739 8075
rect 19073 8041 19107 8075
rect 20269 8041 20303 8075
rect 23029 8041 23063 8075
rect 25697 8041 25731 8075
rect 29561 8041 29595 8075
rect 9781 7973 9815 8007
rect 9873 7973 9907 8007
rect 12256 7973 12290 8007
rect 13737 7973 13771 8007
rect 13829 7973 13863 8007
rect 16865 7973 16899 8007
rect 18613 7973 18647 8007
rect 19349 7973 19383 8007
rect 19809 7973 19843 8007
rect 20361 7973 20395 8007
rect 27353 7973 27387 8007
rect 29837 7973 29871 8007
rect 4813 7905 4847 7939
rect 5181 7905 5215 7939
rect 5365 7905 5399 7939
rect 6009 7905 6043 7939
rect 6469 7905 6503 7939
rect 6745 7905 6779 7939
rect 7113 7905 7147 7939
rect 7205 7905 7239 7939
rect 7921 7905 7955 7939
rect 9597 7905 9631 7939
rect 9965 7905 9999 7939
rect 10229 7911 10263 7945
rect 11161 7905 11195 7939
rect 11529 7905 11563 7939
rect 11621 7905 11655 7939
rect 11805 7905 11839 7939
rect 13640 7905 13674 7939
rect 13957 7905 13991 7939
rect 14105 7905 14139 7939
rect 15025 7905 15059 7939
rect 15209 7905 15243 7939
rect 15485 7905 15519 7939
rect 15669 7905 15703 7939
rect 16313 7905 16347 7939
rect 16405 7905 16439 7939
rect 16497 7905 16531 7939
rect 16681 7905 16715 7939
rect 17509 7905 17543 7939
rect 17877 7905 17911 7939
rect 18822 7905 18856 7939
rect 19257 7905 19291 7939
rect 20478 7905 20512 7939
rect 22405 7905 22439 7939
rect 22937 7905 22971 7939
rect 23121 7905 23155 7939
rect 23397 7905 23431 7939
rect 23765 7905 23799 7939
rect 23949 7905 23983 7939
rect 24041 7905 24075 7939
rect 24225 7905 24259 7939
rect 24317 7905 24351 7939
rect 24573 7905 24607 7939
rect 27261 7905 27295 7939
rect 27623 7905 27657 7939
rect 27721 7905 27755 7939
rect 27997 7905 28031 7939
rect 28089 7905 28123 7939
rect 28345 7905 28379 7939
rect 29745 7905 29779 7939
rect 29929 7905 29963 7939
rect 30113 7905 30147 7939
rect 30757 7905 30791 7939
rect 7665 7837 7699 7871
rect 10333 7837 10367 7871
rect 11437 7837 11471 7871
rect 11989 7837 12023 7871
rect 15853 7837 15887 7871
rect 18337 7837 18371 7871
rect 19993 7837 20027 7871
rect 22661 7837 22695 7871
rect 23673 7837 23707 7871
rect 31033 7837 31067 7871
rect 11253 7769 11287 7803
rect 11529 7769 11563 7803
rect 19809 7769 19843 7803
rect 23213 7769 23247 7803
rect 27537 7769 27571 7803
rect 27905 7769 27939 7803
rect 27997 7769 28031 7803
rect 29469 7769 29503 7803
rect 5641 7701 5675 7735
rect 10425 7701 10459 7735
rect 15209 7701 15243 7735
rect 16129 7701 16163 7735
rect 17417 7701 17451 7735
rect 18981 7701 19015 7735
rect 20637 7701 20671 7735
rect 21281 7701 21315 7735
rect 23765 7701 23799 7735
rect 24225 7701 24259 7735
rect 27077 7701 27111 7735
rect 27445 7701 27479 7735
rect 6653 7497 6687 7531
rect 6929 7497 6963 7531
rect 7481 7497 7515 7531
rect 7757 7497 7791 7531
rect 10425 7497 10459 7531
rect 10517 7497 10551 7531
rect 11805 7497 11839 7531
rect 14197 7497 14231 7531
rect 16221 7497 16255 7531
rect 16497 7497 16531 7531
rect 16957 7497 16991 7531
rect 21925 7497 21959 7531
rect 24409 7497 24443 7531
rect 25605 7497 25639 7531
rect 28089 7497 28123 7531
rect 30389 7497 30423 7531
rect 7849 7429 7883 7463
rect 17509 7429 17543 7463
rect 23305 7429 23339 7463
rect 23397 7429 23431 7463
rect 23857 7429 23891 7463
rect 23949 7429 23983 7463
rect 2789 7361 2823 7395
rect 3065 7361 3099 7395
rect 3525 7361 3559 7395
rect 17049 7361 17083 7395
rect 17877 7361 17911 7395
rect 23581 7361 23615 7395
rect 24133 7361 24167 7395
rect 26341 7361 26375 7395
rect 29009 7361 29043 7395
rect 2697 7293 2731 7327
rect 3249 7293 3283 7327
rect 5089 7293 5123 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 7565 7289 7599 7323
rect 8033 7293 8067 7327
rect 8401 7293 8435 7327
rect 9873 7293 9907 7327
rect 10149 7293 10183 7327
rect 10241 7293 10275 7327
rect 10701 7293 10735 7327
rect 10977 7293 11011 7327
rect 11713 7293 11747 7327
rect 11805 7293 11839 7327
rect 11989 7293 12023 7327
rect 13553 7293 13587 7327
rect 13646 7293 13680 7327
rect 13829 7293 13863 7327
rect 14018 7293 14052 7327
rect 14841 7293 14875 7327
rect 15108 7293 15142 7327
rect 16503 7293 16537 7327
rect 16681 7293 16715 7327
rect 16773 7293 16807 7327
rect 16865 7293 16899 7327
rect 17325 7293 17359 7327
rect 17417 7293 17451 7327
rect 17693 7293 17727 7327
rect 17785 7293 17819 7327
rect 17969 7293 18003 7327
rect 18061 7293 18095 7327
rect 18705 7293 18739 7327
rect 18889 7293 18923 7327
rect 21281 7293 21315 7327
rect 21429 7293 21463 7327
rect 21649 7293 21683 7327
rect 21746 7293 21780 7327
rect 23305 7293 23339 7327
rect 23857 7293 23891 7327
rect 24225 7293 24259 7327
rect 24961 7293 24995 7327
rect 25054 7293 25088 7327
rect 25467 7293 25501 7327
rect 26065 7293 26099 7327
rect 26249 7293 26283 7327
rect 27905 7293 27939 7327
rect 28181 7293 28215 7327
rect 5334 7225 5368 7259
rect 8646 7225 8680 7259
rect 10057 7225 10091 7259
rect 13921 7225 13955 7259
rect 17141 7225 17175 7259
rect 21557 7225 21591 7259
rect 25237 7225 25271 7259
rect 25329 7225 25363 7259
rect 26709 7225 26743 7259
rect 27353 7225 27387 7259
rect 27721 7225 27755 7259
rect 29254 7225 29288 7259
rect 4997 7157 5031 7191
rect 6469 7157 6503 7191
rect 9781 7157 9815 7191
rect 10885 7157 10919 7191
rect 17417 7157 17451 7191
rect 18797 7157 18831 7191
rect 26157 7157 26191 7191
rect 26801 7157 26835 7191
rect 28365 7157 28399 7191
rect 4261 6953 4295 6987
rect 7481 6953 7515 6987
rect 12725 6953 12759 6987
rect 17233 6953 17267 6987
rect 17417 6953 17451 6987
rect 17785 6953 17819 6987
rect 19809 6953 19843 6987
rect 22845 6953 22879 6987
rect 25421 6953 25455 6987
rect 28641 6953 28675 6987
rect 18061 6885 18095 6919
rect 25973 6885 26007 6919
rect 27506 6885 27540 6919
rect 29009 6885 29043 6919
rect 4353 6817 4387 6851
rect 6081 6817 6115 6851
rect 7481 6817 7515 6851
rect 7849 6817 7883 6851
rect 7941 6817 7975 6851
rect 8401 6817 8435 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 8769 6817 8803 6851
rect 8953 6817 8987 6851
rect 11437 6817 11471 6851
rect 11713 6817 11747 6851
rect 12541 6817 12575 6851
rect 12817 6817 12851 6851
rect 13277 6817 13311 6851
rect 13544 6817 13578 6851
rect 15025 6817 15059 6851
rect 17141 6817 17175 6851
rect 17325 6817 17359 6851
rect 17417 6817 17451 6851
rect 17785 6817 17819 6851
rect 17877 6817 17911 6851
rect 18153 6817 18187 6851
rect 18685 6817 18719 6851
rect 20085 6817 20119 6851
rect 20453 6817 20487 6851
rect 20601 6817 20635 6851
rect 20729 6817 20763 6851
rect 20821 6817 20855 6851
rect 20918 6817 20952 6851
rect 21925 6817 21959 6851
rect 22845 6817 22879 6851
rect 23213 6817 23247 6851
rect 23305 6817 23339 6851
rect 23581 6817 23615 6851
rect 23765 6817 23799 6851
rect 24041 6817 24075 6851
rect 24297 6817 24331 6851
rect 25697 6817 25731 6851
rect 25881 6817 25915 6851
rect 26249 6817 26283 6851
rect 26617 6817 26651 6851
rect 26985 6817 27019 6851
rect 27169 6817 27203 6851
rect 28733 6817 28767 6851
rect 28826 6817 28860 6851
rect 29101 6817 29135 6851
rect 29239 6817 29273 6851
rect 5825 6749 5859 6783
rect 7757 6749 7791 6783
rect 8125 6749 8159 6783
rect 8861 6749 8895 6783
rect 11805 6749 11839 6783
rect 12909 6749 12943 6783
rect 13093 6749 13127 6783
rect 17693 6749 17727 6783
rect 18429 6749 18463 6783
rect 21741 6749 21775 6783
rect 22201 6749 22235 6783
rect 22753 6749 22787 6783
rect 23121 6749 23155 6783
rect 23489 6749 23523 6783
rect 26893 6749 26927 6783
rect 27077 6749 27111 6783
rect 27261 6749 27295 6783
rect 7573 6681 7607 6715
rect 7849 6681 7883 6715
rect 8493 6681 8527 6715
rect 12817 6681 12851 6715
rect 14657 6681 14691 6715
rect 17509 6681 17543 6715
rect 18337 6681 18371 6715
rect 21097 6681 21131 6715
rect 22937 6681 22971 6715
rect 23213 6681 23247 6715
rect 23581 6681 23615 6715
rect 26157 6681 26191 6715
rect 26249 6681 26283 6715
rect 26709 6681 26743 6715
rect 29377 6681 29411 6715
rect 7205 6613 7239 6647
rect 11253 6613 11287 6647
rect 11713 6613 11747 6647
rect 12081 6613 12115 6647
rect 14841 6613 14875 6647
rect 15117 6613 15151 6647
rect 20269 6613 20303 6647
rect 25697 6613 25731 6647
rect 26801 6613 26835 6647
rect 12265 6409 12299 6443
rect 13185 6409 13219 6443
rect 13553 6409 13587 6443
rect 14565 6409 14599 6443
rect 16681 6409 16715 6443
rect 21465 6409 21499 6443
rect 23489 6409 23523 6443
rect 24041 6409 24075 6443
rect 24685 6409 24719 6443
rect 26893 6409 26927 6443
rect 27353 6409 27387 6443
rect 15209 6341 15243 6375
rect 18705 6341 18739 6375
rect 19165 6341 19199 6375
rect 26801 6341 26835 6375
rect 5089 6273 5123 6307
rect 8769 6273 8803 6307
rect 20085 6273 20119 6307
rect 3341 6205 3375 6239
rect 5365 6205 5399 6239
rect 5733 6205 5767 6239
rect 6837 6205 6871 6239
rect 8493 6205 8527 6239
rect 10793 6205 10827 6239
rect 11060 6205 11094 6239
rect 12449 6205 12483 6239
rect 12817 6205 12851 6239
rect 13185 6205 13219 6239
rect 13369 6205 13403 6239
rect 13737 6205 13771 6239
rect 14197 6205 14231 6239
rect 14381 6205 14415 6239
rect 14657 6205 14691 6239
rect 14749 6205 14783 6239
rect 15025 6205 15059 6239
rect 15301 6205 15335 6239
rect 18705 6205 18739 6239
rect 18797 6205 18831 6239
rect 18981 6205 19015 6239
rect 19073 6205 19107 6239
rect 20352 6205 20386 6239
rect 22569 6205 22603 6239
rect 22661 6205 22695 6239
rect 22845 6205 22879 6239
rect 22937 6205 22971 6239
rect 23397 6205 23431 6239
rect 23489 6205 23523 6239
rect 23673 6205 23707 6239
rect 23857 6205 23891 6239
rect 24133 6205 24167 6239
rect 24317 6205 24351 6239
rect 24501 6205 24535 6239
rect 25973 6205 26007 6239
rect 26157 6205 26191 6239
rect 26249 6205 26283 6239
rect 26433 6205 26467 6239
rect 26617 6205 26651 6239
rect 27169 6205 27203 6239
rect 3617 6137 3651 6171
rect 5273 6137 5307 6171
rect 6009 6137 6043 6171
rect 7082 6137 7116 6171
rect 9014 6137 9048 6171
rect 12541 6137 12575 6171
rect 12633 6137 12667 6171
rect 14289 6137 14323 6171
rect 14473 6137 14507 6171
rect 15546 6137 15580 6171
rect 19349 6137 19383 6171
rect 24409 6137 24443 6171
rect 26065 6137 26099 6171
rect 26525 6137 26559 6171
rect 5457 6069 5491 6103
rect 5641 6069 5675 6103
rect 5825 6069 5859 6103
rect 8217 6069 8251 6103
rect 8677 6069 8711 6103
rect 10149 6069 10183 6103
rect 12173 6069 12207 6103
rect 19073 6069 19107 6103
rect 22753 6069 22787 6103
rect 23121 6069 23155 6103
rect 3617 5865 3651 5899
rect 6101 5865 6135 5899
rect 10517 5865 10551 5899
rect 12817 5865 12851 5899
rect 18245 5865 18279 5899
rect 20821 5865 20855 5899
rect 23213 5865 23247 5899
rect 24685 5865 24719 5899
rect 26157 5865 26191 5899
rect 27261 5865 27295 5899
rect 28733 5865 28767 5899
rect 10241 5797 10275 5831
rect 13952 5797 13986 5831
rect 25022 5797 25056 5831
rect 27598 5797 27632 5831
rect 3525 5729 3559 5763
rect 3709 5729 3743 5763
rect 5825 5729 5859 5763
rect 6193 5729 6227 5763
rect 9965 5729 9999 5763
rect 10149 5729 10183 5763
rect 10333 5729 10367 5763
rect 14749 5729 14783 5763
rect 15117 5729 15151 5763
rect 16313 5729 16347 5763
rect 16865 5729 16899 5763
rect 17121 5729 17155 5763
rect 19697 5729 19731 5763
rect 22089 5729 22123 5763
rect 23305 5729 23339 5763
rect 23572 5729 23606 5763
rect 24777 5729 24811 5763
rect 27077 5729 27111 5763
rect 27353 5729 27387 5763
rect 6009 5661 6043 5695
rect 14197 5661 14231 5695
rect 14473 5661 14507 5695
rect 19441 5661 19475 5695
rect 21833 5661 21867 5695
rect 5825 5593 5859 5627
rect 14565 5525 14599 5559
rect 14933 5525 14967 5559
rect 15209 5525 15243 5559
rect 16221 5525 16255 5559
rect 9965 5321 9999 5355
rect 11437 5321 11471 5355
rect 13185 5321 13219 5355
rect 16497 5321 16531 5355
rect 20085 5321 20119 5355
rect 21741 5321 21775 5355
rect 27721 5321 27755 5355
rect 27077 5253 27111 5287
rect 27353 5253 27387 5287
rect 3341 5185 3375 5219
rect 5089 5185 5123 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 11805 5185 11839 5219
rect 14657 5185 14691 5219
rect 15025 5185 15059 5219
rect 5549 5117 5583 5151
rect 5825 5117 5859 5151
rect 5917 5117 5951 5151
rect 6101 5117 6135 5151
rect 6469 5117 6503 5151
rect 7205 5117 7239 5151
rect 7941 5117 7975 5151
rect 8585 5117 8619 5151
rect 8841 5117 8875 5151
rect 10057 5117 10091 5151
rect 14749 5117 14783 5151
rect 17969 5117 18003 5151
rect 18705 5117 18739 5151
rect 20361 5117 20395 5151
rect 20617 5117 20651 5151
rect 26617 5117 26651 5151
rect 26893 5117 26927 5151
rect 27169 5117 27203 5151
rect 27629 5117 27663 5151
rect 27905 5117 27939 5151
rect 3617 5049 3651 5083
rect 10302 5049 10336 5083
rect 12072 5049 12106 5083
rect 14381 5049 14415 5083
rect 18950 5049 18984 5083
rect 5365 4981 5399 5015
rect 5733 4981 5767 5015
rect 5917 4981 5951 5015
rect 7021 4981 7055 5015
rect 8033 4981 8067 5015
rect 14105 4981 14139 5015
rect 14289 4981 14323 5015
rect 14473 4981 14507 5015
rect 17877 4981 17911 5015
rect 26801 4981 26835 5015
rect 27445 4981 27479 5015
rect 4445 4777 4479 4811
rect 10241 4777 10275 4811
rect 10425 4777 10459 4811
rect 13553 4777 13587 4811
rect 14121 4777 14155 4811
rect 14381 4777 14415 4811
rect 14657 4777 14691 4811
rect 18429 4777 18463 4811
rect 20361 4777 20395 4811
rect 24869 4777 24903 4811
rect 5181 4709 5215 4743
rect 7205 4709 7239 4743
rect 8953 4709 8987 4743
rect 13921 4709 13955 4743
rect 14933 4709 14967 4743
rect 16957 4709 16991 4743
rect 20637 4709 20671 4743
rect 20853 4709 20887 4743
rect 21557 4709 21591 4743
rect 21649 4709 21683 4743
rect 23734 4709 23768 4743
rect 4353 4641 4387 4675
rect 5365 4641 5399 4675
rect 5549 4641 5583 4675
rect 6929 4641 6963 4675
rect 9045 4641 9079 4675
rect 9413 4641 9447 4675
rect 9965 4641 9999 4675
rect 10149 4641 10183 4675
rect 10517 4641 10551 4675
rect 10609 4641 10643 4675
rect 11161 4641 11195 4675
rect 12173 4641 12207 4675
rect 12440 4641 12474 4675
rect 14565 4641 14599 4675
rect 14749 4641 14783 4675
rect 15577 4641 15611 4675
rect 18613 4641 18647 4675
rect 21281 4641 21315 4675
rect 21465 4641 21499 4675
rect 21833 4641 21867 4675
rect 22017 4641 22051 4675
rect 22281 4641 22315 4675
rect 22477 4641 22511 4675
rect 22569 4641 22603 4675
rect 22753 4641 22787 4675
rect 22845 4641 22879 4675
rect 23489 4641 23523 4675
rect 5641 4573 5675 4607
rect 9781 4573 9815 4607
rect 15485 4573 15519 4607
rect 16681 4573 16715 4607
rect 18889 4573 18923 4607
rect 22385 4573 22419 4607
rect 10793 4505 10827 4539
rect 14289 4505 14323 4539
rect 15945 4505 15979 4539
rect 21005 4505 21039 4539
rect 11253 4437 11287 4471
rect 14105 4437 14139 4471
rect 20821 4437 20855 4471
rect 22109 4437 22143 4471
rect 22569 4437 22603 4471
rect 22937 4437 22971 4471
rect 8217 4233 8251 4267
rect 10793 4233 10827 4267
rect 10977 4233 11011 4267
rect 11253 4233 11287 4267
rect 12633 4233 12667 4267
rect 19625 4233 19659 4267
rect 20913 4233 20947 4267
rect 23673 4233 23707 4267
rect 15669 4165 15703 4199
rect 20361 4165 20395 4199
rect 6469 4097 6503 4131
rect 9045 4097 9079 4131
rect 15209 4097 15243 4131
rect 21925 4097 21959 4131
rect 22201 4097 22235 4131
rect 24869 4097 24903 4131
rect 8401 4029 8435 4063
rect 9137 4029 9171 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 9965 4029 9999 4063
rect 12265 4029 12299 4063
rect 12449 4029 12483 4063
rect 12541 4029 12575 4063
rect 12725 4029 12759 4063
rect 15117 4029 15151 4063
rect 15577 4029 15611 4063
rect 15761 4029 15795 4063
rect 16497 4029 16531 4063
rect 18889 4029 18923 4063
rect 19533 4029 19567 4063
rect 20361 4029 20395 4063
rect 20637 4029 20671 4063
rect 20729 4029 20763 4063
rect 20913 4029 20947 4063
rect 6745 3961 6779 3995
rect 8677 3961 8711 3995
rect 10609 3961 10643 3995
rect 10809 3961 10843 3995
rect 11437 3961 11471 3995
rect 16773 3961 16807 3995
rect 18797 3961 18831 3995
rect 25114 3961 25148 3995
rect 9321 3893 9355 3927
rect 11069 3893 11103 3927
rect 11237 3893 11271 3927
rect 12081 3893 12115 3927
rect 15485 3893 15519 3927
rect 18245 3893 18279 3927
rect 20545 3893 20579 3927
rect 26249 3893 26283 3927
rect 11989 3689 12023 3723
rect 15117 3689 15151 3723
rect 23305 3689 23339 3723
rect 10977 3621 11011 3655
rect 15393 3621 15427 3655
rect 18889 3621 18923 3655
rect 19349 3621 19383 3655
rect 21097 3621 21131 3655
rect 23581 3621 23615 3655
rect 8125 3553 8159 3587
rect 10149 3553 10183 3587
rect 10333 3553 10367 3587
rect 10425 3553 10459 3587
rect 10609 3553 10643 3587
rect 11161 3553 11195 3587
rect 11437 3553 11471 3587
rect 11621 3553 11655 3587
rect 11897 3553 11931 3587
rect 12173 3553 12207 3587
rect 12909 3553 12943 3587
rect 15485 3553 15519 3587
rect 16313 3553 16347 3587
rect 18797 3553 18831 3587
rect 21557 3553 21591 3587
rect 23489 3553 23523 3587
rect 8401 3485 8435 3519
rect 10241 3485 10275 3519
rect 11345 3485 11379 3519
rect 12817 3485 12851 3519
rect 13369 3485 13403 3519
rect 13645 3485 13679 3519
rect 16405 3485 16439 3519
rect 19073 3485 19107 3519
rect 21833 3485 21867 3519
rect 10425 3417 10459 3451
rect 12173 3417 12207 3451
rect 13277 3417 13311 3451
rect 9873 3349 9907 3383
rect 11621 3349 11655 3383
rect 16681 3349 16715 3383
rect 9137 3145 9171 3179
rect 12725 3145 12759 3179
rect 20177 3145 20211 3179
rect 21281 3145 21315 3179
rect 18429 3077 18463 3111
rect 10977 3009 11011 3043
rect 11253 3009 11287 3043
rect 16681 3009 16715 3043
rect 21005 3009 21039 3043
rect 9045 2941 9079 2975
rect 13001 2941 13035 2975
rect 18889 2941 18923 2975
rect 20085 2941 20119 2975
rect 20913 2941 20947 2975
rect 12909 2873 12943 2907
rect 16957 2873 16991 2907
rect 18797 2873 18831 2907
rect 15761 969 15795 1003
rect 16405 969 16439 1003
rect 16865 969 16899 1003
rect 6561 765 6595 799
rect 14289 765 14323 799
rect 15577 765 15611 799
rect 16221 765 16255 799
rect 17049 765 17083 799
rect 18797 765 18831 799
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10413 18819 10471 18825
rect 10413 18816 10425 18819
rect 10376 18788 10425 18816
rect 10376 18776 10382 18788
rect 10413 18785 10425 18788
rect 10459 18785 10471 18819
rect 10413 18779 10471 18785
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 11057 18819 11115 18825
rect 11057 18816 11069 18819
rect 11020 18788 11069 18816
rect 11020 18776 11026 18788
rect 11057 18785 11069 18788
rect 11103 18785 11115 18819
rect 11057 18779 11115 18785
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 12308 18788 12357 18816
rect 12308 18776 12314 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 12989 18819 13047 18825
rect 12989 18816 13001 18819
rect 12952 18788 13001 18816
rect 12952 18776 12958 18788
rect 12989 18785 13001 18788
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 16206 18776 16212 18828
rect 16264 18776 16270 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 18104 18788 18153 18816
rect 18104 18776 18110 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 18690 18776 18696 18828
rect 18748 18816 18754 18828
rect 18785 18819 18843 18825
rect 18785 18816 18797 18819
rect 18748 18788 18797 18816
rect 18748 18776 18754 18788
rect 18785 18785 18797 18788
rect 18831 18785 18843 18819
rect 18785 18779 18843 18785
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19392 18788 19441 18816
rect 19392 18776 19398 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 19429 18779 19487 18785
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 20036 18788 20085 18816
rect 20036 18776 20042 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 20073 18779 20131 18785
rect 20622 18776 20628 18828
rect 20680 18816 20686 18828
rect 20717 18819 20775 18825
rect 20717 18816 20729 18819
rect 20680 18788 20729 18816
rect 20680 18776 20686 18788
rect 20717 18785 20729 18788
rect 20763 18785 20775 18819
rect 20717 18779 20775 18785
rect 21266 18776 21272 18828
rect 21324 18816 21330 18828
rect 21361 18819 21419 18825
rect 21361 18816 21373 18819
rect 21324 18788 21373 18816
rect 21324 18776 21330 18788
rect 21361 18785 21373 18788
rect 21407 18785 21419 18819
rect 21361 18779 21419 18785
rect 21910 18776 21916 18828
rect 21968 18816 21974 18828
rect 22005 18819 22063 18825
rect 22005 18816 22017 18819
rect 21968 18788 22017 18816
rect 21968 18776 21974 18788
rect 22005 18785 22017 18788
rect 22051 18785 22063 18819
rect 22005 18779 22063 18785
rect 31018 18572 31024 18624
rect 31076 18572 31082 18624
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 18230 16776 18236 16788
rect 11532 16748 18236 16776
rect 11532 16720 11560 16748
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 11514 16708 11520 16720
rect 11348 16680 11520 16708
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8996 16612 9045 16640
rect 8996 16600 9002 16612
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 9033 16603 9091 16609
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 10318 16640 10324 16652
rect 9815 16612 10324 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 11348 16649 11376 16680
rect 11514 16668 11520 16680
rect 11572 16668 11578 16720
rect 12618 16668 12624 16720
rect 12676 16668 12682 16720
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 18049 16643 18107 16649
rect 18049 16640 18061 16643
rect 15160 16612 18061 16640
rect 15160 16600 15166 16612
rect 18049 16609 18061 16612
rect 18095 16609 18107 16643
rect 18049 16603 18107 16609
rect 21453 16643 21511 16649
rect 21453 16609 21465 16643
rect 21499 16609 21511 16643
rect 21453 16603 21511 16609
rect 11606 16532 11612 16584
rect 11664 16532 11670 16584
rect 19150 16532 19156 16584
rect 19208 16572 19214 16584
rect 21468 16572 21496 16603
rect 22462 16572 22468 16584
rect 19208 16544 22468 16572
rect 19208 16532 19214 16544
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 9766 16396 9772 16448
rect 9824 16396 9830 16448
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 13081 16439 13139 16445
rect 13081 16436 13093 16439
rect 11480 16408 13093 16436
rect 11480 16396 11486 16408
rect 13081 16405 13093 16408
rect 13127 16405 13139 16439
rect 13081 16399 13139 16405
rect 21542 16396 21548 16448
rect 21600 16396 21606 16448
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 6638 16192 6644 16244
rect 6696 16232 6702 16244
rect 6696 16204 10180 16232
rect 6696 16192 6702 16204
rect 10152 16164 10180 16204
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10413 16235 10471 16241
rect 10413 16232 10425 16235
rect 10376 16204 10425 16232
rect 10376 16192 10382 16204
rect 10413 16201 10425 16204
rect 10459 16201 10471 16235
rect 10413 16195 10471 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11606 16232 11612 16244
rect 11379 16204 11612 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 12529 16235 12587 16241
rect 12529 16201 12541 16235
rect 12575 16232 12587 16235
rect 12618 16232 12624 16244
rect 12575 16204 12624 16232
rect 12575 16201 12587 16204
rect 12529 16195 12587 16201
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 15378 16232 15384 16244
rect 13004 16204 15384 16232
rect 11514 16164 11520 16176
rect 10152 16136 11520 16164
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10152 16105 10180 16136
rect 11514 16124 11520 16136
rect 11572 16124 11578 16176
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9824 16068 9873 16096
rect 9824 16056 9830 16068
rect 9861 16065 9873 16068
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10928 16068 11069 16096
rect 10928 16056 10934 16068
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 12710 16096 12716 16108
rect 11103 16068 12716 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 10229 16031 10287 16037
rect 10229 15997 10241 16031
rect 10275 15997 10287 16031
rect 10229 15991 10287 15997
rect 9122 15920 9128 15972
rect 9180 15920 9186 15972
rect 8389 15895 8447 15901
rect 8389 15861 8401 15895
rect 8435 15892 8447 15895
rect 9030 15892 9036 15904
rect 8435 15864 9036 15892
rect 8435 15861 8447 15864
rect 8389 15855 8447 15861
rect 9030 15852 9036 15864
rect 9088 15892 9094 15904
rect 10244 15892 10272 15991
rect 10410 15988 10416 16040
rect 10468 15988 10474 16040
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11422 16028 11428 16040
rect 11011 16000 11428 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 11422 15988 11428 16000
rect 11480 15988 11486 16040
rect 12621 16031 12679 16037
rect 12621 15997 12633 16031
rect 12667 16028 12679 16031
rect 12802 16028 12808 16040
rect 12667 16000 12808 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 12802 15988 12808 16000
rect 12860 15988 12866 16040
rect 11054 15920 11060 15972
rect 11112 15960 11118 15972
rect 12912 15960 12940 16059
rect 13004 16037 13032 16204
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16558 16235 16616 16241
rect 16558 16232 16570 16235
rect 16163 16204 16570 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16558 16201 16570 16204
rect 16604 16201 16616 16235
rect 16558 16195 16616 16201
rect 15010 16124 15016 16176
rect 15068 16164 15074 16176
rect 15068 16136 16344 16164
rect 15068 16124 15074 16136
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16096 13415 16099
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 13403 16068 13921 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 13909 16065 13921 16068
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 15654 16056 15660 16108
rect 15712 16096 15718 16108
rect 16316 16105 16344 16136
rect 17604 16136 18828 16164
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15712 16068 15761 16096
rect 15712 16056 15718 16068
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 17218 16096 17224 16108
rect 16347 16068 17224 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 17218 16056 17224 16068
rect 17276 16096 17282 16108
rect 17604 16096 17632 16136
rect 17276 16068 17632 16096
rect 17276 16056 17282 16068
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 18288 16068 18705 16096
rect 18288 16056 18294 16068
rect 18693 16065 18705 16068
rect 18739 16065 18751 16099
rect 18800 16096 18828 16136
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 18800 16068 20637 16096
rect 18693 16059 18751 16065
rect 20625 16065 20637 16068
rect 20671 16096 20683 16099
rect 21450 16096 21456 16108
rect 20671 16068 21456 16096
rect 20671 16065 20683 16068
rect 20625 16059 20683 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 22520 16068 22784 16096
rect 22520 16056 22526 16068
rect 12989 16031 13047 16037
rect 12989 15997 13001 16031
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 15997 15899 16031
rect 15841 15991 15899 15997
rect 13538 15960 13544 15972
rect 11112 15932 13544 15960
rect 11112 15920 11118 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 9088 15864 10272 15892
rect 13648 15892 13676 15991
rect 14642 15920 14648 15972
rect 14700 15920 14706 15972
rect 14918 15892 14924 15904
rect 13648 15864 14924 15892
rect 9088 15852 9094 15864
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15856 15892 15884 15991
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 22756 16037 22784 16068
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 18012 16000 18337 16028
rect 18012 15988 18018 16000
rect 18325 15997 18337 16000
rect 18371 16028 18383 16031
rect 22741 16031 22799 16037
rect 18371 16000 18736 16028
rect 18371 15997 18383 16000
rect 18325 15991 18383 15997
rect 18233 15963 18291 15969
rect 18233 15960 18245 15963
rect 17802 15932 18245 15960
rect 18233 15929 18245 15932
rect 18279 15929 18291 15963
rect 18233 15923 18291 15929
rect 18049 15895 18107 15901
rect 18049 15892 18061 15895
rect 15856 15864 18061 15892
rect 18049 15861 18061 15864
rect 18095 15892 18107 15895
rect 18322 15892 18328 15904
rect 18095 15864 18328 15892
rect 18095 15861 18107 15864
rect 18049 15855 18107 15861
rect 18322 15852 18328 15864
rect 18380 15852 18386 15904
rect 18708 15892 18736 16000
rect 22741 15997 22753 16031
rect 22787 15997 22799 16031
rect 22741 15991 22799 15997
rect 18966 15920 18972 15972
rect 19024 15920 19030 15972
rect 19426 15920 19432 15972
rect 19484 15920 19490 15972
rect 20898 15920 20904 15972
rect 20956 15920 20962 15972
rect 21542 15920 21548 15972
rect 21600 15920 21606 15972
rect 19150 15892 19156 15904
rect 18708 15864 19156 15892
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 20441 15895 20499 15901
rect 20441 15892 20453 15895
rect 20312 15864 20453 15892
rect 20312 15852 20318 15864
rect 20441 15861 20453 15864
rect 20487 15861 20499 15895
rect 20441 15855 20499 15861
rect 20530 15852 20536 15904
rect 20588 15892 20594 15904
rect 22373 15895 22431 15901
rect 22373 15892 22385 15895
rect 20588 15864 22385 15892
rect 20588 15852 20594 15864
rect 22373 15861 22385 15864
rect 22419 15861 22431 15895
rect 22373 15855 22431 15861
rect 22830 15852 22836 15904
rect 22888 15852 22894 15904
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 8389 15691 8447 15697
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 8435 15660 8892 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 7926 15580 7932 15632
rect 7984 15580 7990 15632
rect 8665 15555 8723 15561
rect 8665 15521 8677 15555
rect 8711 15552 8723 15555
rect 8711 15524 8800 15552
rect 8711 15521 8723 15524
rect 8665 15515 8723 15521
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6638 15484 6644 15496
rect 6144 15456 6644 15484
rect 6144 15444 6150 15456
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15484 6975 15487
rect 8481 15487 8539 15493
rect 8481 15484 8493 15487
rect 6963 15456 8493 15484
rect 6963 15453 6975 15456
rect 6917 15447 6975 15453
rect 8481 15453 8493 15456
rect 8527 15453 8539 15487
rect 8481 15447 8539 15453
rect 8772 15416 8800 15524
rect 8864 15484 8892 15660
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9088 15660 9904 15688
rect 9088 15648 9094 15660
rect 9876 15629 9904 15660
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 10689 15691 10747 15697
rect 10689 15688 10701 15691
rect 10468 15660 10701 15688
rect 10468 15648 10474 15660
rect 10689 15657 10701 15660
rect 10735 15657 10747 15691
rect 10689 15651 10747 15657
rect 9661 15623 9719 15629
rect 8956 15592 9628 15620
rect 8956 15561 8984 15592
rect 8941 15555 8999 15561
rect 8941 15521 8953 15555
rect 8987 15521 8999 15555
rect 9122 15552 9128 15564
rect 8941 15515 8999 15521
rect 9048 15524 9128 15552
rect 9048 15484 9076 15524
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 9600 15496 9628 15592
rect 9661 15589 9673 15623
rect 9707 15620 9719 15623
rect 9861 15623 9919 15629
rect 9707 15592 9812 15620
rect 9707 15589 9719 15592
rect 9661 15583 9719 15589
rect 9784 15552 9812 15592
rect 9861 15589 9873 15623
rect 9907 15589 9919 15623
rect 10704 15620 10732 15651
rect 11422 15648 11428 15700
rect 11480 15648 11486 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 12618 15688 12624 15700
rect 11756 15660 12624 15688
rect 11756 15648 11762 15660
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 12710 15648 12716 15700
rect 12768 15648 12774 15700
rect 14642 15648 14648 15700
rect 14700 15688 14706 15700
rect 14737 15691 14795 15697
rect 14737 15688 14749 15691
rect 14700 15660 14749 15688
rect 14700 15648 14706 15660
rect 14737 15657 14749 15660
rect 14783 15657 14795 15691
rect 14737 15651 14795 15657
rect 15654 15648 15660 15700
rect 15712 15688 15718 15700
rect 15749 15691 15807 15697
rect 15749 15688 15761 15691
rect 15712 15660 15761 15688
rect 15712 15648 15718 15660
rect 15749 15657 15761 15660
rect 15795 15657 15807 15691
rect 15749 15651 15807 15657
rect 18233 15691 18291 15697
rect 18233 15657 18245 15691
rect 18279 15688 18291 15691
rect 18966 15688 18972 15700
rect 18279 15660 18972 15688
rect 18279 15657 18291 15660
rect 18233 15651 18291 15657
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 19153 15691 19211 15697
rect 19153 15657 19165 15691
rect 19199 15688 19211 15691
rect 19426 15688 19432 15700
rect 19199 15660 19432 15688
rect 19199 15657 19211 15660
rect 19153 15651 19211 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 21361 15691 21419 15697
rect 21361 15657 21373 15691
rect 21407 15688 21419 15691
rect 21407 15660 22140 15688
rect 21407 15657 21419 15660
rect 21361 15651 21419 15657
rect 12728 15620 12756 15648
rect 10704 15592 11744 15620
rect 12728 15592 15332 15620
rect 9861 15583 9919 15589
rect 10502 15552 10508 15564
rect 9784 15524 10508 15552
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 10928 15524 11345 15552
rect 10928 15512 10934 15524
rect 11333 15521 11345 15524
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 11606 15512 11612 15564
rect 11664 15512 11670 15564
rect 11716 15561 11744 15592
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15521 11943 15555
rect 11885 15515 11943 15521
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15521 14703 15555
rect 14645 15515 14703 15521
rect 8864 15456 9076 15484
rect 9582 15444 9588 15496
rect 9640 15444 9646 15496
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 10888 15484 10916 15512
rect 10376 15456 10916 15484
rect 10376 15444 10382 15456
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 11900 15484 11928 15515
rect 11624 15456 11928 15484
rect 11072 15416 11100 15444
rect 11624 15425 11652 15456
rect 8772 15388 11100 15416
rect 11609 15419 11667 15425
rect 11609 15385 11621 15419
rect 11655 15385 11667 15419
rect 11609 15379 11667 15385
rect 12802 15376 12808 15428
rect 12860 15416 12866 15428
rect 13722 15416 13728 15428
rect 12860 15388 13728 15416
rect 12860 15376 12866 15388
rect 13722 15376 13728 15388
rect 13780 15416 13786 15428
rect 14660 15416 14688 15515
rect 15304 15484 15332 15592
rect 15378 15580 15384 15632
rect 15436 15620 15442 15632
rect 22112 15629 22140 15660
rect 20441 15623 20499 15629
rect 20441 15620 20453 15623
rect 15436 15592 15884 15620
rect 15436 15580 15442 15592
rect 15654 15512 15660 15564
rect 15712 15512 15718 15564
rect 15856 15561 15884 15592
rect 18064 15592 20453 15620
rect 15841 15555 15899 15561
rect 15841 15521 15853 15555
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 18064 15484 18092 15592
rect 20441 15589 20453 15592
rect 20487 15620 20499 15623
rect 22097 15623 22155 15629
rect 20487 15592 21312 15620
rect 20487 15589 20499 15592
rect 20441 15583 20499 15589
rect 18325 15555 18383 15561
rect 18325 15552 18337 15555
rect 15304 15456 18092 15484
rect 18156 15524 18337 15552
rect 17954 15416 17960 15428
rect 13780 15388 17960 15416
rect 13780 15376 13786 15388
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 18156 15360 18184 15524
rect 18325 15521 18337 15524
rect 18371 15521 18383 15555
rect 18325 15515 18383 15521
rect 19061 15555 19119 15561
rect 19061 15521 19073 15555
rect 19107 15552 19119 15555
rect 19150 15552 19156 15564
rect 19107 15524 19156 15552
rect 19107 15521 19119 15524
rect 19061 15515 19119 15521
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 19889 15555 19947 15561
rect 19889 15521 19901 15555
rect 19935 15552 19947 15555
rect 20070 15552 20076 15564
rect 19935 15524 20076 15552
rect 19935 15521 19947 15524
rect 19889 15515 19947 15521
rect 20070 15512 20076 15524
rect 20128 15552 20134 15564
rect 20254 15552 20260 15564
rect 20128 15524 20260 15552
rect 20128 15512 20134 15524
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 20622 15512 20628 15564
rect 20680 15512 20686 15564
rect 20806 15512 20812 15564
rect 20864 15512 20870 15564
rect 20990 15512 20996 15564
rect 21048 15512 21054 15564
rect 21284 15561 21312 15592
rect 22097 15589 22109 15623
rect 22143 15589 22155 15623
rect 22097 15583 22155 15589
rect 22830 15580 22836 15632
rect 22888 15580 22894 15632
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15521 21327 15555
rect 21453 15555 21511 15561
rect 21453 15552 21465 15555
rect 21269 15515 21327 15521
rect 21376 15524 21465 15552
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20530 15484 20536 15496
rect 20027 15456 20536 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 20898 15444 20904 15496
rect 20956 15444 20962 15496
rect 21376 15484 21404 15524
rect 21453 15521 21465 15524
rect 21499 15521 21511 15555
rect 21453 15515 21511 15521
rect 23658 15512 23664 15564
rect 23716 15512 23722 15564
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 21008 15456 21404 15484
rect 21468 15456 21833 15484
rect 20257 15419 20315 15425
rect 20257 15385 20269 15419
rect 20303 15416 20315 15419
rect 20916 15416 20944 15444
rect 21008 15425 21036 15456
rect 21468 15428 21496 15456
rect 21821 15453 21833 15456
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 20303 15388 20944 15416
rect 20993 15419 21051 15425
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 20993 15385 21005 15419
rect 21039 15385 21051 15419
rect 20993 15379 21051 15385
rect 21450 15376 21456 15428
rect 21508 15376 21514 15428
rect 23290 15376 23296 15428
rect 23348 15416 23354 15428
rect 23845 15419 23903 15425
rect 23845 15416 23857 15419
rect 23348 15388 23857 15416
rect 23348 15376 23354 15388
rect 23845 15385 23857 15388
rect 23891 15385 23903 15419
rect 23845 15379 23903 15385
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9582 15348 9588 15360
rect 9539 15320 9588 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 9677 15351 9735 15357
rect 9677 15317 9689 15351
rect 9723 15348 9735 15351
rect 10318 15348 10324 15360
rect 9723 15320 10324 15348
rect 9723 15317 9735 15320
rect 9677 15311 9735 15317
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 11790 15308 11796 15360
rect 11848 15348 11854 15360
rect 11885 15351 11943 15357
rect 11885 15348 11897 15351
rect 11848 15320 11897 15348
rect 11848 15308 11854 15320
rect 11885 15317 11897 15320
rect 11931 15317 11943 15351
rect 11885 15311 11943 15317
rect 18138 15308 18144 15360
rect 18196 15308 18202 15360
rect 20346 15308 20352 15360
rect 20404 15348 20410 15360
rect 20806 15348 20812 15360
rect 20404 15320 20812 15348
rect 20404 15308 20410 15320
rect 20806 15308 20812 15320
rect 20864 15348 20870 15360
rect 23569 15351 23627 15357
rect 23569 15348 23581 15351
rect 20864 15320 23581 15348
rect 20864 15308 20870 15320
rect 23569 15317 23581 15320
rect 23615 15348 23627 15351
rect 24118 15348 24124 15360
rect 23615 15320 24124 15348
rect 23615 15317 23627 15320
rect 23569 15311 23627 15317
rect 24118 15308 24124 15320
rect 24176 15308 24182 15360
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 7926 15104 7932 15156
rect 7984 15104 7990 15156
rect 10413 15147 10471 15153
rect 9048 15116 9674 15144
rect 9048 15076 9076 15116
rect 6196 15048 9076 15076
rect 6086 15008 6092 15020
rect 3804 14980 6092 15008
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3804 14949 3832 14980
rect 6086 14968 6092 14980
rect 6144 14968 6150 15020
rect 6196 15017 6224 15048
rect 9122 15036 9128 15088
rect 9180 15036 9186 15088
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6181 14971 6239 14977
rect 9030 14968 9036 15020
rect 9088 14968 9094 15020
rect 9140 15008 9168 15036
rect 9646 15008 9674 15116
rect 10413 15113 10425 15147
rect 10459 15144 10471 15147
rect 10502 15144 10508 15156
rect 10459 15116 10508 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10502 15104 10508 15116
rect 10560 15144 10566 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 10560 15116 11161 15144
rect 10560 15104 10566 15116
rect 11149 15113 11161 15116
rect 11195 15113 11207 15147
rect 15289 15147 15347 15153
rect 11149 15107 11207 15113
rect 11716 15116 15056 15144
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 11716 15076 11744 15116
rect 10192 15048 11744 15076
rect 10192 15036 10198 15048
rect 14918 15008 14924 15020
rect 9140 14980 9352 15008
rect 9646 14980 14924 15008
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 3292 14912 3801 14940
rect 3292 14900 3298 14912
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 6270 14900 6276 14952
rect 6328 14900 6334 14952
rect 6454 14900 6460 14952
rect 6512 14900 6518 14952
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8938 14940 8944 14952
rect 8067 14912 8944 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 8938 14900 8944 14912
rect 8996 14900 9002 14952
rect 9048 14940 9076 14968
rect 9324 14949 9352 14980
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 9048 14912 9137 14940
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 10502 14940 10508 14952
rect 9999 14912 10508 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 10502 14900 10508 14912
rect 10560 14900 10566 14952
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14940 11023 14943
rect 11054 14940 11060 14952
rect 11011 14912 11060 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11333 14943 11391 14949
rect 11333 14909 11345 14943
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 4062 14832 4068 14884
rect 4120 14832 4126 14884
rect 4798 14832 4804 14884
rect 4856 14832 4862 14884
rect 9493 14875 9551 14881
rect 9493 14841 9505 14875
rect 9539 14872 9551 14875
rect 9861 14875 9919 14881
rect 9861 14872 9873 14875
rect 9539 14844 9873 14872
rect 9539 14841 9551 14844
rect 9493 14835 9551 14841
rect 9861 14841 9873 14844
rect 9907 14872 9919 14875
rect 10137 14875 10195 14881
rect 9907 14844 10088 14872
rect 9907 14841 9919 14844
rect 9861 14835 9919 14841
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 5537 14807 5595 14813
rect 5537 14804 5549 14807
rect 4764 14776 5549 14804
rect 4764 14764 4770 14776
rect 5537 14773 5549 14776
rect 5583 14804 5595 14807
rect 6362 14804 6368 14816
rect 5583 14776 6368 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6638 14764 6644 14816
rect 6696 14764 6702 14816
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 9585 14807 9643 14813
rect 9585 14804 9597 14807
rect 7064 14776 9597 14804
rect 7064 14764 7070 14776
rect 9585 14773 9597 14776
rect 9631 14773 9643 14807
rect 9585 14767 9643 14773
rect 9769 14807 9827 14813
rect 9769 14773 9781 14807
rect 9815 14804 9827 14807
rect 9950 14804 9956 14816
rect 9815 14776 9956 14804
rect 9815 14773 9827 14776
rect 9769 14767 9827 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10060 14804 10088 14844
rect 10137 14841 10149 14875
rect 10183 14872 10195 14875
rect 10229 14875 10287 14881
rect 10229 14872 10241 14875
rect 10183 14844 10241 14872
rect 10183 14841 10195 14844
rect 10137 14835 10195 14841
rect 10229 14841 10241 14844
rect 10275 14872 10287 14875
rect 10318 14872 10324 14884
rect 10275 14844 10324 14872
rect 10275 14841 10287 14844
rect 10229 14835 10287 14841
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 10612 14844 10793 14872
rect 10612 14813 10640 14844
rect 10781 14841 10793 14844
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 10429 14807 10487 14813
rect 10429 14804 10441 14807
rect 10060 14776 10441 14804
rect 10429 14773 10441 14776
rect 10475 14773 10487 14807
rect 10429 14767 10487 14773
rect 10597 14807 10655 14813
rect 10597 14773 10609 14807
rect 10643 14773 10655 14807
rect 11348 14804 11376 14903
rect 11422 14900 11428 14952
rect 11480 14900 11486 14952
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 11609 14943 11667 14949
rect 11609 14940 11621 14943
rect 11572 14912 11621 14940
rect 11572 14900 11578 14912
rect 11609 14909 11621 14912
rect 11655 14909 11667 14943
rect 11609 14903 11667 14909
rect 13722 14900 13728 14952
rect 13780 14900 13786 14952
rect 15028 14949 15056 15116
rect 15289 15113 15301 15147
rect 15335 15144 15347 15147
rect 15930 15144 15936 15156
rect 15335 15116 15936 15144
rect 15335 15113 15347 15116
rect 15289 15107 15347 15113
rect 15930 15104 15936 15116
rect 15988 15104 15994 15156
rect 20438 15144 20444 15156
rect 19873 15116 20444 15144
rect 15378 15036 15384 15088
rect 15436 15036 15442 15088
rect 15473 15079 15531 15085
rect 15473 15045 15485 15079
rect 15519 15076 15531 15079
rect 15519 15048 16712 15076
rect 15519 15045 15531 15048
rect 15473 15039 15531 15045
rect 15396 15008 15424 15036
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15396 14980 16129 15008
rect 16117 14977 16129 14980
rect 16163 15008 16175 15011
rect 16298 15008 16304 15020
rect 16163 14980 16304 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 16684 15017 16712 15048
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 19873 15008 19901 15116
rect 20088 15088 20116 15116
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 20530 15104 20536 15156
rect 20588 15104 20594 15156
rect 20622 15104 20628 15156
rect 20680 15104 20686 15156
rect 20901 15147 20959 15153
rect 20901 15113 20913 15147
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 19981 15079 20039 15085
rect 19981 15045 19993 15079
rect 20027 15045 20039 15079
rect 19981 15039 20039 15045
rect 18156 14980 19901 15008
rect 18156 14952 18184 14980
rect 14829 14943 14887 14949
rect 14829 14940 14841 14943
rect 14476 14912 14841 14940
rect 11790 14832 11796 14884
rect 11848 14872 11854 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11848 14844 11897 14872
rect 11848 14832 11854 14844
rect 11885 14841 11897 14844
rect 11931 14841 11943 14875
rect 13633 14875 13691 14881
rect 13633 14872 13645 14875
rect 13110 14844 13645 14872
rect 11885 14835 11943 14841
rect 13633 14841 13645 14844
rect 13679 14841 13691 14875
rect 13633 14835 13691 14841
rect 11606 14804 11612 14816
rect 11348 14776 11612 14804
rect 10597 14767 10655 14773
rect 11606 14764 11612 14776
rect 11664 14804 11670 14816
rect 13354 14804 13360 14816
rect 11664 14776 13360 14804
rect 11664 14764 11670 14776
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 14476 14804 14504 14912
rect 14829 14909 14841 14912
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 15013 14943 15071 14949
rect 15013 14909 15025 14943
rect 15059 14940 15071 14943
rect 16206 14940 16212 14952
rect 15059 14912 16212 14940
rect 15059 14909 15071 14912
rect 15013 14903 15071 14909
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 16758 14900 16764 14952
rect 16816 14900 16822 14952
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14940 17463 14943
rect 17494 14940 17500 14952
rect 17451 14912 17500 14940
rect 17451 14909 17463 14912
rect 17405 14903 17463 14909
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 18138 14900 18144 14952
rect 18196 14900 18202 14952
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 18693 14943 18751 14949
rect 18693 14940 18705 14943
rect 18555 14912 18705 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 18693 14909 18705 14912
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 15105 14875 15163 14881
rect 15105 14841 15117 14875
rect 15151 14872 15163 14875
rect 15194 14872 15200 14884
rect 15151 14844 15200 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 15654 14872 15660 14884
rect 15488 14844 15660 14872
rect 15305 14807 15363 14813
rect 15305 14804 15317 14807
rect 13596 14776 15317 14804
rect 13596 14764 13602 14776
rect 15305 14773 15317 14776
rect 15351 14804 15363 14807
rect 15488 14804 15516 14844
rect 15654 14832 15660 14844
rect 15712 14872 15718 14884
rect 15749 14875 15807 14881
rect 15749 14872 15761 14875
rect 15712 14844 15761 14872
rect 15712 14832 15718 14844
rect 15749 14841 15761 14844
rect 15795 14841 15807 14875
rect 15749 14835 15807 14841
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14872 15899 14875
rect 16776 14872 16804 14900
rect 15887 14844 16804 14872
rect 15887 14841 15899 14844
rect 15841 14835 15899 14841
rect 15351 14776 15516 14804
rect 15351 14773 15363 14776
rect 15305 14767 15363 14773
rect 15562 14764 15568 14816
rect 15620 14764 15626 14816
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16574 14804 16580 14816
rect 15988 14776 16580 14804
rect 15988 14764 15994 14776
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 17313 14807 17371 14813
rect 17313 14773 17325 14807
rect 17359 14804 17371 14807
rect 17586 14804 17592 14816
rect 17359 14776 17592 14804
rect 17359 14773 17371 14776
rect 17313 14767 17371 14773
rect 17586 14764 17592 14776
rect 17644 14764 17650 14816
rect 18414 14764 18420 14816
rect 18472 14764 18478 14816
rect 18708 14804 18736 14903
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 19812 14949 19840 14980
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 18840 14912 19257 14940
rect 18840 14900 18846 14912
rect 19245 14909 19257 14912
rect 19291 14909 19303 14943
rect 19245 14903 19303 14909
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14909 19763 14943
rect 19705 14903 19763 14909
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 18969 14875 19027 14881
rect 18969 14841 18981 14875
rect 19015 14872 19027 14875
rect 19150 14872 19156 14884
rect 19015 14844 19156 14872
rect 19015 14841 19027 14844
rect 18969 14835 19027 14841
rect 19150 14832 19156 14844
rect 19208 14832 19214 14884
rect 19720 14872 19748 14903
rect 19886 14900 19892 14952
rect 19944 14900 19950 14952
rect 19996 14940 20024 15039
rect 20070 15036 20076 15088
rect 20128 15036 20134 15088
rect 20254 15036 20260 15088
rect 20312 15076 20318 15088
rect 20548 15076 20576 15104
rect 20916 15076 20944 15107
rect 20990 15104 20996 15156
rect 21048 15144 21054 15156
rect 21085 15147 21143 15153
rect 21085 15144 21097 15147
rect 21048 15116 21097 15144
rect 21048 15104 21054 15116
rect 21085 15113 21097 15116
rect 21131 15113 21143 15147
rect 21085 15107 21143 15113
rect 20312 15048 20944 15076
rect 20312 15036 20318 15048
rect 21100 15008 21128 15107
rect 20732 14980 20944 15008
rect 21100 14980 21404 15008
rect 20732 14940 20760 14980
rect 19996 14934 20576 14940
rect 20664 14934 20760 14940
rect 19996 14912 20760 14934
rect 20916 14940 20944 14980
rect 21376 14949 21404 14980
rect 21450 14968 21456 15020
rect 21508 15008 21514 15020
rect 21637 15011 21695 15017
rect 21637 15008 21649 15011
rect 21508 14980 21649 15008
rect 21508 14968 21514 14980
rect 21637 14977 21649 14980
rect 21683 14977 21695 15011
rect 21637 14971 21695 14977
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 20916 14912 21189 14940
rect 20548 14906 20692 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14909 21419 14943
rect 21361 14903 21419 14909
rect 23845 14943 23903 14949
rect 23845 14909 23857 14943
rect 23891 14940 23903 14943
rect 23934 14940 23940 14952
rect 23891 14912 23940 14940
rect 23891 14909 23903 14912
rect 23845 14903 23903 14909
rect 23934 14900 23940 14912
rect 23992 14900 23998 14952
rect 24118 14949 24124 14952
rect 24112 14903 24124 14949
rect 24118 14900 24124 14903
rect 24176 14900 24182 14952
rect 19904 14872 19932 14900
rect 19720 14844 19932 14872
rect 19981 14875 20039 14881
rect 19981 14841 19993 14875
rect 20027 14872 20039 14875
rect 20349 14875 20407 14881
rect 20349 14872 20361 14875
rect 20027 14844 20361 14872
rect 20027 14841 20039 14844
rect 19981 14835 20039 14841
rect 20349 14841 20361 14844
rect 20395 14872 20407 14875
rect 20395 14844 20576 14872
rect 20395 14841 20407 14844
rect 20349 14835 20407 14841
rect 19426 14804 19432 14816
rect 18708 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 20254 14764 20260 14816
rect 20312 14764 20318 14816
rect 20438 14764 20444 14816
rect 20496 14764 20502 14816
rect 20548 14804 20576 14844
rect 20714 14832 20720 14884
rect 20772 14832 20778 14884
rect 21269 14875 21327 14881
rect 21269 14841 21281 14875
rect 21315 14872 21327 14875
rect 21913 14875 21971 14881
rect 21913 14872 21925 14875
rect 21315 14844 21925 14872
rect 21315 14841 21327 14844
rect 21269 14835 21327 14841
rect 21913 14841 21925 14844
rect 21959 14841 21971 14875
rect 21913 14835 21971 14841
rect 22646 14832 22652 14884
rect 22704 14832 22710 14884
rect 20927 14807 20985 14813
rect 20927 14804 20939 14807
rect 20548 14776 20939 14804
rect 20927 14773 20939 14776
rect 20973 14804 20985 14807
rect 23385 14807 23443 14813
rect 23385 14804 23397 14807
rect 20973 14776 23397 14804
rect 20973 14773 20985 14776
rect 20927 14767 20985 14773
rect 23385 14773 23397 14776
rect 23431 14804 23443 14807
rect 23842 14804 23848 14816
rect 23431 14776 23848 14804
rect 23431 14773 23443 14776
rect 23385 14767 23443 14773
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 25038 14764 25044 14816
rect 25096 14804 25102 14816
rect 25225 14807 25283 14813
rect 25225 14804 25237 14807
rect 25096 14776 25237 14804
rect 25096 14764 25102 14776
rect 25225 14773 25237 14776
rect 25271 14773 25283 14807
rect 25225 14767 25283 14773
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 4893 14603 4951 14609
rect 4893 14600 4905 14603
rect 4856 14572 4905 14600
rect 4856 14560 4862 14572
rect 4893 14569 4905 14572
rect 4939 14569 4951 14603
rect 4893 14563 4951 14569
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6270 14600 6276 14612
rect 6227 14572 6276 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 6362 14560 6368 14612
rect 6420 14560 6426 14612
rect 6638 14600 6644 14612
rect 6564 14572 6644 14600
rect 3418 14532 3424 14544
rect 2608 14504 3424 14532
rect 842 14424 848 14476
rect 900 14424 906 14476
rect 2608 14473 2636 14504
rect 3418 14492 3424 14504
rect 3476 14532 3482 14544
rect 6380 14532 6408 14560
rect 6564 14541 6592 14572
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 6788 14572 8064 14600
rect 6788 14560 6794 14572
rect 3476 14504 6132 14532
rect 3476 14492 3482 14504
rect 2593 14467 2651 14473
rect 2593 14433 2605 14467
rect 2639 14433 2651 14467
rect 2593 14427 2651 14433
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 3142 14464 3148 14476
rect 2823 14436 3148 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3605 14467 3663 14473
rect 3605 14433 3617 14467
rect 3651 14464 3663 14467
rect 3651 14436 3924 14464
rect 3651 14433 3663 14436
rect 3605 14427 3663 14433
rect 3694 14356 3700 14408
rect 3752 14356 3758 14408
rect 2406 14288 2412 14340
rect 2464 14328 2470 14340
rect 2961 14331 3019 14337
rect 2961 14328 2973 14331
rect 2464 14300 2973 14328
rect 2464 14288 2470 14300
rect 2961 14297 2973 14300
rect 3007 14297 3019 14331
rect 3896 14328 3924 14436
rect 4062 14424 4068 14476
rect 4120 14424 4126 14476
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14464 4859 14467
rect 4890 14464 4896 14476
rect 4847 14436 4896 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 5997 14467 6055 14473
rect 5997 14433 6009 14467
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4080 14396 4108 14424
rect 4019 14368 4108 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4706 14328 4712 14340
rect 3896 14300 4712 14328
rect 2961 14291 3019 14297
rect 1029 14263 1087 14269
rect 1029 14260 1041 14263
rect 492 14232 1041 14260
rect 492 14056 520 14232
rect 1029 14229 1041 14232
rect 1075 14229 1087 14263
rect 2976 14260 3004 14291
rect 4706 14288 4712 14300
rect 4764 14288 4770 14340
rect 4798 14260 4804 14272
rect 2976 14232 4804 14260
rect 1029 14223 1087 14229
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 6012 14260 6040 14427
rect 6104 14396 6132 14504
rect 6196 14504 6408 14532
rect 6549 14535 6607 14541
rect 6196 14473 6224 14504
rect 6549 14501 6561 14535
rect 6595 14501 6607 14535
rect 6549 14495 6607 14501
rect 7558 14492 7564 14544
rect 7616 14492 7622 14544
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14433 6239 14467
rect 6181 14427 6239 14433
rect 6270 14424 6276 14476
rect 6328 14424 6334 14476
rect 8036 14464 8064 14572
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 8996 14572 10272 14600
rect 8996 14560 9002 14572
rect 8472 14535 8530 14541
rect 8472 14501 8484 14535
rect 8518 14532 8530 14535
rect 9122 14532 9128 14544
rect 8518 14504 9128 14532
rect 8518 14501 8530 14504
rect 8472 14495 8530 14501
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 8036 14436 10149 14464
rect 6638 14396 6644 14408
rect 6104 14368 6644 14396
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 8205 14399 8263 14405
rect 8205 14396 8217 14399
rect 6972 14368 8217 14396
rect 6972 14356 6978 14368
rect 8205 14365 8217 14368
rect 8251 14365 8263 14399
rect 10060 14396 10088 14436
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 10244 14464 10272 14572
rect 11422 14560 11428 14612
rect 11480 14560 11486 14612
rect 13354 14560 13360 14612
rect 13412 14560 13418 14612
rect 15010 14560 15016 14612
rect 15068 14560 15074 14612
rect 16114 14560 16120 14612
rect 16172 14560 16178 14612
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 16264 14572 16681 14600
rect 16264 14560 16270 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 16669 14563 16727 14569
rect 17126 14560 17132 14612
rect 17184 14600 17190 14612
rect 17184 14572 17724 14600
rect 17184 14560 17190 14572
rect 11440 14532 11468 14560
rect 11578 14535 11636 14541
rect 11578 14532 11590 14535
rect 11440 14504 11590 14532
rect 11578 14501 11590 14504
rect 11624 14501 11636 14535
rect 13372 14532 13400 14560
rect 13510 14535 13568 14541
rect 13510 14532 13522 14535
rect 13372 14504 13522 14532
rect 11578 14495 11636 14501
rect 13510 14501 13522 14504
rect 13556 14501 13568 14535
rect 13510 14495 13568 14501
rect 14936 14504 15516 14532
rect 14936 14476 14964 14504
rect 12802 14464 12808 14476
rect 10244 14436 12808 14464
rect 10137 14427 10195 14433
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 14918 14424 14924 14476
rect 14976 14424 14982 14476
rect 15102 14424 15108 14476
rect 15160 14424 15166 14476
rect 15488 14473 15516 14504
rect 15562 14492 15568 14544
rect 15620 14492 15626 14544
rect 16132 14532 16160 14560
rect 16301 14535 16359 14541
rect 16301 14532 16313 14535
rect 16132 14504 16313 14532
rect 16301 14501 16313 14504
rect 16347 14501 16359 14535
rect 16301 14495 16359 14501
rect 16393 14535 16451 14541
rect 16393 14501 16405 14535
rect 16439 14532 16451 14535
rect 16758 14532 16764 14544
rect 16439 14504 16764 14532
rect 16439 14501 16451 14504
rect 16393 14495 16451 14501
rect 16758 14492 16764 14504
rect 16816 14532 16822 14544
rect 17586 14532 17592 14544
rect 16816 14504 17172 14532
rect 16816 14492 16822 14504
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 11238 14396 11244 14408
rect 10060 14368 11244 14396
rect 8205 14359 8263 14365
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 13262 14396 13268 14408
rect 11333 14359 11391 14365
rect 12406 14368 13268 14396
rect 7650 14260 7656 14272
rect 6012 14232 7656 14260
rect 7650 14220 7656 14232
rect 7708 14260 7714 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 7708 14232 8033 14260
rect 7708 14220 7714 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8021 14223 8079 14229
rect 9585 14263 9643 14269
rect 9585 14229 9597 14263
rect 9631 14260 9643 14263
rect 9766 14260 9772 14272
rect 9631 14232 9772 14260
rect 9631 14229 9643 14232
rect 9585 14223 9643 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 9953 14263 10011 14269
rect 9953 14260 9965 14263
rect 9916 14232 9965 14260
rect 9916 14220 9922 14232
rect 9953 14229 9965 14232
rect 9999 14260 10011 14263
rect 11348 14260 11376 14359
rect 12406 14260 12434 14368
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 15580 14396 15608 14492
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 16206 14464 16212 14476
rect 16163 14436 16212 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16482 14464 16488 14476
rect 16408 14436 16488 14464
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 15580 14368 15669 14396
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 16408 14396 16436 14436
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 15795 14368 16436 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 15194 14328 15200 14340
rect 14660 14300 15200 14328
rect 9999 14232 12434 14260
rect 9999 14229 10011 14232
rect 9953 14223 10011 14229
rect 12710 14220 12716 14272
rect 12768 14220 12774 14272
rect 14660 14269 14688 14300
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 17144 14328 17172 14504
rect 17328 14504 17592 14532
rect 17218 14424 17224 14476
rect 17276 14424 17282 14476
rect 17328 14473 17356 14504
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 17696 14541 17724 14572
rect 22646 14560 22652 14612
rect 22704 14560 22710 14612
rect 17681 14535 17739 14541
rect 17681 14501 17693 14535
rect 17727 14501 17739 14535
rect 17681 14495 17739 14501
rect 18414 14492 18420 14544
rect 18472 14492 18478 14544
rect 23216 14504 23796 14532
rect 23216 14476 23244 14504
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14433 17371 14467
rect 17313 14427 17371 14433
rect 22462 14424 22468 14476
rect 22520 14464 22526 14476
rect 22557 14467 22615 14473
rect 22557 14464 22569 14467
rect 22520 14436 22569 14464
rect 22520 14424 22526 14436
rect 22557 14433 22569 14436
rect 22603 14433 22615 14467
rect 22557 14427 22615 14433
rect 23198 14424 23204 14476
rect 23256 14424 23262 14476
rect 23290 14424 23296 14476
rect 23348 14424 23354 14476
rect 23400 14473 23428 14504
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14433 23443 14467
rect 23641 14467 23699 14473
rect 23641 14464 23653 14467
rect 23385 14427 23443 14433
rect 23483 14436 23653 14464
rect 17236 14396 17264 14424
rect 17405 14399 17463 14405
rect 17405 14396 17417 14399
rect 17236 14368 17417 14396
rect 17405 14365 17417 14368
rect 17451 14365 17463 14399
rect 19153 14399 19211 14405
rect 19153 14396 19165 14399
rect 17405 14359 17463 14365
rect 17512 14368 19165 14396
rect 17512 14328 17540 14368
rect 19153 14365 19165 14368
rect 19199 14396 19211 14399
rect 23483 14396 23511 14436
rect 23641 14433 23653 14436
rect 23687 14433 23699 14467
rect 23768 14464 23796 14504
rect 23842 14492 23848 14544
rect 23900 14532 23906 14544
rect 25102 14535 25160 14541
rect 25102 14532 25114 14535
rect 23900 14504 25114 14532
rect 23900 14492 23906 14504
rect 25102 14501 25114 14504
rect 25148 14501 25160 14535
rect 25102 14495 25160 14501
rect 23934 14464 23940 14476
rect 23768 14436 23940 14464
rect 23641 14427 23699 14433
rect 23934 14424 23940 14436
rect 23992 14464 23998 14476
rect 24857 14467 24915 14473
rect 24857 14464 24869 14467
rect 23992 14436 24869 14464
rect 23992 14424 23998 14436
rect 24857 14433 24869 14436
rect 24903 14433 24915 14467
rect 24857 14427 24915 14433
rect 19199 14368 23511 14396
rect 19199 14365 19211 14368
rect 19153 14359 19211 14365
rect 17144 14300 17540 14328
rect 14645 14263 14703 14269
rect 14645 14229 14657 14263
rect 14691 14229 14703 14263
rect 14645 14223 14703 14229
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15102 14260 15108 14272
rect 14884 14232 15108 14260
rect 14884 14220 14890 14232
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 15286 14220 15292 14272
rect 15344 14220 15350 14272
rect 17129 14263 17187 14269
rect 17129 14229 17141 14263
rect 17175 14260 17187 14263
rect 18690 14260 18696 14272
rect 17175 14232 18696 14260
rect 17175 14229 17187 14232
rect 17129 14223 17187 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 23109 14263 23167 14269
rect 23109 14229 23121 14263
rect 23155 14260 23167 14263
rect 23198 14260 23204 14272
rect 23155 14232 23204 14260
rect 23155 14229 23167 14232
rect 23109 14223 23167 14229
rect 23198 14220 23204 14232
rect 23256 14220 23262 14272
rect 24765 14263 24823 14269
rect 24765 14229 24777 14263
rect 24811 14260 24823 14263
rect 25498 14260 25504 14272
rect 24811 14232 25504 14260
rect 24811 14229 24823 14232
rect 24765 14223 24823 14229
rect 25498 14220 25504 14232
rect 25556 14220 25562 14272
rect 26234 14220 26240 14272
rect 26292 14220 26298 14272
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 492 14028 3280 14056
rect 2406 13948 2412 14000
rect 2464 13948 2470 14000
rect 2501 13991 2559 13997
rect 2501 13957 2513 13991
rect 2547 13957 2559 13991
rect 2501 13951 2559 13957
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2424 13852 2452 13948
rect 2363 13824 2452 13852
rect 2516 13852 2544 13951
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 2516 13824 2605 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 3252 13861 3280 14028
rect 3418 14016 3424 14068
rect 3476 14016 3482 14068
rect 3694 14016 3700 14068
rect 3752 14056 3758 14068
rect 4338 14056 4344 14068
rect 3752 14028 4344 14056
rect 3752 14016 3758 14028
rect 4338 14016 4344 14028
rect 4396 14056 4402 14068
rect 7006 14056 7012 14068
rect 4396 14028 7012 14056
rect 4396 14016 4402 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 7558 14056 7564 14068
rect 7515 14028 7564 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 13262 14016 13268 14068
rect 13320 14016 13326 14068
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 15378 14056 15384 14068
rect 13964 14028 14964 14056
rect 13964 14016 13970 14028
rect 3712 13861 3740 14016
rect 4706 13988 4712 14000
rect 3896 13960 4712 13988
rect 3896 13929 3924 13960
rect 4706 13948 4712 13960
rect 4764 13948 4770 14000
rect 6365 13991 6423 13997
rect 6365 13957 6377 13991
rect 6411 13988 6423 13991
rect 8018 13988 8024 14000
rect 6411 13960 8024 13988
rect 6411 13957 6423 13960
rect 6365 13951 6423 13957
rect 8018 13948 8024 13960
rect 8076 13948 8082 14000
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 3988 13892 5120 13920
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13821 3295 13855
rect 3237 13815 3295 13821
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 3789 13787 3847 13793
rect 3789 13753 3801 13787
rect 3835 13784 3847 13787
rect 3988 13784 4016 13892
rect 4540 13861 4568 13892
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4525 13855 4583 13861
rect 4111 13824 4476 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 3835 13756 4016 13784
rect 3835 13753 3847 13756
rect 3789 13747 3847 13753
rect 4338 13744 4344 13796
rect 4396 13744 4402 13796
rect 4448 13793 4476 13824
rect 4525 13821 4537 13855
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 4798 13812 4804 13864
rect 4856 13852 4862 13864
rect 4982 13852 4988 13864
rect 4856 13824 4988 13852
rect 4856 13812 4862 13824
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5092 13852 5120 13892
rect 6454 13880 6460 13932
rect 6512 13880 6518 13932
rect 13280 13920 13308 14016
rect 14936 13997 14964 14028
rect 15028 14028 15384 14056
rect 14921 13991 14979 13997
rect 14921 13957 14933 13991
rect 14967 13957 14979 13991
rect 14921 13951 14979 13957
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 6656 13892 7696 13920
rect 6656 13861 6684 13892
rect 7668 13864 7696 13892
rect 9048 13892 9996 13920
rect 13280 13892 13553 13920
rect 9048 13864 9076 13892
rect 6641 13855 6699 13861
rect 6641 13852 6653 13855
rect 5092 13824 6653 13852
rect 6641 13821 6653 13824
rect 6687 13821 6699 13855
rect 6641 13815 6699 13821
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13852 6975 13855
rect 7006 13852 7012 13864
rect 6963 13824 7012 13852
rect 6963 13821 6975 13824
rect 6917 13815 6975 13821
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 7156 13824 7389 13852
rect 7156 13812 7162 13824
rect 7377 13821 7389 13824
rect 7423 13821 7435 13855
rect 7377 13815 7435 13821
rect 7650 13812 7656 13864
rect 7708 13812 7714 13864
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9858 13812 9864 13864
rect 9916 13812 9922 13864
rect 9968 13852 9996 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 15028 13920 15056 14028
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 18690 14016 18696 14068
rect 18748 14056 18754 14068
rect 19058 14056 19064 14068
rect 18748 14028 19064 14056
rect 18748 14016 18754 14028
rect 19058 14016 19064 14028
rect 19116 14056 19122 14068
rect 19116 14028 21588 14056
rect 19116 14016 19122 14028
rect 16482 13948 16488 14000
rect 16540 13988 16546 14000
rect 16540 13960 16712 13988
rect 16540 13948 16546 13960
rect 13541 13883 13599 13889
rect 14936 13892 15056 13920
rect 10117 13855 10175 13861
rect 10117 13852 10129 13855
rect 9968 13824 10129 13852
rect 10117 13821 10129 13824
rect 10163 13821 10175 13855
rect 10117 13815 10175 13821
rect 13808 13855 13866 13861
rect 13808 13821 13820 13855
rect 13854 13852 13866 13855
rect 14936 13852 14964 13892
rect 15286 13880 15292 13932
rect 15344 13880 15350 13932
rect 13854 13824 14964 13852
rect 13854 13821 13866 13824
rect 13808 13815 13866 13821
rect 15010 13812 15016 13864
rect 15068 13812 15074 13864
rect 16684 13852 16712 13960
rect 21560 13929 21588 14028
rect 23017 13991 23075 13997
rect 23017 13957 23029 13991
rect 23063 13957 23075 13991
rect 23017 13951 23075 13957
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13889 16819 13923
rect 21545 13923 21603 13929
rect 16761 13883 16819 13889
rect 18340 13892 18828 13920
rect 16776 13852 16804 13883
rect 18340 13852 18368 13892
rect 16684 13824 18368 13852
rect 18417 13855 18475 13861
rect 18417 13821 18429 13855
rect 18463 13852 18475 13855
rect 18690 13852 18696 13864
rect 18463 13824 18696 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 18800 13852 18828 13892
rect 21545 13889 21557 13923
rect 21591 13920 21603 13923
rect 21637 13923 21695 13929
rect 21637 13920 21649 13923
rect 21591 13892 21649 13920
rect 21591 13889 21603 13892
rect 21545 13883 21603 13889
rect 21637 13889 21649 13892
rect 21683 13889 21695 13923
rect 23032 13920 23060 13951
rect 23032 13892 24808 13920
rect 21637 13883 21695 13889
rect 21893 13855 21951 13861
rect 21893 13852 21905 13855
rect 18800 13824 21496 13852
rect 4433 13787 4491 13793
rect 4433 13753 4445 13787
rect 4479 13784 4491 13787
rect 5230 13787 5288 13793
rect 5230 13784 5242 13787
rect 4479 13756 4666 13784
rect 4479 13753 4491 13756
rect 4433 13747 4491 13753
rect 2774 13676 2780 13728
rect 2832 13676 2838 13728
rect 3050 13676 3056 13728
rect 3108 13676 3114 13728
rect 3973 13719 4031 13725
rect 3973 13685 3985 13719
rect 4019 13716 4031 13719
rect 4062 13716 4068 13728
rect 4019 13688 4068 13716
rect 4019 13685 4031 13688
rect 3973 13679 4031 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4157 13719 4215 13725
rect 4157 13685 4169 13719
rect 4203 13716 4215 13719
rect 4246 13716 4252 13728
rect 4203 13688 4252 13716
rect 4203 13685 4215 13688
rect 4157 13679 4215 13685
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 4638 13716 4666 13756
rect 5000 13756 5242 13784
rect 5000 13728 5028 13756
rect 5230 13753 5242 13756
rect 5276 13753 5288 13787
rect 5230 13747 5288 13753
rect 12894 13744 12900 13796
rect 12952 13784 12958 13796
rect 15562 13784 15568 13796
rect 12952 13756 15568 13784
rect 12952 13744 12958 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 15746 13744 15752 13796
rect 15804 13744 15810 13796
rect 18138 13744 18144 13796
rect 18196 13793 18202 13796
rect 18196 13747 18208 13793
rect 18196 13744 18202 13747
rect 18322 13744 18328 13796
rect 18380 13784 18386 13796
rect 18938 13787 18996 13793
rect 18938 13784 18950 13787
rect 18380 13756 18950 13784
rect 18380 13744 18386 13756
rect 18938 13753 18950 13756
rect 18984 13753 18996 13787
rect 18938 13747 18996 13753
rect 20254 13744 20260 13796
rect 20312 13784 20318 13796
rect 21278 13787 21336 13793
rect 21278 13784 21290 13787
rect 20312 13756 21290 13784
rect 20312 13744 20318 13756
rect 21278 13753 21290 13756
rect 21324 13753 21336 13787
rect 21468 13784 21496 13824
rect 21744 13824 21905 13852
rect 21744 13784 21772 13824
rect 21893 13821 21905 13824
rect 21939 13821 21951 13855
rect 21893 13815 21951 13821
rect 24486 13812 24492 13864
rect 24544 13852 24550 13864
rect 24780 13861 24808 13892
rect 24673 13855 24731 13861
rect 24673 13852 24685 13855
rect 24544 13824 24685 13852
rect 24544 13812 24550 13824
rect 24673 13821 24685 13824
rect 24719 13821 24731 13855
rect 24673 13815 24731 13821
rect 24766 13855 24824 13861
rect 24766 13821 24778 13855
rect 24812 13821 24824 13855
rect 24766 13815 24824 13821
rect 25038 13812 25044 13864
rect 25096 13812 25102 13864
rect 25130 13812 25136 13864
rect 25188 13861 25194 13864
rect 25188 13852 25196 13861
rect 25188 13824 25233 13852
rect 25188 13815 25196 13824
rect 25188 13812 25194 13815
rect 21468 13756 21772 13784
rect 21278 13747 21336 13753
rect 23290 13744 23296 13796
rect 23348 13784 23354 13796
rect 24394 13784 24400 13796
rect 23348 13756 24400 13784
rect 23348 13744 23354 13756
rect 24394 13744 24400 13756
rect 24452 13744 24458 13796
rect 24946 13744 24952 13796
rect 25004 13744 25010 13796
rect 4982 13716 4988 13728
rect 4638 13688 4988 13716
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6822 13716 6828 13728
rect 6420 13688 6828 13716
rect 6420 13676 6426 13688
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 11241 13719 11299 13725
rect 11241 13685 11253 13719
rect 11287 13716 11299 13719
rect 11514 13716 11520 13728
rect 11287 13688 11520 13716
rect 11287 13685 11299 13688
rect 11241 13679 11299 13685
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 14734 13676 14740 13728
rect 14792 13716 14798 13728
rect 17037 13719 17095 13725
rect 17037 13716 17049 13719
rect 14792 13688 17049 13716
rect 14792 13676 14798 13688
rect 17037 13685 17049 13688
rect 17083 13685 17095 13719
rect 17037 13679 17095 13685
rect 20070 13676 20076 13728
rect 20128 13676 20134 13728
rect 20165 13719 20223 13725
rect 20165 13685 20177 13719
rect 20211 13716 20223 13719
rect 20530 13716 20536 13728
rect 20211 13688 20536 13716
rect 20211 13685 20223 13688
rect 20165 13679 20223 13685
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 20622 13676 20628 13728
rect 20680 13716 20686 13728
rect 24854 13716 24860 13728
rect 20680 13688 24860 13716
rect 20680 13676 20686 13688
rect 24854 13676 24860 13688
rect 24912 13676 24918 13728
rect 25317 13719 25375 13725
rect 25317 13685 25329 13719
rect 25363 13716 25375 13719
rect 25590 13716 25596 13728
rect 25363 13688 25596 13716
rect 25363 13685 25375 13688
rect 25317 13679 25375 13685
rect 25590 13676 25596 13688
rect 25648 13676 25654 13728
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 2774 13472 2780 13524
rect 2832 13472 2838 13524
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2924 13484 2973 13512
rect 2924 13472 2930 13484
rect 2961 13481 2973 13484
rect 3007 13481 3019 13515
rect 2961 13475 3019 13481
rect 3050 13472 3056 13524
rect 3108 13472 3114 13524
rect 3329 13515 3387 13521
rect 3329 13481 3341 13515
rect 3375 13481 3387 13515
rect 3329 13475 3387 13481
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10091 13484 10272 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 2792 13385 2820 13472
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13345 2835 13379
rect 3068 13376 3096 13472
rect 3344 13444 3372 13475
rect 3881 13447 3939 13453
rect 3881 13444 3893 13447
rect 3344 13416 3893 13444
rect 3881 13413 3893 13416
rect 3927 13413 3939 13447
rect 3881 13407 3939 13413
rect 7460 13447 7518 13453
rect 7460 13413 7472 13447
rect 7506 13444 7518 13447
rect 7650 13444 7656 13456
rect 7506 13416 7656 13444
rect 7506 13413 7518 13416
rect 7460 13407 7518 13413
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 8036 13416 10180 13444
rect 8036 13388 8064 13416
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 3068 13348 3157 13376
rect 2777 13339 2835 13345
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 3697 13379 3755 13385
rect 3697 13345 3709 13379
rect 3743 13376 3755 13379
rect 3743 13348 4108 13376
rect 3743 13345 3755 13348
rect 3697 13339 3755 13345
rect 4080 13252 4108 13348
rect 4154 13336 4160 13388
rect 4212 13336 4218 13388
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4341 13379 4399 13385
rect 4341 13376 4353 13379
rect 4304 13348 4353 13376
rect 4304 13336 4310 13348
rect 4341 13345 4353 13348
rect 4387 13376 4399 13379
rect 4706 13376 4712 13388
rect 4387 13348 4712 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 8018 13336 8024 13388
rect 8076 13336 8082 13388
rect 8754 13336 8760 13388
rect 8812 13376 8818 13388
rect 8921 13379 8979 13385
rect 8921 13376 8933 13379
rect 8812 13348 8933 13376
rect 8812 13336 8818 13348
rect 8921 13345 8933 13348
rect 8967 13345 8979 13379
rect 8921 13339 8979 13345
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 10152 13385 10180 13416
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10244 13376 10272 13484
rect 10594 13472 10600 13524
rect 10652 13512 10658 13524
rect 14921 13515 14979 13521
rect 10652 13484 12848 13512
rect 10652 13472 10658 13484
rect 10318 13404 10324 13456
rect 10376 13444 10382 13456
rect 10376 13416 12664 13444
rect 10376 13404 10382 13416
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10244 13348 10425 13376
rect 10137 13339 10195 13345
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 10505 13379 10563 13385
rect 10505 13345 10517 13379
rect 10551 13376 10563 13379
rect 10778 13376 10784 13388
rect 10551 13348 10784 13376
rect 10551 13345 10563 13348
rect 10505 13339 10563 13345
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 11238 13385 11244 13388
rect 11232 13339 11244 13385
rect 11238 13336 11244 13339
rect 11296 13336 11302 13388
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 12636 13385 12664 13416
rect 12710 13404 12716 13456
rect 12768 13404 12774 13456
rect 12820 13444 12848 13484
rect 14921 13481 14933 13515
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 14936 13444 14964 13475
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 15620 13484 19334 13512
rect 15620 13472 15626 13484
rect 15289 13447 15347 13453
rect 15289 13444 15301 13447
rect 12820 13416 14228 13444
rect 14936 13416 15301 13444
rect 12437 13382 12495 13385
rect 12360 13379 12495 13382
rect 12360 13376 12449 13379
rect 11664 13354 12449 13376
rect 11664 13348 12388 13354
rect 11664 13336 11670 13348
rect 12437 13345 12449 13354
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12621 13379 12679 13385
rect 12621 13345 12633 13379
rect 12667 13345 12679 13379
rect 12621 13339 12679 13345
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13376 13599 13379
rect 13630 13376 13636 13388
rect 13587 13348 13636 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 6972 13280 7205 13308
rect 6972 13268 6978 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 8662 13268 8668 13320
rect 8720 13268 8726 13320
rect 9876 13308 9904 13336
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 9876 13280 10977 13308
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 4062 13200 4068 13252
rect 4120 13200 4126 13252
rect 12636 13240 12664 13339
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 12820 13308 12848 13339
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 13808 13379 13866 13385
rect 13808 13345 13820 13379
rect 13854 13376 13866 13379
rect 14090 13376 14096 13388
rect 13854 13348 14096 13376
rect 13854 13345 13866 13348
rect 13808 13339 13866 13345
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 14200 13376 14228 13416
rect 15289 13413 15301 13416
rect 15335 13413 15347 13447
rect 19306 13444 19334 13484
rect 24854 13472 24860 13524
rect 24912 13512 24918 13524
rect 25130 13512 25136 13524
rect 24912 13484 25136 13512
rect 24912 13472 24918 13484
rect 25130 13472 25136 13484
rect 25188 13512 25194 13524
rect 25188 13484 26832 13512
rect 25188 13472 25194 13484
rect 20346 13444 20352 13456
rect 15289 13407 15347 13413
rect 16316 13416 16804 13444
rect 19306 13416 20352 13444
rect 16316 13388 16344 13416
rect 15013 13379 15071 13385
rect 15013 13376 15025 13379
rect 14200 13348 15025 13376
rect 15013 13345 15025 13348
rect 15059 13345 15071 13379
rect 15013 13339 15071 13345
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13376 15255 13379
rect 15243 13348 15332 13376
rect 15243 13345 15255 13348
rect 15197 13339 15255 13345
rect 12768 13280 13216 13308
rect 12768 13268 12774 13280
rect 12894 13240 12900 13252
rect 12636 13212 12900 13240
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 3510 13132 3516 13184
rect 3568 13132 3574 13184
rect 4154 13132 4160 13184
rect 4212 13132 4218 13184
rect 4798 13132 4804 13184
rect 4856 13172 4862 13184
rect 5261 13175 5319 13181
rect 5261 13172 5273 13175
rect 4856 13144 5273 13172
rect 4856 13132 4862 13144
rect 5261 13141 5273 13144
rect 5307 13141 5319 13175
rect 5261 13135 5319 13141
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5408 13144 5825 13172
rect 5408 13132 5414 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 5813 13135 5871 13141
rect 6638 13132 6644 13184
rect 6696 13132 6702 13184
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 10594 13172 10600 13184
rect 8619 13144 10600 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10686 13132 10692 13184
rect 10744 13132 10750 13184
rect 12342 13132 12348 13184
rect 12400 13132 12406 13184
rect 12986 13132 12992 13184
rect 13044 13132 13050 13184
rect 13078 13132 13084 13184
rect 13136 13132 13142 13184
rect 13188 13172 13216 13280
rect 15304 13240 15332 13348
rect 15378 13336 15384 13388
rect 15436 13336 15442 13388
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16298 13376 16304 13388
rect 15896 13348 16304 13376
rect 15896 13336 15902 13348
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 16482 13336 16488 13388
rect 16540 13376 16546 13388
rect 16649 13379 16707 13385
rect 16649 13376 16661 13379
rect 16540 13348 16661 13376
rect 16540 13336 16546 13348
rect 16649 13345 16661 13348
rect 16695 13345 16707 13379
rect 16776 13376 16804 13416
rect 20346 13404 20352 13416
rect 20404 13404 20410 13456
rect 20438 13404 20444 13456
rect 20496 13404 20502 13456
rect 23198 13404 23204 13456
rect 23256 13444 23262 13456
rect 23256 13416 26188 13444
rect 23256 13404 23262 13416
rect 18690 13376 18696 13388
rect 16776 13348 18696 13376
rect 16649 13339 16707 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 18782 13336 18788 13388
rect 18840 13336 18846 13388
rect 18966 13336 18972 13388
rect 19024 13336 19030 13388
rect 19061 13379 19119 13385
rect 19061 13345 19073 13379
rect 19107 13345 19119 13379
rect 19061 13339 19119 13345
rect 15562 13268 15568 13320
rect 15620 13268 15626 13320
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 19076 13308 19104 13339
rect 19150 13336 19156 13388
rect 19208 13376 19214 13388
rect 19208 13348 19334 13376
rect 19208 13336 19214 13348
rect 16393 13271 16451 13277
rect 18984 13280 19104 13308
rect 19306 13308 19334 13348
rect 20162 13336 20168 13388
rect 20220 13336 20226 13388
rect 20254 13336 20260 13388
rect 20312 13376 20318 13388
rect 20312 13348 20357 13376
rect 20312 13336 20318 13348
rect 20530 13336 20536 13388
rect 20588 13336 20594 13388
rect 20622 13336 20628 13388
rect 20680 13385 20686 13388
rect 22002 13385 22008 13388
rect 20680 13376 20688 13385
rect 20680 13348 20725 13376
rect 20680 13339 20688 13348
rect 21996 13339 22008 13385
rect 20680 13336 20686 13339
rect 22002 13336 22008 13339
rect 22060 13336 22066 13388
rect 20714 13308 20720 13320
rect 19306 13280 20720 13308
rect 15580 13240 15608 13268
rect 15304 13212 15608 13240
rect 15654 13200 15660 13252
rect 15712 13240 15718 13252
rect 16209 13243 16267 13249
rect 16209 13240 16221 13243
rect 15712 13212 16221 13240
rect 15712 13200 15718 13212
rect 16209 13209 16221 13212
rect 16255 13209 16267 13243
rect 16209 13203 16267 13209
rect 14642 13172 14648 13184
rect 13188 13144 14648 13172
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 14918 13132 14924 13184
rect 14976 13172 14982 13184
rect 15565 13175 15623 13181
rect 15565 13172 15577 13175
rect 14976 13144 15577 13172
rect 14976 13132 14982 13144
rect 15565 13141 15577 13144
rect 15611 13141 15623 13175
rect 16408 13172 16436 13271
rect 17773 13243 17831 13249
rect 17773 13209 17785 13243
rect 17819 13240 17831 13243
rect 18984 13240 19012 13280
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 23216 13317 23244 13404
rect 23474 13385 23480 13388
rect 23468 13339 23480 13385
rect 23474 13336 23480 13339
rect 23532 13336 23538 13388
rect 24872 13385 24900 13416
rect 26160 13388 26188 13416
rect 26234 13404 26240 13456
rect 26292 13444 26298 13456
rect 26697 13447 26755 13453
rect 26697 13444 26709 13447
rect 26292 13416 26709 13444
rect 26292 13404 26298 13416
rect 26697 13413 26709 13416
rect 26743 13413 26755 13447
rect 26697 13407 26755 13413
rect 25130 13385 25136 13388
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13376 24915 13379
rect 25113 13379 25136 13385
rect 24903 13348 24937 13376
rect 24903 13345 24915 13348
rect 24857 13339 24915 13345
rect 25113 13345 25125 13379
rect 25113 13339 25136 13345
rect 25130 13336 25136 13339
rect 25188 13336 25194 13388
rect 26142 13336 26148 13388
rect 26200 13336 26206 13388
rect 26804 13385 26832 13484
rect 26421 13379 26479 13385
rect 26421 13376 26433 13379
rect 26252 13348 26433 13376
rect 21729 13311 21787 13317
rect 21729 13308 21741 13311
rect 21324 13280 21741 13308
rect 21324 13268 21330 13280
rect 21729 13277 21741 13280
rect 21775 13277 21787 13311
rect 21729 13271 21787 13277
rect 23201 13311 23259 13317
rect 23201 13277 23213 13311
rect 23247 13277 23259 13311
rect 23201 13271 23259 13277
rect 21634 13240 21640 13252
rect 17819 13212 19012 13240
rect 19076 13212 21640 13240
rect 17819 13209 17831 13212
rect 17773 13203 17831 13209
rect 17126 13172 17132 13184
rect 16408 13144 17132 13172
rect 15565 13135 15623 13141
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 17310 13132 17316 13184
rect 17368 13172 17374 13184
rect 19076 13172 19104 13212
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 17368 13144 19104 13172
rect 17368 13132 17374 13144
rect 19334 13132 19340 13184
rect 19392 13132 19398 13184
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 20622 13172 20628 13184
rect 19576 13144 20628 13172
rect 19576 13132 19582 13144
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 20806 13132 20812 13184
rect 20864 13132 20870 13184
rect 23106 13132 23112 13184
rect 23164 13132 23170 13184
rect 23216 13172 23244 13271
rect 26252 13249 26280 13348
rect 26421 13345 26433 13348
rect 26467 13345 26479 13379
rect 26421 13339 26479 13345
rect 26605 13379 26663 13385
rect 26605 13345 26617 13379
rect 26651 13345 26663 13379
rect 26605 13339 26663 13345
rect 26789 13379 26847 13385
rect 26789 13345 26801 13379
rect 26835 13345 26847 13379
rect 26789 13339 26847 13345
rect 26237 13243 26295 13249
rect 24504 13212 24854 13240
rect 23382 13172 23388 13184
rect 23216 13144 23388 13172
rect 23382 13132 23388 13144
rect 23440 13132 23446 13184
rect 23934 13132 23940 13184
rect 23992 13172 23998 13184
rect 24504 13172 24532 13212
rect 23992 13144 24532 13172
rect 23992 13132 23998 13144
rect 24578 13132 24584 13184
rect 24636 13132 24642 13184
rect 24826 13172 24854 13212
rect 26237 13209 26249 13243
rect 26283 13209 26295 13243
rect 26237 13203 26295 13209
rect 26620 13240 26648 13339
rect 27798 13240 27804 13252
rect 26620 13212 27804 13240
rect 26620 13172 26648 13212
rect 27798 13200 27804 13212
rect 27856 13200 27862 13252
rect 24826 13144 26648 13172
rect 26878 13132 26884 13184
rect 26936 13172 26942 13184
rect 26973 13175 27031 13181
rect 26973 13172 26985 13175
rect 26936 13144 26985 13172
rect 26936 13132 26942 13144
rect 26973 13141 26985 13144
rect 27019 13141 27031 13175
rect 26973 13135 27031 13141
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 4982 12928 4988 12980
rect 5040 12928 5046 12980
rect 8754 12928 8760 12980
rect 8812 12928 8818 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 12710 12968 12716 12980
rect 11756 12940 12716 12968
rect 11756 12928 11762 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 13078 12928 13084 12980
rect 13136 12928 13142 12980
rect 13998 12928 14004 12980
rect 14056 12968 14062 12980
rect 14093 12971 14151 12977
rect 14093 12968 14105 12971
rect 14056 12940 14105 12968
rect 14056 12928 14062 12940
rect 14093 12937 14105 12940
rect 14139 12968 14151 12971
rect 15657 12971 15715 12977
rect 14139 12940 15608 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 7561 12903 7619 12909
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 11606 12900 11612 12912
rect 7607 12872 11612 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 11606 12860 11612 12872
rect 11664 12860 11670 12912
rect 12437 12903 12495 12909
rect 12437 12900 12449 12903
rect 11716 12872 12449 12900
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 4154 12832 4160 12844
rect 3559 12804 4160 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5552 12804 5825 12832
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 3068 12696 3096 12727
rect 3234 12724 3240 12776
rect 3292 12724 3298 12776
rect 5258 12724 5264 12776
rect 5316 12724 5322 12776
rect 5552 12773 5580 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 11716 12832 11744 12872
rect 12437 12869 12449 12872
rect 12483 12900 12495 12903
rect 12802 12900 12808 12912
rect 12483 12872 12808 12900
rect 12483 12869 12495 12872
rect 12437 12863 12495 12869
rect 12802 12860 12808 12872
rect 12860 12860 12866 12912
rect 12342 12832 12348 12844
rect 5813 12795 5871 12801
rect 8588 12804 11744 12832
rect 11808 12804 12348 12832
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 5994 12764 6000 12776
rect 5767 12736 6000 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 6181 12767 6239 12773
rect 6181 12733 6193 12767
rect 6227 12733 6239 12767
rect 6181 12727 6239 12733
rect 6448 12767 6506 12773
rect 6448 12733 6460 12767
rect 6494 12764 6506 12767
rect 6822 12764 6828 12776
rect 6494 12736 6828 12764
rect 6494 12733 6506 12736
rect 6448 12727 6506 12733
rect 3068 12668 3648 12696
rect 3620 12640 3648 12668
rect 4154 12656 4160 12708
rect 4212 12656 4218 12708
rect 5074 12656 5080 12708
rect 5132 12696 5138 12708
rect 6196 12696 6224 12727
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7650 12724 7656 12776
rect 7708 12724 7714 12776
rect 7742 12724 7748 12776
rect 7800 12764 7806 12776
rect 8588 12773 8616 12804
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 7800 12736 8585 12764
rect 7800 12724 7806 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 9815 12736 9849 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 6914 12696 6920 12708
rect 5132 12668 6920 12696
rect 5132 12656 5138 12668
rect 6914 12656 6920 12668
rect 6972 12696 6978 12708
rect 7466 12696 7472 12708
rect 6972 12668 7472 12696
rect 6972 12656 6978 12668
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 9784 12696 9812 12727
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 11425 12767 11483 12773
rect 11425 12764 11437 12767
rect 10744 12736 11437 12764
rect 10744 12724 10750 12736
rect 11425 12733 11437 12736
rect 11471 12733 11483 12767
rect 11425 12727 11483 12733
rect 11514 12724 11520 12776
rect 11572 12764 11578 12776
rect 11572 12736 11617 12764
rect 11572 12724 11578 12736
rect 11698 12724 11704 12776
rect 11756 12724 11762 12776
rect 11808 12773 11836 12804
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 13096 12832 13124 12928
rect 15580 12900 15608 12940
rect 15657 12937 15669 12971
rect 15703 12968 15715 12971
rect 16482 12968 16488 12980
rect 15703 12940 16488 12968
rect 15703 12937 15715 12940
rect 15657 12931 15715 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 18509 12971 18567 12977
rect 18509 12937 18521 12971
rect 18555 12968 18567 12971
rect 18782 12968 18788 12980
rect 18555 12940 18788 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19392 12940 20668 12968
rect 19392 12928 19398 12940
rect 15838 12900 15844 12912
rect 12820 12804 13124 12832
rect 13188 12872 14964 12900
rect 15580 12872 15844 12900
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 11931 12767 11989 12773
rect 11931 12733 11943 12767
rect 11977 12764 11989 12767
rect 12066 12764 12072 12776
rect 11977 12736 12072 12764
rect 11977 12733 11989 12736
rect 11931 12727 11989 12733
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 12434 12724 12440 12776
rect 12492 12724 12498 12776
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 12820 12773 12848 12804
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 12544 12696 12572 12724
rect 7852 12668 12572 12696
rect 12713 12699 12771 12705
rect 7852 12640 7880 12668
rect 12713 12665 12725 12699
rect 12759 12696 12771 12699
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 12759 12668 12909 12696
rect 12759 12665 12771 12668
rect 12713 12659 12771 12665
rect 12897 12665 12909 12668
rect 12943 12665 12955 12699
rect 13004 12696 13032 12727
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 13188 12764 13216 12872
rect 14936 12832 14964 12872
rect 15838 12860 15844 12872
rect 15896 12860 15902 12912
rect 15933 12903 15991 12909
rect 15933 12869 15945 12903
rect 15979 12900 15991 12903
rect 17034 12900 17040 12912
rect 15979 12872 17040 12900
rect 15979 12869 15991 12872
rect 15933 12863 15991 12869
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 18138 12860 18144 12912
rect 18196 12900 18202 12912
rect 19518 12900 19524 12912
rect 18196 12872 19524 12900
rect 18196 12860 18202 12872
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 13280 12804 14872 12832
rect 14936 12804 15608 12832
rect 13280 12776 13308 12804
rect 13136 12736 13216 12764
rect 13136 12724 13142 12736
rect 13262 12724 13268 12776
rect 13320 12724 13326 12776
rect 13722 12724 13728 12776
rect 13780 12764 13786 12776
rect 14844 12773 14872 12804
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 13780 12736 14565 12764
rect 13780 12724 13786 12736
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12733 14887 12767
rect 14829 12727 14887 12733
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12733 15531 12767
rect 15580 12764 15608 12804
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 16264 12804 17264 12832
rect 16264 12792 16270 12804
rect 15580 12736 16160 12764
rect 15473 12727 15531 12733
rect 13740 12696 13768 12724
rect 13004 12668 13768 12696
rect 13817 12699 13875 12705
rect 12897 12659 12955 12665
rect 13817 12665 13829 12699
rect 13863 12665 13875 12699
rect 13817 12659 13875 12665
rect 3602 12588 3608 12640
rect 3660 12588 3666 12640
rect 5442 12588 5448 12640
rect 5500 12588 5506 12640
rect 5626 12588 5632 12640
rect 5684 12588 5690 12640
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 7098 12628 7104 12640
rect 5960 12600 7104 12628
rect 5960 12588 5966 12600
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 7834 12588 7840 12640
rect 7892 12588 7898 12640
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12628 9643 12631
rect 9674 12628 9680 12640
rect 9631 12600 9680 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 12066 12588 12072 12640
rect 12124 12588 12130 12640
rect 13170 12588 13176 12640
rect 13228 12588 13234 12640
rect 13538 12588 13544 12640
rect 13596 12628 13602 12640
rect 13832 12628 13860 12659
rect 13596 12600 13860 12628
rect 13596 12588 13602 12600
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 14148 12600 14381 12628
rect 14148 12588 14154 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 14642 12588 14648 12640
rect 14700 12588 14706 12640
rect 15488 12628 15516 12727
rect 15838 12656 15844 12708
rect 15896 12696 15902 12708
rect 16025 12699 16083 12705
rect 16025 12696 16037 12699
rect 15896 12668 16037 12696
rect 15896 12656 15902 12668
rect 16025 12665 16037 12668
rect 16071 12665 16083 12699
rect 16132 12696 16160 12736
rect 16298 12724 16304 12776
rect 16356 12724 16362 12776
rect 17126 12724 17132 12776
rect 17184 12724 17190 12776
rect 17236 12764 17264 12804
rect 19352 12804 19748 12832
rect 19352 12773 19380 12804
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 17236 12736 19349 12764
rect 19337 12733 19349 12736
rect 19383 12764 19395 12767
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19383 12736 19437 12764
rect 19536 12736 19625 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 16393 12699 16451 12705
rect 16393 12696 16405 12699
rect 16132 12668 16405 12696
rect 16025 12659 16083 12665
rect 16393 12665 16405 12668
rect 16439 12696 16451 12699
rect 16574 12696 16580 12708
rect 16439 12668 16580 12696
rect 16439 12665 16451 12668
rect 16393 12659 16451 12665
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 16758 12656 16764 12708
rect 16816 12656 16822 12708
rect 16298 12628 16304 12640
rect 15488 12600 16304 12628
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 17144 12628 17172 12724
rect 17396 12699 17454 12705
rect 17396 12665 17408 12699
rect 17442 12696 17454 12699
rect 17862 12696 17868 12708
rect 17442 12668 17868 12696
rect 17442 12665 17454 12668
rect 17396 12659 17454 12665
rect 17862 12656 17868 12668
rect 17920 12656 17926 12708
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 19058 12696 19064 12708
rect 18472 12668 19064 12696
rect 18472 12656 18478 12668
rect 19058 12656 19064 12668
rect 19116 12696 19122 12708
rect 19536 12696 19564 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19720 12764 19748 12804
rect 20640 12764 20668 12940
rect 20806 12928 20812 12980
rect 20864 12928 20870 12980
rect 21913 12971 21971 12977
rect 21913 12937 21925 12971
rect 21959 12968 21971 12971
rect 22002 12968 22008 12980
rect 21959 12940 22008 12968
rect 21959 12937 21971 12940
rect 21913 12931 21971 12937
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 23106 12928 23112 12980
rect 23164 12928 23170 12980
rect 23474 12928 23480 12980
rect 23532 12928 23538 12980
rect 24486 12928 24492 12980
rect 24544 12928 24550 12980
rect 24949 12971 25007 12977
rect 24949 12937 24961 12971
rect 24995 12968 25007 12971
rect 25130 12968 25136 12980
rect 24995 12940 25136 12968
rect 24995 12937 25007 12940
rect 24949 12931 25007 12937
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 20824 12832 20852 12928
rect 20993 12903 21051 12909
rect 20993 12869 21005 12903
rect 21039 12900 21051 12903
rect 21039 12872 21312 12900
rect 21039 12869 21051 12872
rect 20993 12863 21051 12869
rect 20824 12804 21220 12832
rect 21192 12773 21220 12804
rect 21085 12767 21143 12773
rect 21085 12764 21097 12767
rect 19720 12736 20301 12764
rect 20640 12736 21097 12764
rect 19613 12727 19671 12733
rect 19116 12668 19564 12696
rect 19858 12699 19916 12705
rect 19116 12656 19122 12668
rect 19858 12665 19870 12699
rect 19904 12665 19916 12699
rect 19858 12659 19916 12665
rect 18432 12628 18460 12656
rect 17144 12600 18460 12628
rect 19521 12631 19579 12637
rect 19521 12597 19533 12631
rect 19567 12628 19579 12631
rect 19873 12628 19901 12659
rect 19567 12600 19901 12628
rect 20273 12628 20301 12736
rect 21085 12733 21097 12736
rect 21131 12733 21143 12767
rect 21085 12727 21143 12733
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12733 21235 12767
rect 21284 12764 21312 12872
rect 21634 12860 21640 12912
rect 21692 12900 21698 12912
rect 22922 12900 22928 12912
rect 21692 12872 22928 12900
rect 21692 12860 21698 12872
rect 22922 12860 22928 12872
rect 22980 12860 22986 12912
rect 23014 12832 23020 12844
rect 21560 12804 21864 12832
rect 21361 12767 21419 12773
rect 21361 12764 21373 12767
rect 21284 12736 21373 12764
rect 21177 12727 21235 12733
rect 21361 12733 21373 12736
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 21453 12767 21511 12773
rect 21453 12733 21465 12767
rect 21499 12733 21511 12767
rect 21453 12727 21511 12733
rect 20990 12656 20996 12708
rect 21048 12696 21054 12708
rect 21468 12696 21496 12727
rect 21048 12668 21496 12696
rect 21048 12656 21054 12668
rect 21560 12628 21588 12804
rect 21726 12724 21732 12776
rect 21784 12724 21790 12776
rect 21836 12764 21864 12804
rect 22480 12804 23020 12832
rect 22480 12773 22508 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 23124 12832 23152 12928
rect 23201 12903 23259 12909
rect 23201 12869 23213 12903
rect 23247 12900 23259 12903
rect 23842 12900 23848 12912
rect 23247 12872 23848 12900
rect 23247 12869 23259 12872
rect 23201 12863 23259 12869
rect 23842 12860 23848 12872
rect 23900 12860 23906 12912
rect 24578 12832 24584 12844
rect 23124 12804 23980 12832
rect 22281 12767 22339 12773
rect 22281 12764 22293 12767
rect 21836 12736 22293 12764
rect 22281 12733 22293 12736
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 22465 12767 22523 12773
rect 22465 12733 22477 12767
rect 22511 12733 22523 12767
rect 22465 12727 22523 12733
rect 23032 12736 23250 12764
rect 21637 12699 21695 12705
rect 21637 12665 21649 12699
rect 21683 12696 21695 12699
rect 23032 12696 23060 12736
rect 21683 12668 23060 12696
rect 23222 12696 23250 12736
rect 23290 12724 23296 12776
rect 23348 12724 23354 12776
rect 23952 12773 23980 12804
rect 24228 12804 24584 12832
rect 24228 12773 24256 12804
rect 24578 12792 24584 12804
rect 24636 12792 24642 12844
rect 25976 12804 27384 12832
rect 25976 12776 26004 12804
rect 23937 12767 23995 12773
rect 23937 12733 23949 12767
rect 23983 12733 23995 12767
rect 23937 12727 23995 12733
rect 24213 12767 24271 12773
rect 24213 12733 24225 12767
rect 24259 12733 24271 12767
rect 24213 12727 24271 12733
rect 24302 12724 24308 12776
rect 24360 12724 24366 12776
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 25958 12724 25964 12776
rect 26016 12724 26022 12776
rect 26878 12724 26884 12776
rect 26936 12724 26942 12776
rect 27062 12773 27068 12776
rect 27029 12767 27068 12773
rect 27029 12733 27041 12767
rect 27029 12727 27068 12733
rect 27062 12724 27068 12727
rect 27120 12724 27126 12776
rect 27356 12773 27384 12804
rect 27346 12767 27404 12773
rect 27346 12733 27358 12767
rect 27392 12733 27404 12767
rect 27346 12727 27404 12733
rect 23222 12668 23980 12696
rect 21683 12665 21695 12668
rect 21637 12659 21695 12665
rect 20273 12600 21588 12628
rect 19567 12597 19579 12600
rect 19521 12591 19579 12597
rect 22370 12588 22376 12640
rect 22428 12588 22434 12640
rect 23952 12628 23980 12668
rect 24026 12656 24032 12708
rect 24084 12696 24090 12708
rect 24121 12699 24179 12705
rect 24121 12696 24133 12699
rect 24084 12668 24133 12696
rect 24084 12656 24090 12668
rect 24121 12665 24133 12668
rect 24167 12665 24179 12699
rect 24320 12696 24348 12724
rect 26418 12696 26424 12708
rect 24320 12668 26424 12696
rect 24121 12659 24179 12665
rect 26418 12656 26424 12668
rect 26476 12696 26482 12708
rect 27157 12699 27215 12705
rect 27157 12696 27169 12699
rect 26476 12668 27169 12696
rect 26476 12656 26482 12668
rect 27157 12665 27169 12668
rect 27203 12665 27215 12699
rect 27157 12659 27215 12665
rect 27246 12656 27252 12708
rect 27304 12656 27310 12708
rect 24854 12628 24860 12640
rect 23952 12600 24860 12628
rect 24854 12588 24860 12600
rect 24912 12588 24918 12640
rect 26234 12588 26240 12640
rect 26292 12628 26298 12640
rect 27525 12631 27583 12637
rect 27525 12628 27537 12631
rect 26292 12600 27537 12628
rect 26292 12588 26298 12600
rect 27525 12597 27537 12600
rect 27571 12597 27583 12631
rect 27525 12591 27583 12597
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4154 12424 4160 12436
rect 4019 12396 4160 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 4893 12427 4951 12433
rect 4893 12424 4905 12427
rect 4672 12396 4905 12424
rect 4672 12384 4678 12396
rect 4893 12393 4905 12396
rect 4939 12424 4951 12427
rect 5166 12424 5172 12436
rect 4939 12396 5172 12424
rect 4939 12393 4951 12396
rect 4893 12387 4951 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5718 12424 5724 12436
rect 5316 12396 5724 12424
rect 5316 12384 5322 12396
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 6822 12384 6828 12436
rect 6880 12384 6886 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 6972 12396 7297 12424
rect 6972 12384 6978 12396
rect 7285 12393 7297 12396
rect 7331 12393 7343 12427
rect 7285 12387 7343 12393
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 11149 12427 11207 12433
rect 7524 12396 7972 12424
rect 7524 12384 7530 12396
rect 3510 12316 3516 12368
rect 3568 12356 3574 12368
rect 3697 12359 3755 12365
rect 3697 12356 3709 12359
rect 3568 12328 3709 12356
rect 3568 12316 3574 12328
rect 3697 12325 3709 12328
rect 3743 12325 3755 12359
rect 3697 12319 3755 12325
rect 5000 12328 5396 12356
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12257 3939 12291
rect 3881 12251 3939 12257
rect 3896 12220 3924 12251
rect 4614 12248 4620 12300
rect 4672 12297 4678 12300
rect 4672 12288 4681 12297
rect 4672 12260 4717 12288
rect 4672 12251 4681 12260
rect 4672 12248 4678 12251
rect 4798 12248 4804 12300
rect 4856 12248 4862 12300
rect 4890 12248 4896 12300
rect 4948 12248 4954 12300
rect 5000 12297 5028 12328
rect 5368 12300 5396 12328
rect 5534 12316 5540 12368
rect 5592 12316 5598 12368
rect 6840 12356 6868 12384
rect 7193 12359 7251 12365
rect 6380 12328 6684 12356
rect 6840 12328 7144 12356
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12257 5043 12291
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 4985 12251 5043 12257
rect 5092 12260 5273 12288
rect 4062 12220 4068 12232
rect 3896 12192 4068 12220
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3896 12084 3924 12192
rect 4062 12180 4068 12192
rect 4120 12220 4126 12232
rect 4908 12220 4936 12248
rect 5092 12220 5120 12260
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 4120 12192 5120 12220
rect 4120 12180 4126 12192
rect 5166 12180 5172 12232
rect 5224 12180 5230 12232
rect 5276 12220 5304 12251
rect 5350 12248 5356 12300
rect 5408 12248 5414 12300
rect 5810 12288 5816 12300
rect 5781 12278 5816 12288
rect 5736 12250 5816 12278
rect 5736 12220 5764 12250
rect 5810 12248 5816 12250
rect 5868 12248 5874 12300
rect 5994 12248 6000 12300
rect 6052 12248 6058 12300
rect 6380 12297 6408 12328
rect 6656 12300 6684 12328
rect 6365 12291 6423 12297
rect 6365 12257 6377 12291
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6546 12248 6552 12300
rect 6604 12248 6610 12300
rect 6638 12248 6644 12300
rect 6696 12248 6702 12300
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 7006 12288 7012 12300
rect 6963 12260 7012 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 5813 12247 5825 12248
rect 5859 12247 5871 12248
rect 5813 12241 5871 12247
rect 5276 12192 5764 12220
rect 4798 12112 4804 12164
rect 4856 12112 4862 12164
rect 5258 12112 5264 12164
rect 5316 12152 5322 12164
rect 5353 12155 5411 12161
rect 5353 12152 5365 12155
rect 5316 12124 5365 12152
rect 5316 12112 5322 12124
rect 5353 12121 5365 12124
rect 5399 12152 5411 12155
rect 5399 12124 5764 12152
rect 5399 12121 5411 12124
rect 5353 12115 5411 12121
rect 3660 12056 3924 12084
rect 5736 12084 5764 12124
rect 5810 12112 5816 12164
rect 5868 12152 5874 12164
rect 5905 12155 5963 12161
rect 5905 12152 5917 12155
rect 5868 12124 5917 12152
rect 5868 12112 5874 12124
rect 5905 12121 5917 12124
rect 5951 12121 5963 12155
rect 6012 12152 6040 12248
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 6144 12192 6469 12220
rect 6144 12180 6150 12192
rect 6457 12189 6469 12192
rect 6503 12220 6515 12223
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6503 12192 6745 12220
rect 6503 12189 6515 12192
rect 6457 12183 6515 12189
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 6840 12220 6868 12251
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7116 12288 7144 12328
rect 7193 12325 7205 12359
rect 7239 12356 7251 12359
rect 7745 12359 7803 12365
rect 7745 12356 7757 12359
rect 7239 12328 7757 12356
rect 7239 12325 7251 12328
rect 7193 12319 7251 12325
rect 7745 12325 7757 12328
rect 7791 12325 7803 12359
rect 7745 12319 7803 12325
rect 7282 12288 7288 12300
rect 7116 12260 7288 12288
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 7653 12291 7711 12297
rect 7653 12288 7665 12291
rect 7484 12260 7665 12288
rect 7484 12220 7512 12260
rect 7653 12257 7665 12260
rect 7699 12257 7711 12291
rect 7653 12251 7711 12257
rect 6840 12192 7512 12220
rect 6733 12183 6791 12189
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7668 12220 7696 12251
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 7944 12297 7972 12396
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11238 12424 11244 12436
rect 11195 12396 11244 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 12584 12396 12725 12424
rect 12584 12384 12590 12396
rect 12713 12393 12725 12396
rect 12759 12393 12771 12427
rect 12713 12387 12771 12393
rect 13262 12384 13268 12436
rect 13320 12384 13326 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13372 12396 13645 12424
rect 9674 12365 9680 12368
rect 9668 12356 9680 12365
rect 9635 12328 9680 12356
rect 9668 12319 9680 12328
rect 9674 12316 9680 12319
rect 9732 12316 9738 12368
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 11514 12356 11520 12368
rect 9916 12328 11520 12356
rect 9916 12316 9922 12328
rect 11514 12316 11520 12328
rect 11572 12316 11578 12368
rect 12066 12356 12072 12368
rect 11624 12328 12072 12356
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8018 12248 8024 12300
rect 8076 12248 8082 12300
rect 8196 12291 8254 12297
rect 8196 12257 8208 12291
rect 8242 12288 8254 12291
rect 8662 12288 8668 12300
rect 8242 12260 8668 12288
rect 8242 12257 8254 12260
rect 8196 12251 8254 12257
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 9401 12291 9459 12297
rect 9401 12257 9413 12291
rect 9447 12288 9459 12291
rect 9876 12288 9904 12316
rect 11624 12297 11652 12328
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 12618 12316 12624 12368
rect 12676 12316 12682 12368
rect 12989 12359 13047 12365
rect 12989 12325 13001 12359
rect 13035 12356 13047 12359
rect 13170 12356 13176 12368
rect 13035 12328 13176 12356
rect 13035 12325 13047 12328
rect 12989 12319 13047 12325
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 9447 12260 9904 12288
rect 10704 12260 10977 12288
rect 9447 12257 9459 12260
rect 9401 12251 9459 12257
rect 8036 12220 8064 12248
rect 7668 12192 8064 12220
rect 6914 12152 6920 12164
rect 6012 12124 6920 12152
rect 5905 12115 5963 12121
rect 6914 12112 6920 12124
rect 6972 12152 6978 12164
rect 7009 12155 7067 12161
rect 7009 12152 7021 12155
rect 6972 12124 7021 12152
rect 6972 12112 6978 12124
rect 7009 12121 7021 12124
rect 7055 12121 7067 12155
rect 7377 12155 7435 12161
rect 7377 12152 7389 12155
rect 7009 12115 7067 12121
rect 7116 12124 7389 12152
rect 5997 12087 6055 12093
rect 5997 12084 6009 12087
rect 5736 12056 6009 12084
rect 3660 12044 3666 12056
rect 5997 12053 6009 12056
rect 6043 12053 6055 12087
rect 5997 12047 6055 12053
rect 6638 12044 6644 12096
rect 6696 12084 6702 12096
rect 7116 12093 7144 12124
rect 7377 12121 7389 12124
rect 7423 12121 7435 12155
rect 7377 12115 7435 12121
rect 10704 12096 10732 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 12713 12291 12771 12297
rect 12713 12288 12725 12291
rect 12452 12260 12725 12288
rect 11698 12180 11704 12232
rect 11756 12220 11762 12232
rect 12069 12223 12127 12229
rect 12069 12220 12081 12223
rect 11756 12192 12081 12220
rect 11756 12180 11762 12192
rect 12069 12189 12081 12192
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 12452 12164 12480 12260
rect 12713 12257 12725 12260
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 12802 12248 12808 12300
rect 12860 12248 12866 12300
rect 13372 12297 13400 12396
rect 13633 12393 13645 12396
rect 13679 12424 13691 12427
rect 13722 12424 13728 12436
rect 13679 12396 13728 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 13998 12384 14004 12436
rect 14056 12384 14062 12436
rect 16206 12384 16212 12436
rect 16264 12384 16270 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16356 12396 16896 12424
rect 16356 12384 16362 12396
rect 14016 12356 14044 12384
rect 13648 12328 14044 12356
rect 14360 12359 14418 12365
rect 13648 12297 13676 12328
rect 14360 12325 14372 12359
rect 14406 12356 14418 12359
rect 14642 12356 14648 12368
rect 14406 12328 14648 12356
rect 14406 12325 14418 12328
rect 14360 12319 14418 12325
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 14826 12316 14832 12368
rect 14884 12356 14890 12368
rect 14884 12328 15700 12356
rect 14884 12316 14890 12328
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13633 12291 13691 12297
rect 13633 12288 13645 12291
rect 13357 12251 13415 12257
rect 13464 12260 13645 12288
rect 13280 12220 13308 12251
rect 13464 12220 13492 12260
rect 13633 12257 13645 12260
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 13909 12291 13967 12297
rect 13909 12257 13921 12291
rect 13955 12288 13967 12291
rect 13955 12260 15240 12288
rect 13955 12257 13967 12260
rect 13909 12251 13967 12257
rect 13280 12192 13492 12220
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12189 14151 12223
rect 15212 12220 15240 12260
rect 15212 12192 15608 12220
rect 14093 12183 14151 12189
rect 12434 12112 12440 12164
rect 12492 12112 12498 12164
rect 12802 12112 12808 12164
rect 12860 12152 12866 12164
rect 13078 12152 13084 12164
rect 12860 12124 13084 12152
rect 12860 12112 12866 12124
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 13262 12112 13268 12164
rect 13320 12152 13326 12164
rect 13725 12155 13783 12161
rect 13725 12152 13737 12155
rect 13320 12124 13737 12152
rect 13320 12112 13326 12124
rect 13725 12121 13737 12124
rect 13771 12121 13783 12155
rect 13725 12115 13783 12121
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 6696 12056 7113 12084
rect 6696 12044 6702 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7101 12047 7159 12053
rect 9309 12087 9367 12093
rect 9309 12053 9321 12087
rect 9355 12084 9367 12087
rect 9582 12084 9588 12096
rect 9355 12056 9588 12084
rect 9355 12053 9367 12056
rect 9309 12047 9367 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10686 12084 10692 12096
rect 9732 12056 10692 12084
rect 9732 12044 9738 12056
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 10778 12044 10784 12096
rect 10836 12044 10842 12096
rect 11514 12044 11520 12096
rect 11572 12084 11578 12096
rect 14108 12084 14136 12183
rect 11572 12056 14136 12084
rect 11572 12044 11578 12056
rect 15470 12044 15476 12096
rect 15528 12044 15534 12096
rect 15580 12084 15608 12192
rect 15672 12152 15700 12328
rect 15948 12328 16804 12356
rect 15838 12248 15844 12300
rect 15896 12288 15902 12300
rect 15948 12297 15976 12328
rect 15933 12291 15991 12297
rect 15933 12288 15945 12291
rect 15896 12260 15945 12288
rect 15896 12248 15902 12260
rect 15933 12257 15945 12260
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 16209 12291 16267 12297
rect 16209 12257 16221 12291
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 16224 12220 16252 12251
rect 16298 12248 16304 12300
rect 16356 12248 16362 12300
rect 16390 12248 16396 12300
rect 16448 12248 16454 12300
rect 16574 12248 16580 12300
rect 16632 12248 16638 12300
rect 16776 12297 16804 12328
rect 16868 12297 16896 12396
rect 17862 12384 17868 12436
rect 17920 12384 17926 12436
rect 19429 12427 19487 12433
rect 19429 12393 19441 12427
rect 19475 12424 19487 12427
rect 23109 12427 23167 12433
rect 19475 12396 22232 12424
rect 19475 12393 19487 12396
rect 19429 12387 19487 12393
rect 18233 12359 18291 12365
rect 18233 12325 18245 12359
rect 18279 12356 18291 12359
rect 18877 12359 18935 12365
rect 18877 12356 18889 12359
rect 18279 12328 18889 12356
rect 18279 12325 18291 12328
rect 18233 12319 18291 12325
rect 18877 12325 18889 12328
rect 18923 12325 18935 12359
rect 18877 12319 18935 12325
rect 19168 12328 19472 12356
rect 16761 12291 16819 12297
rect 16761 12257 16773 12291
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 16853 12291 16911 12297
rect 16853 12257 16865 12291
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 17034 12248 17040 12300
rect 17092 12248 17098 12300
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12288 17555 12291
rect 18049 12291 18107 12297
rect 18049 12288 18061 12291
rect 17543 12260 17816 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 16408 12220 16436 12248
rect 16224 12192 16436 12220
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12220 16543 12223
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 16531 12192 16681 12220
rect 16531 12189 16543 12192
rect 16485 12183 16543 12189
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 17328 12220 17356 12251
rect 17589 12223 17647 12229
rect 17589 12220 17601 12223
rect 17328 12192 17601 12220
rect 16669 12183 16727 12189
rect 17589 12189 17601 12192
rect 17635 12189 17647 12223
rect 17589 12183 17647 12189
rect 15749 12155 15807 12161
rect 15749 12152 15761 12155
rect 15672 12124 15761 12152
rect 15749 12121 15761 12124
rect 15795 12121 15807 12155
rect 17313 12155 17371 12161
rect 17313 12152 17325 12155
rect 15749 12115 15807 12121
rect 15856 12124 17325 12152
rect 15856 12084 15884 12124
rect 17313 12121 17325 12124
rect 17359 12121 17371 12155
rect 17788 12152 17816 12260
rect 17880 12260 18061 12288
rect 17880 12232 17908 12260
rect 18049 12257 18061 12260
rect 18095 12288 18107 12291
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 18095 12260 18153 12288
rect 18095 12257 18107 12260
rect 18049 12251 18107 12257
rect 18141 12257 18153 12260
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 18325 12291 18383 12297
rect 18325 12257 18337 12291
rect 18371 12288 18383 12291
rect 18690 12288 18696 12300
rect 18371 12260 18696 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 19168 12297 19196 12328
rect 19444 12300 19472 12328
rect 19720 12328 20484 12356
rect 18785 12291 18843 12297
rect 18785 12257 18797 12291
rect 18831 12288 18843 12291
rect 19153 12291 19211 12297
rect 19153 12288 19165 12291
rect 18831 12260 19165 12288
rect 18831 12257 18843 12260
rect 18785 12251 18843 12257
rect 19153 12257 19165 12260
rect 19199 12257 19211 12291
rect 19153 12251 19211 12257
rect 19245 12291 19303 12297
rect 19245 12257 19257 12291
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 17862 12180 17868 12232
rect 17920 12180 17926 12232
rect 18506 12180 18512 12232
rect 18564 12180 18570 12232
rect 18874 12220 18880 12232
rect 18616 12192 18880 12220
rect 17954 12152 17960 12164
rect 17788 12124 17960 12152
rect 17313 12115 17371 12121
rect 17954 12112 17960 12124
rect 18012 12112 18018 12164
rect 15580 12056 15884 12084
rect 17037 12087 17095 12093
rect 17037 12053 17049 12087
rect 17083 12084 17095 12087
rect 18616 12084 18644 12192
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 19260 12220 19288 12251
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19720 12297 19748 12328
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19484 12260 19717 12288
rect 19484 12248 19490 12260
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12288 19855 12291
rect 20070 12288 20076 12300
rect 19843 12260 20076 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 20254 12248 20260 12300
rect 20312 12288 20318 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 20312 12260 20361 12288
rect 20312 12248 20318 12260
rect 20349 12257 20361 12260
rect 20395 12257 20407 12291
rect 20349 12251 20407 12257
rect 19886 12220 19892 12232
rect 19076 12192 19288 12220
rect 19352 12192 19892 12220
rect 19076 12161 19104 12192
rect 18693 12155 18751 12161
rect 18693 12121 18705 12155
rect 18739 12121 18751 12155
rect 18693 12115 18751 12121
rect 18785 12155 18843 12161
rect 18785 12121 18797 12155
rect 18831 12152 18843 12155
rect 19061 12155 19119 12161
rect 19061 12152 19073 12155
rect 18831 12124 19073 12152
rect 18831 12121 18843 12124
rect 18785 12115 18843 12121
rect 19061 12121 19073 12124
rect 19107 12121 19119 12155
rect 19061 12115 19119 12121
rect 19153 12155 19211 12161
rect 19153 12121 19165 12155
rect 19199 12152 19211 12155
rect 19352 12152 19380 12192
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12220 20039 12223
rect 20027 12192 20392 12220
rect 20027 12189 20039 12192
rect 19981 12183 20039 12189
rect 20364 12161 20392 12192
rect 20349 12155 20407 12161
rect 19199 12124 19380 12152
rect 19444 12124 20300 12152
rect 19199 12121 19211 12124
rect 19153 12115 19211 12121
rect 17083 12056 18644 12084
rect 18708 12084 18736 12115
rect 19168 12084 19196 12115
rect 18708 12056 19196 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19444 12084 19472 12124
rect 20272 12096 20300 12124
rect 20349 12121 20361 12155
rect 20395 12121 20407 12155
rect 20456 12152 20484 12328
rect 20824 12328 21777 12356
rect 20533 12291 20591 12297
rect 20533 12257 20545 12291
rect 20579 12288 20591 12291
rect 20824 12288 20852 12328
rect 21749 12300 21777 12328
rect 21836 12328 22140 12356
rect 20579 12260 20852 12288
rect 20579 12257 20591 12260
rect 20533 12251 20591 12257
rect 20898 12248 20904 12300
rect 20956 12248 20962 12300
rect 21082 12248 21088 12300
rect 21140 12248 21146 12300
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 21453 12291 21511 12297
rect 21453 12288 21465 12291
rect 21416 12260 21465 12288
rect 21416 12248 21422 12260
rect 21453 12257 21465 12260
rect 21499 12257 21511 12291
rect 21453 12251 21511 12257
rect 21545 12291 21603 12297
rect 21545 12257 21557 12291
rect 21591 12257 21603 12291
rect 21545 12251 21603 12257
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12220 21051 12223
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21039 12192 21281 12220
rect 21039 12189 21051 12192
rect 20993 12183 21051 12189
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21560 12220 21588 12251
rect 21634 12248 21640 12300
rect 21692 12248 21698 12300
rect 21726 12248 21732 12300
rect 21784 12248 21790 12300
rect 21269 12183 21327 12189
rect 21468 12192 21588 12220
rect 21468 12164 21496 12192
rect 21450 12152 21456 12164
rect 20456 12124 21456 12152
rect 20349 12115 20407 12121
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 21749 12161 21777 12248
rect 21836 12232 21864 12328
rect 22002 12248 22008 12300
rect 22060 12248 22066 12300
rect 21818 12180 21824 12232
rect 21876 12180 21882 12232
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22112 12220 22140 12328
rect 22204 12297 22232 12396
rect 23109 12393 23121 12427
rect 23155 12424 23167 12427
rect 25225 12427 25283 12433
rect 23155 12396 24992 12424
rect 23155 12393 23167 12396
rect 23109 12387 23167 12393
rect 22370 12316 22376 12368
rect 22428 12356 22434 12368
rect 22465 12359 22523 12365
rect 22465 12356 22477 12359
rect 22428 12328 22477 12356
rect 22428 12316 22434 12328
rect 22465 12325 22477 12328
rect 22511 12325 22523 12359
rect 23124 12356 23152 12387
rect 23842 12356 23848 12368
rect 22465 12319 22523 12325
rect 22664 12328 23152 12356
rect 23492 12328 23848 12356
rect 22189 12291 22247 12297
rect 22189 12257 22201 12291
rect 22235 12288 22247 12291
rect 22554 12288 22560 12300
rect 22235 12260 22560 12288
rect 22235 12257 22247 12260
rect 22189 12251 22247 12257
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 22664 12297 22692 12328
rect 22649 12291 22707 12297
rect 22649 12257 22661 12291
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 22738 12248 22744 12300
rect 22796 12248 22802 12300
rect 23014 12248 23020 12300
rect 23072 12288 23078 12300
rect 23072 12287 23152 12288
rect 23072 12281 23167 12287
rect 23072 12260 23121 12281
rect 23072 12248 23078 12260
rect 23109 12247 23121 12260
rect 23155 12247 23167 12281
rect 23198 12248 23204 12300
rect 23256 12248 23262 12300
rect 23492 12297 23520 12328
rect 23842 12316 23848 12328
rect 23900 12316 23906 12368
rect 23385 12291 23443 12297
rect 23385 12257 23397 12291
rect 23431 12257 23443 12291
rect 23385 12251 23443 12257
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 23109 12241 23167 12247
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 21959 12192 22048 12220
rect 22112 12192 22845 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 22020 12161 22048 12192
rect 22833 12189 22845 12192
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 23400 12220 23428 12251
rect 23566 12248 23572 12300
rect 23624 12248 23630 12300
rect 23661 12291 23719 12297
rect 23661 12257 23673 12291
rect 23707 12288 23719 12291
rect 23952 12288 23980 12396
rect 24118 12297 24124 12300
rect 23707 12260 23980 12288
rect 23707 12257 23719 12260
rect 23661 12251 23719 12257
rect 24112 12251 24124 12297
rect 24118 12248 24124 12251
rect 24176 12248 24182 12300
rect 23584 12220 23612 12248
rect 23400 12192 23612 12220
rect 21545 12155 21603 12161
rect 21545 12121 21557 12155
rect 21591 12152 21603 12155
rect 21729 12155 21787 12161
rect 21729 12152 21741 12155
rect 21591 12124 21741 12152
rect 21591 12121 21603 12124
rect 21545 12115 21603 12121
rect 21729 12121 21741 12124
rect 21775 12121 21787 12155
rect 21729 12115 21787 12121
rect 22005 12155 22063 12161
rect 22005 12121 22017 12155
rect 22051 12121 22063 12155
rect 22005 12115 22063 12121
rect 22741 12155 22799 12161
rect 22741 12121 22753 12155
rect 22787 12152 22799 12155
rect 23017 12155 23075 12161
rect 23017 12152 23029 12155
rect 22787 12124 23029 12152
rect 22787 12121 22799 12124
rect 22741 12115 22799 12121
rect 23017 12121 23029 12124
rect 23063 12152 23075 12155
rect 23400 12152 23428 12192
rect 23842 12180 23848 12232
rect 23900 12180 23906 12232
rect 24964 12220 24992 12396
rect 25225 12393 25237 12427
rect 25271 12424 25283 12427
rect 26237 12427 26295 12433
rect 25271 12396 25728 12424
rect 25271 12393 25283 12396
rect 25225 12387 25283 12393
rect 25038 12316 25044 12368
rect 25096 12356 25102 12368
rect 25700 12365 25728 12396
rect 26237 12393 26249 12427
rect 26283 12393 26295 12427
rect 26237 12387 26295 12393
rect 25593 12359 25651 12365
rect 25593 12356 25605 12359
rect 25096 12328 25605 12356
rect 25096 12316 25102 12328
rect 25593 12325 25605 12328
rect 25639 12325 25651 12359
rect 25593 12319 25651 12325
rect 25685 12359 25743 12365
rect 25685 12325 25697 12359
rect 25731 12325 25743 12359
rect 26252 12356 26280 12387
rect 27246 12384 27252 12436
rect 27304 12424 27310 12436
rect 27893 12427 27951 12433
rect 27893 12424 27905 12427
rect 27304 12396 27905 12424
rect 27304 12384 27310 12396
rect 27893 12393 27905 12396
rect 27939 12393 27951 12427
rect 27893 12387 27951 12393
rect 26666 12359 26724 12365
rect 26666 12356 26678 12359
rect 26252 12328 26678 12356
rect 25685 12319 25743 12325
rect 26666 12325 26678 12328
rect 26712 12325 26724 12359
rect 26666 12319 26724 12325
rect 25222 12248 25228 12300
rect 25280 12288 25286 12300
rect 25317 12291 25375 12297
rect 25317 12288 25329 12291
rect 25280 12260 25329 12288
rect 25280 12248 25286 12260
rect 25317 12257 25329 12260
rect 25363 12257 25375 12291
rect 25317 12251 25375 12257
rect 25410 12291 25468 12297
rect 25410 12257 25422 12291
rect 25456 12288 25468 12291
rect 25498 12288 25504 12300
rect 25456 12260 25504 12288
rect 25456 12257 25468 12260
rect 25410 12251 25468 12257
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 25774 12248 25780 12300
rect 25832 12297 25838 12300
rect 25832 12251 25840 12297
rect 26053 12291 26111 12297
rect 26053 12257 26065 12291
rect 26099 12257 26111 12291
rect 26053 12251 26111 12257
rect 25832 12248 25838 12251
rect 26068 12220 26096 12251
rect 26142 12248 26148 12300
rect 26200 12288 26206 12300
rect 26421 12291 26479 12297
rect 26421 12288 26433 12291
rect 26200 12260 26433 12288
rect 26200 12248 26206 12260
rect 26421 12257 26433 12260
rect 26467 12257 26479 12291
rect 26421 12251 26479 12257
rect 27706 12248 27712 12300
rect 27764 12288 27770 12300
rect 29006 12291 29064 12297
rect 29006 12288 29018 12291
rect 27764 12260 29018 12288
rect 27764 12248 27770 12260
rect 29006 12257 29018 12260
rect 29052 12257 29064 12291
rect 29006 12251 29064 12257
rect 24964 12192 26096 12220
rect 29270 12180 29276 12232
rect 29328 12180 29334 12232
rect 23063 12124 23428 12152
rect 23063 12121 23075 12124
rect 23017 12115 23075 12121
rect 19300 12056 19472 12084
rect 19300 12044 19306 12056
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19576 12056 19717 12084
rect 19576 12044 19582 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 20254 12044 20260 12096
rect 20312 12044 20318 12096
rect 20622 12044 20628 12096
rect 20680 12044 20686 12096
rect 21266 12044 21272 12096
rect 21324 12084 21330 12096
rect 21821 12087 21879 12093
rect 21821 12084 21833 12087
rect 21324 12056 21833 12084
rect 21324 12044 21330 12056
rect 21821 12053 21833 12056
rect 21867 12084 21879 12087
rect 22830 12084 22836 12096
rect 21867 12056 22836 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 23198 12044 23204 12096
rect 23256 12044 23262 12096
rect 23474 12044 23480 12096
rect 23532 12044 23538 12096
rect 25961 12087 26019 12093
rect 25961 12053 25973 12087
rect 26007 12084 26019 12087
rect 26326 12084 26332 12096
rect 26007 12056 26332 12084
rect 26007 12053 26019 12056
rect 25961 12047 26019 12053
rect 26326 12044 26332 12056
rect 26384 12044 26390 12096
rect 27062 12044 27068 12096
rect 27120 12084 27126 12096
rect 27801 12087 27859 12093
rect 27801 12084 27813 12087
rect 27120 12056 27813 12084
rect 27120 12044 27126 12056
rect 27801 12053 27813 12056
rect 27847 12053 27859 12087
rect 27801 12047 27859 12053
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 6086 11880 6092 11892
rect 5224 11852 6092 11880
rect 5224 11840 5230 11852
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7653 11883 7711 11889
rect 7653 11880 7665 11883
rect 7616 11852 7665 11880
rect 7616 11840 7622 11852
rect 7653 11849 7665 11852
rect 7699 11849 7711 11883
rect 7653 11843 7711 11849
rect 8662 11840 8668 11892
rect 8720 11840 8726 11892
rect 11701 11883 11759 11889
rect 11701 11849 11713 11883
rect 11747 11880 11759 11883
rect 11790 11880 11796 11892
rect 11747 11852 11796 11880
rect 11747 11849 11759 11852
rect 11701 11843 11759 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 12710 11880 12716 11892
rect 11940 11852 12716 11880
rect 11940 11840 11946 11852
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 18230 11880 18236 11892
rect 15320 11852 18236 11880
rect 4706 11812 4712 11824
rect 3528 11784 4712 11812
rect 3528 11753 3556 11784
rect 4706 11772 4712 11784
rect 4764 11772 4770 11824
rect 6638 11772 6644 11824
rect 6696 11772 6702 11824
rect 7742 11812 7748 11824
rect 7484 11784 7748 11812
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3786 11704 3792 11756
rect 3844 11704 3850 11756
rect 4614 11704 4620 11756
rect 4672 11704 4678 11756
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3467 11648 3556 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3528 11552 3556 11648
rect 4062 11636 4068 11688
rect 4120 11636 4126 11688
rect 4632 11661 4660 11704
rect 4893 11679 4951 11685
rect 4617 11655 4675 11661
rect 4617 11621 4629 11655
rect 4663 11621 4675 11655
rect 4893 11645 4905 11679
rect 4939 11676 4951 11679
rect 6656 11676 6684 11772
rect 7484 11685 7512 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 7929 11815 7987 11821
rect 7929 11781 7941 11815
rect 7975 11812 7987 11815
rect 8570 11812 8576 11824
rect 7975 11784 8576 11812
rect 7975 11781 7987 11784
rect 7929 11775 7987 11781
rect 8570 11772 8576 11784
rect 8628 11772 8634 11824
rect 9214 11772 9220 11824
rect 9272 11812 9278 11824
rect 11054 11812 11060 11824
rect 9272 11784 11060 11812
rect 9272 11772 9278 11784
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 11296 11784 11561 11812
rect 11296 11772 11302 11784
rect 8389 11747 8447 11753
rect 8389 11744 8401 11747
rect 7944 11716 8401 11744
rect 6917 11679 6975 11685
rect 6917 11676 6929 11679
rect 4939 11648 5304 11676
rect 6656 11648 6929 11676
rect 4939 11645 4951 11648
rect 4893 11639 4951 11645
rect 4617 11615 4675 11621
rect 5276 11620 5304 11648
rect 6917 11645 6929 11648
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 7650 11636 7656 11688
rect 7708 11636 7714 11688
rect 7742 11636 7748 11688
rect 7800 11636 7806 11688
rect 7944 11685 7972 11716
rect 8389 11713 8401 11716
rect 8435 11713 8447 11747
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 8389 11707 8447 11713
rect 9508 11716 9781 11744
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 8018 11636 8024 11688
rect 8076 11636 8082 11688
rect 9508 11685 9536 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11533 11744 11561 11784
rect 12544 11784 13952 11812
rect 12544 11756 12572 11784
rect 10836 11716 11468 11744
rect 11533 11716 12112 11744
rect 10836 11704 10842 11716
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 8251 11648 8861 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 4982 11608 4988 11620
rect 4816 11580 4988 11608
rect 3510 11500 3516 11552
rect 3568 11500 3574 11552
rect 3970 11500 3976 11552
rect 4028 11500 4034 11552
rect 4816 11549 4844 11580
rect 4982 11568 4988 11580
rect 5040 11608 5046 11620
rect 5138 11611 5196 11617
rect 5138 11608 5150 11611
rect 5040 11580 5150 11608
rect 5040 11568 5046 11580
rect 5138 11577 5150 11580
rect 5184 11577 5196 11611
rect 5138 11571 5196 11577
rect 5258 11568 5264 11620
rect 5316 11568 5322 11620
rect 6288 11580 7512 11608
rect 6288 11549 6316 11580
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 6273 11543 6331 11549
rect 6273 11509 6285 11543
rect 6319 11509 6331 11543
rect 6273 11503 6331 11509
rect 6730 11500 6736 11552
rect 6788 11500 6794 11552
rect 7484 11540 7512 11580
rect 7558 11568 7564 11620
rect 7616 11608 7622 11620
rect 8113 11611 8171 11617
rect 8113 11608 8125 11611
rect 7616 11580 8125 11608
rect 7616 11568 7622 11580
rect 8113 11577 8125 11580
rect 8159 11577 8171 11611
rect 8864 11608 8892 11639
rect 9582 11636 9588 11688
rect 9640 11636 9646 11688
rect 9674 11636 9680 11688
rect 9732 11636 9738 11688
rect 11054 11636 11060 11688
rect 11112 11636 11118 11688
rect 11440 11685 11468 11716
rect 11150 11679 11208 11685
rect 11150 11645 11162 11679
rect 11196 11645 11208 11679
rect 11150 11639 11208 11645
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 11563 11679 11621 11685
rect 11563 11645 11575 11679
rect 11609 11676 11621 11679
rect 11882 11676 11888 11688
rect 11609 11648 11888 11676
rect 11609 11645 11621 11648
rect 11563 11639 11621 11645
rect 9398 11608 9404 11620
rect 8864 11580 9404 11608
rect 8113 11571 8171 11577
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 9600 11608 9628 11636
rect 11164 11608 11192 11639
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 12084 11685 12112 11716
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 12986 11704 12992 11756
rect 13044 11704 13050 11756
rect 13170 11704 13176 11756
rect 13228 11704 13234 11756
rect 11977 11679 12035 11685
rect 11977 11645 11989 11679
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11676 12127 11679
rect 12434 11676 12440 11688
rect 12115 11648 12440 11676
rect 12115 11645 12127 11648
rect 12069 11639 12127 11645
rect 9600 11580 11192 11608
rect 11330 11568 11336 11620
rect 11388 11568 11394 11620
rect 11790 11568 11796 11620
rect 11848 11568 11854 11620
rect 11992 11608 12020 11639
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 12618 11636 12624 11688
rect 12676 11636 12682 11688
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11676 12863 11679
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12851 11648 12909 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 13004 11676 13032 11704
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13004 11648 13645 11676
rect 12897 11639 12955 11645
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 13814 11676 13820 11688
rect 13771 11648 13820 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 13924 11685 13952 11784
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 15320 11676 15348 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 18325 11883 18383 11889
rect 18325 11849 18337 11883
rect 18371 11880 18383 11883
rect 18506 11880 18512 11892
rect 18371 11852 18512 11880
rect 18371 11849 18383 11852
rect 18325 11843 18383 11849
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 19150 11840 19156 11892
rect 19208 11840 19214 11892
rect 19705 11883 19763 11889
rect 19705 11880 19717 11883
rect 19260 11852 19717 11880
rect 17497 11815 17555 11821
rect 17497 11781 17509 11815
rect 17543 11812 17555 11815
rect 17957 11815 18015 11821
rect 17957 11812 17969 11815
rect 17543 11784 17969 11812
rect 17543 11781 17555 11784
rect 17497 11775 17555 11781
rect 17957 11781 17969 11784
rect 18003 11812 18015 11815
rect 18003 11784 18092 11812
rect 18003 11781 18015 11784
rect 17957 11775 18015 11781
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 15948 11716 17693 11744
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 13955 11648 15393 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 15381 11645 15393 11648
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 15470 11636 15476 11688
rect 15528 11676 15534 11688
rect 15565 11679 15623 11685
rect 15565 11676 15577 11679
rect 15528 11648 15577 11676
rect 15528 11636 15534 11648
rect 15565 11645 15577 11648
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11676 15715 11679
rect 15838 11676 15844 11688
rect 15703 11648 15844 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 11905 11580 12020 11608
rect 12713 11611 12771 11617
rect 7650 11540 7656 11552
rect 7484 11512 7656 11540
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 7984 11512 9597 11540
rect 7984 11500 7990 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9858 11540 9864 11552
rect 9732 11512 9864 11540
rect 9732 11500 9738 11512
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 11905 11540 11933 11580
rect 12713 11577 12725 11611
rect 12759 11608 12771 11611
rect 15948 11608 15976 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17788 11716 18000 11744
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 16448 11648 17601 11676
rect 16448 11636 16454 11648
rect 17589 11645 17601 11648
rect 17635 11676 17647 11679
rect 17788 11676 17816 11716
rect 17635 11648 17816 11676
rect 17635 11645 17647 11648
rect 17589 11639 17647 11645
rect 17862 11636 17868 11688
rect 17920 11636 17926 11688
rect 17972 11685 18000 11716
rect 17957 11679 18015 11685
rect 17957 11645 17969 11679
rect 18003 11645 18015 11679
rect 18064 11676 18092 11784
rect 18138 11772 18144 11824
rect 18196 11812 18202 11824
rect 19260 11812 19288 11852
rect 19705 11849 19717 11852
rect 19751 11880 19763 11883
rect 20070 11880 20076 11892
rect 19751 11852 20076 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 21082 11880 21088 11892
rect 20312 11852 21088 11880
rect 20312 11840 20318 11852
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21450 11840 21456 11892
rect 21508 11840 21514 11892
rect 21545 11883 21603 11889
rect 21545 11849 21557 11883
rect 21591 11880 21603 11883
rect 22002 11880 22008 11892
rect 21591 11852 22008 11880
rect 21591 11849 21603 11852
rect 21545 11843 21603 11849
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 23290 11880 23296 11892
rect 23032 11852 23296 11880
rect 18196 11784 19288 11812
rect 18196 11772 18202 11784
rect 19518 11772 19524 11824
rect 19576 11812 19582 11824
rect 19613 11815 19671 11821
rect 19613 11812 19625 11815
rect 19576 11784 19625 11812
rect 19576 11772 19582 11784
rect 19613 11781 19625 11784
rect 19659 11781 19671 11815
rect 21468 11812 21496 11840
rect 22738 11812 22744 11824
rect 21468 11784 22744 11812
rect 19613 11775 19671 11781
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 22833 11815 22891 11821
rect 22833 11781 22845 11815
rect 22879 11812 22891 11815
rect 23032 11812 23060 11852
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 23474 11840 23480 11892
rect 23532 11840 23538 11892
rect 24029 11883 24087 11889
rect 24029 11849 24041 11883
rect 24075 11880 24087 11883
rect 24118 11880 24124 11892
rect 24075 11852 24124 11880
rect 24075 11849 24087 11852
rect 24029 11843 24087 11849
rect 24118 11840 24124 11852
rect 24176 11840 24182 11892
rect 27706 11840 27712 11892
rect 27764 11840 27770 11892
rect 22879 11784 23060 11812
rect 22879 11781 22891 11784
rect 22833 11775 22891 11781
rect 19536 11744 19564 11772
rect 22848 11744 22876 11775
rect 23106 11772 23112 11824
rect 23164 11812 23170 11824
rect 23201 11815 23259 11821
rect 23201 11812 23213 11815
rect 23164 11784 23213 11812
rect 23164 11772 23170 11784
rect 23201 11781 23213 11784
rect 23247 11781 23259 11815
rect 23201 11775 23259 11781
rect 19352 11716 19564 11744
rect 19653 11716 20024 11744
rect 18138 11676 18144 11688
rect 18064 11648 18144 11676
rect 17957 11639 18015 11645
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11676 18383 11679
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18371 11648 18705 11676
rect 18371 11645 18383 11648
rect 18325 11639 18383 11645
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18874 11636 18880 11688
rect 18932 11676 18938 11688
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 18932 11648 19165 11676
rect 18932 11636 18938 11648
rect 19153 11645 19165 11648
rect 19199 11676 19211 11679
rect 19242 11676 19248 11688
rect 19199 11648 19248 11676
rect 19199 11645 19211 11648
rect 19153 11639 19211 11645
rect 19242 11636 19248 11648
rect 19300 11636 19306 11688
rect 19352 11685 19380 11716
rect 19337 11679 19395 11685
rect 19337 11645 19349 11679
rect 19383 11645 19395 11679
rect 19337 11639 19395 11645
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 19484 11648 19533 11676
rect 19484 11636 19490 11648
rect 19521 11645 19533 11648
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 12759 11580 15976 11608
rect 17313 11611 17371 11617
rect 12759 11577 12771 11580
rect 12713 11571 12771 11577
rect 17313 11577 17325 11611
rect 17359 11577 17371 11611
rect 17880 11608 17908 11636
rect 17313 11571 17371 11577
rect 17604 11580 17908 11608
rect 10744 11512 11933 11540
rect 10744 11500 10750 11512
rect 12066 11500 12072 11552
rect 12124 11500 12130 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 13814 11540 13820 11552
rect 12492 11512 13820 11540
rect 12492 11500 12498 11512
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14093 11543 14151 11549
rect 14093 11509 14105 11543
rect 14139 11540 14151 11543
rect 14274 11540 14280 11552
rect 14139 11512 14280 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 15197 11543 15255 11549
rect 15197 11509 15209 11543
rect 15243 11540 15255 11543
rect 15378 11540 15384 11552
rect 15243 11512 15384 11540
rect 15243 11509 15255 11512
rect 15197 11503 15255 11509
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 17328 11540 17356 11571
rect 17604 11549 17632 11580
rect 18046 11568 18052 11620
rect 18104 11608 18110 11620
rect 19653 11608 19681 11716
rect 19886 11676 19892 11688
rect 18104 11580 19681 11608
rect 19720 11648 19892 11676
rect 18104 11568 18110 11580
rect 15528 11512 17356 11540
rect 17589 11543 17647 11549
rect 15528 11500 15534 11512
rect 17589 11509 17601 11543
rect 17635 11509 17647 11543
rect 17589 11503 17647 11509
rect 17678 11500 17684 11552
rect 17736 11540 17742 11552
rect 19720 11540 19748 11648
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 19996 11676 20024 11716
rect 22664 11716 22876 11744
rect 22186 11676 22192 11688
rect 19996 11648 22192 11676
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 22664 11685 22692 11716
rect 22922 11704 22928 11756
rect 22980 11704 22986 11756
rect 23017 11747 23075 11753
rect 23017 11713 23029 11747
rect 23063 11744 23075 11747
rect 23385 11747 23443 11753
rect 23063 11716 23244 11744
rect 23063 11713 23075 11716
rect 23017 11707 23075 11713
rect 22373 11679 22431 11685
rect 22373 11645 22385 11679
rect 22419 11676 22431 11679
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 22419 11648 22477 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 22465 11645 22477 11648
rect 22511 11645 22523 11679
rect 22465 11639 22523 11645
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11645 22707 11679
rect 22649 11639 22707 11645
rect 22738 11636 22744 11688
rect 22796 11636 22802 11688
rect 22940 11676 22968 11704
rect 23216 11688 23244 11716
rect 23385 11713 23397 11747
rect 23431 11744 23443 11747
rect 23492 11744 23520 11840
rect 23431 11716 23520 11744
rect 23431 11713 23443 11716
rect 23385 11707 23443 11713
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 23716 11716 27568 11744
rect 23716 11704 23722 11716
rect 23109 11679 23167 11685
rect 23109 11676 23121 11679
rect 22940 11648 23121 11676
rect 23109 11645 23121 11648
rect 23155 11645 23167 11679
rect 23109 11639 23167 11645
rect 23198 11636 23204 11688
rect 23256 11636 23262 11688
rect 23566 11636 23572 11688
rect 23624 11676 23630 11688
rect 23845 11679 23903 11685
rect 23845 11676 23857 11679
rect 23624 11648 23857 11676
rect 23624 11636 23630 11648
rect 23845 11645 23857 11648
rect 23891 11645 23903 11679
rect 25961 11679 26019 11685
rect 25961 11676 25973 11679
rect 23845 11639 23903 11645
rect 24826 11648 25973 11676
rect 20162 11617 20168 11620
rect 19797 11611 19855 11617
rect 19797 11577 19809 11611
rect 19843 11577 19855 11611
rect 19797 11571 19855 11577
rect 20156 11571 20168 11617
rect 17736 11512 19748 11540
rect 19812 11540 19840 11571
rect 20162 11568 20168 11571
rect 20220 11568 20226 11620
rect 23014 11608 23020 11620
rect 22756 11580 23020 11608
rect 20254 11540 20260 11552
rect 19812 11512 20260 11540
rect 17736 11500 17742 11512
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21818 11540 21824 11552
rect 21315 11512 21824 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 22554 11500 22560 11552
rect 22612 11500 22618 11552
rect 22756 11549 22784 11580
rect 23014 11568 23020 11580
rect 23072 11568 23078 11620
rect 22741 11543 22799 11549
rect 22741 11509 22753 11543
rect 22787 11509 22799 11543
rect 22741 11503 22799 11509
rect 22830 11500 22836 11552
rect 22888 11540 22894 11552
rect 24826 11540 24854 11648
rect 25961 11645 25973 11648
rect 26007 11645 26019 11679
rect 25961 11639 26019 11645
rect 26234 11636 26240 11688
rect 26292 11636 26298 11688
rect 26326 11636 26332 11688
rect 26384 11676 26390 11688
rect 26421 11679 26479 11685
rect 26421 11676 26433 11679
rect 26384 11648 26433 11676
rect 26384 11636 26390 11648
rect 26421 11645 26433 11648
rect 26467 11645 26479 11679
rect 26421 11639 26479 11645
rect 26694 11636 26700 11688
rect 26752 11636 26758 11688
rect 27246 11636 27252 11688
rect 27304 11636 27310 11688
rect 27540 11685 27568 11716
rect 27525 11679 27583 11685
rect 27525 11645 27537 11679
rect 27571 11645 27583 11679
rect 27525 11639 27583 11645
rect 22888 11512 24854 11540
rect 22888 11500 22894 11512
rect 26142 11500 26148 11552
rect 26200 11500 26206 11552
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 2225 11339 2283 11345
rect 2225 11305 2237 11339
rect 2271 11336 2283 11339
rect 3418 11336 3424 11348
rect 2271 11308 3424 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 3970 11336 3976 11348
rect 3528 11308 3976 11336
rect 3528 11268 3556 11308
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4614 11296 4620 11348
rect 4672 11296 4678 11348
rect 4982 11296 4988 11348
rect 5040 11296 5046 11348
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 7098 11296 7104 11348
rect 7156 11296 7162 11348
rect 7282 11296 7288 11348
rect 7340 11296 7346 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 7742 11336 7748 11348
rect 7699 11308 7748 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 8665 11339 8723 11345
rect 8352 11308 8616 11336
rect 8352 11296 8358 11308
rect 3266 11240 3556 11268
rect 3697 11271 3755 11277
rect 3697 11237 3709 11271
rect 3743 11268 3755 11271
rect 3786 11268 3792 11280
rect 3743 11240 3792 11268
rect 3743 11237 3755 11240
rect 3697 11231 3755 11237
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 4632 11200 4660 11296
rect 6012 11209 6040 11296
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 4632 11172 5181 11200
rect 5169 11169 5181 11172
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5997 11203 6055 11209
rect 5997 11169 6009 11203
rect 6043 11169 6055 11203
rect 7116 11200 7144 11296
rect 7300 11268 7328 11296
rect 8588 11268 8616 11308
rect 8665 11305 8677 11339
rect 8711 11336 8723 11339
rect 9309 11339 9367 11345
rect 8711 11308 9168 11336
rect 8711 11305 8723 11308
rect 8665 11299 8723 11305
rect 8849 11271 8907 11277
rect 8849 11268 8861 11271
rect 7300 11240 7696 11268
rect 8588 11240 8861 11268
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 7116 11172 7297 11200
rect 5997 11163 6055 11169
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7558 11160 7564 11212
rect 7616 11160 7622 11212
rect 7668 11209 7696 11240
rect 8849 11237 8861 11240
rect 8895 11237 8907 11271
rect 8849 11231 8907 11237
rect 9140 11268 9168 11308
rect 9309 11305 9321 11339
rect 9355 11305 9367 11339
rect 9309 11299 9367 11305
rect 9214 11268 9220 11280
rect 9140 11240 9220 11268
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 8021 11203 8079 11209
rect 8202 11206 8208 11212
rect 8021 11200 8033 11203
rect 7699 11172 8033 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 8021 11169 8033 11172
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8128 11178 8208 11206
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3292 11104 3985 11132
rect 3292 11092 3298 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 7834 11132 7840 11144
rect 7423 11104 7840 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 8128 11141 8156 11178
rect 8202 11160 8208 11178
rect 8260 11160 8266 11212
rect 8294 11160 8300 11212
rect 8352 11160 8358 11212
rect 8662 11160 8668 11212
rect 8720 11160 8726 11212
rect 8754 11160 8760 11212
rect 8812 11160 8818 11212
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11200 8999 11203
rect 9030 11200 9036 11212
rect 8987 11172 9036 11200
rect 8987 11169 8999 11172
rect 8941 11163 8999 11169
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 9140 11209 9168 11240
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 9324 11268 9352 11299
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 9456 11308 9812 11336
rect 9456 11296 9462 11308
rect 9646 11271 9704 11277
rect 9646 11268 9658 11271
rect 9324 11240 9658 11268
rect 9646 11237 9658 11240
rect 9692 11237 9704 11271
rect 9784 11268 9812 11308
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 10744 11308 11253 11336
rect 10744 11296 10750 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 11885 11339 11943 11345
rect 11885 11336 11897 11339
rect 11848 11308 11897 11336
rect 11848 11296 11854 11308
rect 11885 11305 11897 11308
rect 11931 11305 11943 11339
rect 11885 11299 11943 11305
rect 12066 11296 12072 11348
rect 12124 11296 12130 11348
rect 13170 11336 13176 11348
rect 12544 11308 13176 11336
rect 12084 11268 12112 11296
rect 9784 11240 12112 11268
rect 9646 11231 9704 11237
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11169 9183 11203
rect 10594 11200 10600 11212
rect 9125 11163 9183 11169
rect 9232 11172 10600 11200
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8435 11104 8524 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8496 11076 8524 11104
rect 7285 11067 7343 11073
rect 7285 11064 7297 11067
rect 5184 11036 7297 11064
rect 5184 11008 5212 11036
rect 7285 11033 7297 11036
rect 7331 11064 7343 11067
rect 7745 11067 7803 11073
rect 7745 11064 7757 11067
rect 7331 11036 7757 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 7745 11033 7757 11036
rect 7791 11033 7803 11067
rect 7745 11027 7803 11033
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 5166 10956 5172 11008
rect 5224 10956 5230 11008
rect 5813 10999 5871 11005
rect 5813 10965 5825 10999
rect 5859 10996 5871 10999
rect 5902 10996 5908 11008
rect 5859 10968 5908 10996
rect 5859 10965 5871 10968
rect 5813 10959 5871 10965
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 7760 10996 7788 11027
rect 7926 10996 7932 11008
rect 7760 10968 7932 10996
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8036 10996 8064 11027
rect 8478 11024 8484 11076
rect 8536 11024 8542 11076
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 9232 11064 9260 11172
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 11238 11200 11244 11212
rect 10704 11172 11244 11200
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 8619 11036 9260 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 8110 10996 8116 11008
rect 8036 10968 8116 10996
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8588 10996 8616 11027
rect 8352 10968 8616 10996
rect 8352 10956 8358 10968
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 10704 10996 10732 11172
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11348 11209 11376 11240
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11480 11172 11805 11200
rect 11480 11160 11486 11172
rect 11793 11169 11805 11172
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 12434 11200 12440 11212
rect 12023 11172 12440 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 12544 11209 12572 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13633 11339 13691 11345
rect 13633 11305 13645 11339
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 13648 11268 13676 11299
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 16114 11336 16120 11348
rect 13872 11308 16120 11336
rect 13872 11296 13878 11308
rect 16114 11296 16120 11308
rect 16172 11336 16178 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 16172 11308 16221 11336
rect 16172 11296 16178 11308
rect 16209 11305 16221 11308
rect 16255 11336 16267 11339
rect 18046 11336 18052 11348
rect 16255 11308 16712 11336
rect 16255 11305 16267 11308
rect 16209 11299 16267 11305
rect 13970 11271 14028 11277
rect 13970 11268 13982 11271
rect 12728 11240 13492 11268
rect 13648 11240 13982 11268
rect 12728 11209 12756 11240
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11169 12587 11203
rect 12529 11163 12587 11169
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11169 12771 11203
rect 12713 11163 12771 11169
rect 12805 11203 12863 11209
rect 12805 11169 12817 11203
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 13354 11200 13360 11212
rect 13035 11172 13360 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11132 11575 11135
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 11563 11104 12633 11132
rect 11563 11101 11575 11104
rect 11517 11095 11575 11101
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 12820 11064 12848 11163
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 13464 11209 13492 11240
rect 13970 11237 13982 11240
rect 14016 11237 14028 11271
rect 15473 11271 15531 11277
rect 15473 11268 15485 11271
rect 13970 11231 14028 11237
rect 15120 11240 15485 11268
rect 15120 11212 15148 11240
rect 15473 11237 15485 11240
rect 15519 11237 15531 11271
rect 16298 11268 16304 11280
rect 15473 11231 15531 11237
rect 15580 11240 16304 11268
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11200 13507 11203
rect 13495 11172 14780 11200
rect 13495 11169 13507 11172
rect 13449 11163 13507 11169
rect 13725 11135 13783 11141
rect 13725 11132 13737 11135
rect 11440 11036 12848 11064
rect 12912 11104 13737 11132
rect 11440 11008 11468 11036
rect 8720 10968 10732 10996
rect 8720 10956 8726 10968
rect 10778 10956 10784 11008
rect 10836 10956 10842 11008
rect 11422 10956 11428 11008
rect 11480 10956 11486 11008
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 12912 10996 12940 11104
rect 13725 11101 13737 11104
rect 13771 11101 13783 11135
rect 14752 11132 14780 11172
rect 15102 11160 15108 11212
rect 15160 11160 15166 11212
rect 15194 11160 15200 11212
rect 15252 11160 15258 11212
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 15580 11209 15608 11240
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 16390 11228 16396 11280
rect 16448 11228 16454 11280
rect 16482 11228 16488 11280
rect 16540 11228 16546 11280
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 15344 11172 15393 11200
rect 15344 11160 15350 11172
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 16408 11200 16436 11228
rect 16684 11209 16712 11308
rect 17052 11308 18052 11336
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 16255 11172 16589 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 16577 11169 16589 11172
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11169 16727 11203
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 16669 11163 16727 11169
rect 16776 11172 16957 11200
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 14752 11104 16313 11132
rect 13725 11095 13783 11101
rect 16301 11101 16313 11104
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 12989 11067 13047 11073
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 15470 11064 15476 11076
rect 13035 11036 13768 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 11572 10968 12940 10996
rect 13740 10996 13768 11036
rect 14660 11036 15476 11064
rect 14660 10996 14688 11036
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 16316 11064 16344 11095
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 16316 11036 16589 11064
rect 16577 11033 16589 11036
rect 16623 11033 16635 11067
rect 16776 11064 16804 11172
rect 16945 11169 16957 11172
rect 16991 11169 17003 11203
rect 17052 11204 17080 11308
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18138 11296 18144 11348
rect 18196 11296 18202 11348
rect 18325 11339 18383 11345
rect 18325 11305 18337 11339
rect 18371 11305 18383 11339
rect 18325 11299 18383 11305
rect 18156 11268 18184 11296
rect 17880 11240 18184 11268
rect 18340 11268 18368 11299
rect 19518 11296 19524 11348
rect 19576 11296 19582 11348
rect 20073 11339 20131 11345
rect 20073 11305 20085 11339
rect 20119 11336 20131 11339
rect 20162 11336 20168 11348
rect 20119 11308 20168 11336
rect 20119 11305 20131 11308
rect 20073 11299 20131 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20254 11296 20260 11348
rect 20312 11336 20318 11348
rect 20349 11339 20407 11345
rect 20349 11336 20361 11339
rect 20312 11308 20361 11336
rect 20312 11296 20318 11308
rect 20349 11305 20361 11308
rect 20395 11305 20407 11339
rect 20349 11299 20407 11305
rect 20622 11296 20628 11348
rect 20680 11296 20686 11348
rect 21450 11296 21456 11348
rect 21508 11296 21514 11348
rect 22741 11339 22799 11345
rect 22741 11336 22753 11339
rect 22204 11308 22753 11336
rect 18662 11271 18720 11277
rect 18662 11268 18674 11271
rect 18340 11240 18674 11268
rect 17129 11204 17187 11209
rect 17052 11203 17187 11204
rect 17052 11176 17141 11203
rect 16945 11163 17003 11169
rect 17129 11169 17141 11176
rect 17175 11169 17187 11203
rect 17129 11163 17187 11169
rect 17218 11160 17224 11212
rect 17276 11160 17282 11212
rect 17880 11209 17908 11240
rect 18662 11237 18674 11240
rect 18708 11237 18720 11271
rect 18662 11231 18720 11237
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 17405 11163 17463 11169
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 16853 11135 16911 11141
rect 16853 11101 16865 11135
rect 16899 11132 16911 11135
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 16899 11104 17049 11132
rect 16899 11101 16911 11104
rect 16853 11095 16911 11101
rect 17037 11101 17049 11104
rect 17083 11101 17095 11135
rect 17420 11132 17448 11163
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18141 11203 18199 11209
rect 18141 11200 18153 11203
rect 18012 11172 18153 11200
rect 18012 11160 18018 11172
rect 18141 11169 18153 11172
rect 18187 11169 18199 11203
rect 19536 11200 19564 11296
rect 20640 11268 20668 11296
rect 20272 11240 20668 11268
rect 20272 11209 20300 11240
rect 19889 11203 19947 11209
rect 19889 11200 19901 11203
rect 18141 11163 18199 11169
rect 18340 11172 19472 11200
rect 19536 11172 19901 11200
rect 18340 11132 18368 11172
rect 17420 11104 18368 11132
rect 17037 11095 17095 11101
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 19444 11132 19472 11172
rect 19889 11169 19901 11172
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 20257 11203 20315 11209
rect 20257 11169 20269 11203
rect 20303 11169 20315 11203
rect 20257 11163 20315 11169
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11200 20499 11203
rect 21266 11200 21272 11212
rect 20487 11172 21272 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 21468 11200 21496 11296
rect 22204 11212 22232 11308
rect 22741 11305 22753 11308
rect 22787 11336 22799 11339
rect 22830 11336 22836 11348
rect 22787 11308 22836 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 22922 11296 22928 11348
rect 22980 11296 22986 11348
rect 23014 11296 23020 11348
rect 23072 11296 23078 11348
rect 23937 11339 23995 11345
rect 23937 11305 23949 11339
rect 23983 11305 23995 11339
rect 23937 11299 23995 11305
rect 25409 11339 25467 11345
rect 25409 11305 25421 11339
rect 25455 11305 25467 11339
rect 26421 11339 26479 11345
rect 26421 11336 26433 11339
rect 25409 11299 25467 11305
rect 25884 11308 26433 11336
rect 22465 11271 22523 11277
rect 22465 11237 22477 11271
rect 22511 11268 22523 11271
rect 22554 11268 22560 11280
rect 22511 11240 22560 11268
rect 22511 11237 22523 11240
rect 22465 11231 22523 11237
rect 22554 11228 22560 11240
rect 22612 11228 22618 11280
rect 22940 11268 22968 11296
rect 22756 11240 22968 11268
rect 23032 11268 23060 11296
rect 23952 11268 23980 11299
rect 24274 11271 24332 11277
rect 24274 11268 24286 11271
rect 23032 11240 23336 11268
rect 23952 11240 24286 11268
rect 22097 11203 22155 11209
rect 22097 11200 22109 11203
rect 21468 11172 22109 11200
rect 22097 11169 22109 11172
rect 22143 11169 22155 11203
rect 22097 11163 22155 11169
rect 22186 11160 22192 11212
rect 22244 11160 22250 11212
rect 22756 11209 22784 11240
rect 22649 11203 22707 11209
rect 22649 11200 22661 11203
rect 22296 11172 22661 11200
rect 20806 11132 20812 11144
rect 19444 11104 20812 11132
rect 20806 11092 20812 11104
rect 20864 11132 20870 11144
rect 22296 11132 22324 11172
rect 22649 11169 22661 11172
rect 22695 11169 22707 11203
rect 22649 11163 22707 11169
rect 22741 11203 22799 11209
rect 22741 11169 22753 11203
rect 22787 11169 22799 11203
rect 22741 11163 22799 11169
rect 22830 11160 22836 11212
rect 22888 11160 22894 11212
rect 23308 11209 23336 11240
rect 24274 11237 24286 11240
rect 24320 11237 24332 11271
rect 25424 11268 25452 11299
rect 25424 11240 25636 11268
rect 24274 11231 24332 11237
rect 23109 11203 23167 11209
rect 23109 11169 23121 11203
rect 23155 11169 23167 11203
rect 23109 11163 23167 11169
rect 23293 11203 23351 11209
rect 23293 11169 23305 11203
rect 23339 11200 23351 11203
rect 23753 11203 23811 11209
rect 23753 11200 23765 11203
rect 23339 11172 23765 11200
rect 23339 11169 23351 11172
rect 23293 11163 23351 11169
rect 23753 11169 23765 11172
rect 23799 11169 23811 11203
rect 23753 11163 23811 11169
rect 20864 11104 22324 11132
rect 22373 11135 22431 11141
rect 20864 11092 20870 11104
rect 17497 11067 17555 11073
rect 17497 11064 17509 11067
rect 16776 11036 17509 11064
rect 16577 11027 16635 11033
rect 17497 11033 17509 11036
rect 17543 11033 17555 11067
rect 17497 11027 17555 11033
rect 19797 11067 19855 11073
rect 19797 11033 19809 11067
rect 19843 11064 19855 11067
rect 20162 11064 20168 11076
rect 19843 11036 20168 11064
rect 19843 11033 19855 11036
rect 19797 11027 19855 11033
rect 20162 11024 20168 11036
rect 20220 11024 20226 11076
rect 22112 11073 22140 11104
rect 22373 11101 22385 11135
rect 22419 11132 22431 11135
rect 23014 11132 23020 11144
rect 22419 11104 23020 11132
rect 22419 11101 22431 11104
rect 22373 11095 22431 11101
rect 23014 11092 23020 11104
rect 23072 11092 23078 11144
rect 23124 11132 23152 11163
rect 25222 11160 25228 11212
rect 25280 11200 25286 11212
rect 25608 11209 25636 11240
rect 25774 11228 25780 11280
rect 25832 11228 25838 11280
rect 25884 11277 25912 11308
rect 26421 11305 26433 11308
rect 26467 11305 26479 11339
rect 26421 11299 26479 11305
rect 25869 11271 25927 11277
rect 25869 11237 25881 11271
rect 25915 11237 25927 11271
rect 25869 11231 25927 11237
rect 26142 11228 26148 11280
rect 26200 11268 26206 11280
rect 27534 11271 27592 11277
rect 27534 11268 27546 11271
rect 26200 11240 27546 11268
rect 26200 11228 26206 11240
rect 27534 11237 27546 11240
rect 27580 11237 27592 11271
rect 27534 11231 27592 11237
rect 25501 11203 25559 11209
rect 25501 11200 25513 11203
rect 25280 11172 25513 11200
rect 25280 11160 25286 11172
rect 25501 11169 25513 11172
rect 25547 11169 25559 11203
rect 25501 11163 25559 11169
rect 25594 11203 25652 11209
rect 25594 11169 25606 11203
rect 25640 11169 25652 11203
rect 25594 11163 25652 11169
rect 25958 11160 25964 11212
rect 26016 11209 26022 11212
rect 26016 11200 26024 11209
rect 28074 11200 28080 11212
rect 26016 11172 28080 11200
rect 26016 11163 26024 11172
rect 26016 11160 26022 11163
rect 28074 11160 28080 11172
rect 28132 11160 28138 11212
rect 29270 11160 29276 11212
rect 29328 11160 29334 11212
rect 23124 11104 23244 11132
rect 22097 11067 22155 11073
rect 22097 11033 22109 11067
rect 22143 11064 22155 11067
rect 23216 11064 23244 11104
rect 23658 11092 23664 11144
rect 23716 11132 23722 11144
rect 23842 11132 23848 11144
rect 23716 11104 23848 11132
rect 23716 11092 23722 11104
rect 23842 11092 23848 11104
rect 23900 11132 23906 11144
rect 24029 11135 24087 11141
rect 24029 11132 24041 11135
rect 23900 11104 24041 11132
rect 23900 11092 23906 11104
rect 24029 11101 24041 11104
rect 24075 11101 24087 11135
rect 24029 11095 24087 11101
rect 27801 11135 27859 11141
rect 27801 11101 27813 11135
rect 27847 11132 27859 11135
rect 27982 11132 27988 11144
rect 27847 11104 27988 11132
rect 27847 11101 27859 11104
rect 27801 11095 27859 11101
rect 27982 11092 27988 11104
rect 28040 11132 28046 11144
rect 28994 11132 29000 11144
rect 28040 11104 29000 11132
rect 28040 11092 28046 11104
rect 28994 11092 29000 11104
rect 29052 11132 29058 11144
rect 29288 11132 29316 11160
rect 29052 11104 29316 11132
rect 29052 11092 29058 11104
rect 22143 11036 22177 11064
rect 22296 11036 23244 11064
rect 22143 11033 22155 11036
rect 22097 11027 22155 11033
rect 13740 10968 14688 10996
rect 11572 10956 11578 10968
rect 15102 10956 15108 11008
rect 15160 10956 15166 11008
rect 15746 10956 15752 11008
rect 15804 10956 15810 11008
rect 16482 10956 16488 11008
rect 16540 10996 16546 11008
rect 17221 10999 17279 11005
rect 17221 10996 17233 10999
rect 16540 10968 17233 10996
rect 16540 10956 16546 10968
rect 17221 10965 17233 10968
rect 17267 10965 17279 10999
rect 17221 10959 17279 10965
rect 18049 10999 18107 11005
rect 18049 10965 18061 10999
rect 18095 10996 18107 10999
rect 18782 10996 18788 11008
rect 18095 10968 18788 10996
rect 18095 10965 18107 10968
rect 18049 10959 18107 10965
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 21082 10956 21088 11008
rect 21140 10996 21146 11008
rect 22296 10996 22324 11036
rect 21140 10968 22324 10996
rect 21140 10956 21146 10968
rect 23014 10956 23020 11008
rect 23072 10956 23078 11008
rect 23106 10956 23112 11008
rect 23164 10956 23170 11008
rect 23216 10996 23244 11036
rect 26068 11036 26924 11064
rect 26068 10996 26096 11036
rect 23216 10968 26096 10996
rect 26142 10956 26148 11008
rect 26200 10956 26206 11008
rect 26896 10996 26924 11036
rect 27154 10996 27160 11008
rect 26896 10968 27160 10996
rect 27154 10956 27160 10968
rect 27212 10956 27218 11008
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 1029 10795 1087 10801
rect 1029 10761 1041 10795
rect 1075 10792 1087 10795
rect 4801 10795 4859 10801
rect 1075 10764 2774 10792
rect 1075 10761 1087 10764
rect 1029 10755 1087 10761
rect 842 10548 848 10600
rect 900 10548 906 10600
rect 2746 10520 2774 10764
rect 3436 10764 4384 10792
rect 3436 10665 3464 10764
rect 4356 10724 4384 10764
rect 4801 10761 4813 10795
rect 4847 10792 4859 10795
rect 10134 10792 10140 10804
rect 4847 10764 10140 10792
rect 4847 10761 4859 10764
rect 4801 10755 4859 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10594 10752 10600 10804
rect 10652 10792 10658 10804
rect 11241 10795 11299 10801
rect 10652 10764 11193 10792
rect 10652 10752 10658 10764
rect 7009 10727 7067 10733
rect 4356 10696 5304 10724
rect 5276 10668 5304 10696
rect 7009 10693 7021 10727
rect 7055 10724 7067 10727
rect 10413 10727 10471 10733
rect 7055 10696 10088 10724
rect 7055 10693 7067 10696
rect 7009 10687 7067 10693
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5316 10628 5641 10656
rect 5316 10616 5322 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8754 10656 8760 10668
rect 7984 10628 8760 10656
rect 7984 10616 7990 10628
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 10060 10665 10088 10696
rect 10413 10693 10425 10727
rect 10459 10724 10471 10727
rect 10686 10724 10692 10736
rect 10459 10696 10692 10724
rect 10459 10693 10471 10696
rect 10413 10687 10471 10693
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10625 10103 10659
rect 11165 10656 11193 10764
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 11287 10764 14197 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 14185 10755 14243 10761
rect 15565 10795 15623 10801
rect 15565 10761 15577 10795
rect 15611 10792 15623 10795
rect 15746 10792 15752 10804
rect 15611 10764 15752 10792
rect 15611 10761 15623 10764
rect 15565 10755 15623 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 22278 10792 22284 10804
rect 18288 10764 22284 10792
rect 18288 10752 18294 10764
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 14093 10727 14151 10733
rect 14093 10693 14105 10727
rect 14139 10693 14151 10727
rect 14093 10687 14151 10693
rect 10045 10619 10103 10625
rect 10244 10628 11100 10656
rect 11165 10628 11376 10656
rect 3510 10548 3516 10600
rect 3568 10588 3574 10600
rect 3677 10591 3735 10597
rect 3677 10588 3689 10591
rect 3568 10560 3689 10588
rect 3568 10548 3574 10560
rect 3677 10557 3689 10560
rect 3723 10557 3735 10591
rect 3677 10551 3735 10557
rect 5166 10548 5172 10600
rect 5224 10548 5230 10600
rect 5902 10597 5908 10600
rect 5896 10588 5908 10597
rect 5863 10560 5908 10588
rect 5896 10551 5908 10560
rect 5902 10548 5908 10551
rect 5960 10548 5966 10600
rect 7760 10573 7788 10616
rect 7745 10567 7803 10573
rect 7745 10533 7757 10567
rect 7791 10533 7803 10567
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 10244 10597 10272 10628
rect 10229 10591 10287 10597
rect 7892 10560 10180 10588
rect 7892 10548 7898 10560
rect 7745 10527 7803 10533
rect 8478 10520 8484 10532
rect 2746 10492 7696 10520
rect 4982 10412 4988 10464
rect 5040 10412 5046 10464
rect 7668 10452 7696 10492
rect 7852 10492 8484 10520
rect 7852 10452 7880 10492
rect 8478 10480 8484 10492
rect 8536 10480 8542 10532
rect 10152 10520 10180 10560
rect 10229 10557 10241 10591
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 10704 10520 10732 10551
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 11072 10597 11100 10628
rect 10965 10591 11023 10597
rect 10965 10588 10977 10591
rect 10836 10560 10977 10588
rect 10836 10548 10842 10560
rect 10965 10557 10977 10560
rect 11011 10557 11023 10591
rect 10965 10551 11023 10557
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11146 10588 11152 10600
rect 11103 10560 11152 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11348 10588 11376 10628
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11572 10628 11713 10656
rect 11572 10616 11578 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11422 10588 11428 10600
rect 11348 10560 11428 10588
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 13541 10591 13599 10597
rect 13541 10588 13553 10591
rect 13096 10560 13553 10588
rect 10152 10492 10732 10520
rect 10873 10523 10931 10529
rect 10873 10489 10885 10523
rect 10919 10520 10931 10523
rect 11514 10520 11520 10532
rect 10919 10492 11520 10520
rect 10919 10489 10931 10492
rect 10873 10483 10931 10489
rect 7668 10424 7880 10452
rect 7926 10412 7932 10464
rect 7984 10412 7990 10464
rect 10594 10412 10600 10464
rect 10652 10452 10658 10464
rect 10888 10452 10916 10483
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 11946 10523 12004 10529
rect 11946 10520 11958 10523
rect 11624 10492 11958 10520
rect 11624 10461 11652 10492
rect 11946 10489 11958 10492
rect 11992 10489 12004 10523
rect 11946 10483 12004 10489
rect 13096 10461 13124 10560
rect 13541 10557 13553 10560
rect 13587 10557 13599 10591
rect 13541 10551 13599 10557
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 13998 10588 14004 10600
rect 13955 10560 14004 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14108 10588 14136 10687
rect 20714 10684 20720 10736
rect 20772 10684 20778 10736
rect 14274 10616 14280 10668
rect 14332 10616 14338 10668
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15436 10628 15485 10656
rect 15436 10616 15442 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 20732 10656 20760 10684
rect 16172 10628 16252 10656
rect 20732 10628 21588 10656
rect 16172 10616 16178 10628
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 14108 10560 14197 10588
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14734 10548 14740 10600
rect 14792 10548 14798 10600
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 16224 10597 16252 10628
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 14976 10560 15577 10588
rect 14976 10548 14982 10560
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 18693 10591 18751 10597
rect 18693 10557 18705 10591
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 13725 10523 13783 10529
rect 13725 10489 13737 10523
rect 13771 10489 13783 10523
rect 13725 10483 13783 10489
rect 13817 10523 13875 10529
rect 13817 10489 13829 10523
rect 13863 10520 13875 10523
rect 14752 10520 14780 10548
rect 13863 10492 14780 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 10652 10424 10916 10452
rect 11609 10455 11667 10461
rect 10652 10412 10658 10424
rect 11609 10421 11621 10455
rect 11655 10421 11667 10455
rect 11609 10415 11667 10421
rect 13081 10455 13139 10461
rect 13081 10421 13093 10455
rect 13127 10421 13139 10455
rect 13740 10452 13768 10483
rect 15378 10480 15384 10532
rect 15436 10520 15442 10532
rect 15841 10523 15899 10529
rect 15841 10520 15853 10523
rect 15436 10492 15853 10520
rect 15436 10480 15442 10492
rect 15841 10489 15853 10492
rect 15887 10489 15899 10523
rect 18414 10520 18420 10532
rect 15841 10483 15899 10489
rect 16224 10492 18420 10520
rect 16224 10464 16252 10492
rect 18414 10480 18420 10492
rect 18472 10520 18478 10532
rect 18708 10520 18736 10551
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 18949 10591 19007 10597
rect 18949 10588 18961 10591
rect 18840 10560 18961 10588
rect 18840 10548 18846 10560
rect 18949 10557 18961 10560
rect 18995 10557 19007 10591
rect 18949 10551 19007 10557
rect 20717 10591 20775 10597
rect 20717 10557 20729 10591
rect 20763 10588 20775 10591
rect 20806 10588 20812 10600
rect 20763 10560 20812 10588
rect 20763 10557 20775 10560
rect 20717 10551 20775 10557
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 21560 10597 21588 10628
rect 25590 10616 25596 10668
rect 25648 10616 25654 10668
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10557 21603 10591
rect 21545 10551 21603 10557
rect 21726 10548 21732 10600
rect 21784 10548 21790 10600
rect 21818 10548 21824 10600
rect 21876 10588 21882 10600
rect 21913 10591 21971 10597
rect 21913 10588 21925 10591
rect 21876 10560 21925 10588
rect 21876 10548 21882 10560
rect 21913 10557 21925 10560
rect 21959 10557 21971 10591
rect 21913 10551 21971 10557
rect 23014 10548 23020 10600
rect 23072 10588 23078 10600
rect 23394 10591 23452 10597
rect 23394 10588 23406 10591
rect 23072 10560 23406 10588
rect 23072 10548 23078 10560
rect 23394 10557 23406 10560
rect 23440 10557 23452 10591
rect 23394 10551 23452 10557
rect 23658 10548 23664 10600
rect 23716 10548 23722 10600
rect 25130 10548 25136 10600
rect 25188 10548 25194 10600
rect 25314 10548 25320 10600
rect 25372 10548 25378 10600
rect 25685 10591 25743 10597
rect 25685 10557 25697 10591
rect 25731 10588 25743 10591
rect 26142 10588 26148 10600
rect 25731 10560 26148 10588
rect 25731 10557 25743 10560
rect 25685 10551 25743 10557
rect 26142 10548 26148 10560
rect 26200 10548 26206 10600
rect 18472 10492 18736 10520
rect 21637 10523 21695 10529
rect 18472 10480 18478 10492
rect 21637 10489 21649 10523
rect 21683 10489 21695 10523
rect 21637 10483 21695 10489
rect 14274 10452 14280 10464
rect 13740 10424 14280 10452
rect 13081 10415 13139 10421
rect 14274 10412 14280 10424
rect 14332 10412 14338 10464
rect 14553 10455 14611 10461
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 14642 10452 14648 10464
rect 14599 10424 14648 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 15197 10455 15255 10461
rect 15197 10421 15209 10455
rect 15243 10452 15255 10455
rect 15470 10452 15476 10464
rect 15243 10424 15476 10452
rect 15243 10421 15255 10424
rect 15197 10415 15255 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 15749 10455 15807 10461
rect 15749 10452 15761 10455
rect 15620 10424 15761 10452
rect 15620 10412 15626 10424
rect 15749 10421 15761 10424
rect 15795 10421 15807 10455
rect 15749 10415 15807 10421
rect 16206 10412 16212 10464
rect 16264 10412 16270 10464
rect 16390 10412 16396 10464
rect 16448 10412 16454 10464
rect 20070 10412 20076 10464
rect 20128 10412 20134 10464
rect 20898 10412 20904 10464
rect 20956 10412 20962 10464
rect 21358 10412 21364 10464
rect 21416 10412 21422 10464
rect 21652 10452 21680 10483
rect 23106 10480 23112 10532
rect 23164 10520 23170 10532
rect 23676 10520 23704 10548
rect 23164 10492 23704 10520
rect 26329 10523 26387 10529
rect 23164 10480 23170 10492
rect 26329 10489 26341 10523
rect 26375 10520 26387 10523
rect 31662 10520 31668 10532
rect 26375 10492 31668 10520
rect 26375 10489 26387 10492
rect 26329 10483 26387 10489
rect 31662 10480 31668 10492
rect 31720 10480 31726 10532
rect 22281 10455 22339 10461
rect 22281 10452 22293 10455
rect 21652 10424 22293 10452
rect 22281 10421 22293 10424
rect 22327 10421 22339 10455
rect 22281 10415 22339 10421
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 4982 10208 4988 10260
rect 5040 10208 5046 10260
rect 9692 10220 13124 10248
rect 3142 10140 3148 10192
rect 3200 10180 3206 10192
rect 3237 10183 3295 10189
rect 3237 10180 3249 10183
rect 3200 10152 3249 10180
rect 3200 10140 3206 10152
rect 3237 10149 3249 10152
rect 3283 10149 3295 10183
rect 3237 10143 3295 10149
rect 4516 10183 4574 10189
rect 4516 10149 4528 10183
rect 4562 10180 4574 10183
rect 5000 10180 5028 10208
rect 9692 10192 9720 10220
rect 4562 10152 5028 10180
rect 6448 10183 6506 10189
rect 4562 10149 4574 10152
rect 4516 10143 4574 10149
rect 6448 10149 6460 10183
rect 6494 10180 6506 10183
rect 6730 10180 6736 10192
rect 6494 10152 6736 10180
rect 6494 10149 6506 10152
rect 6448 10143 6506 10149
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 3252 9908 3280 10143
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 8846 10180 8852 10192
rect 7668 10152 8852 10180
rect 4249 10115 4307 10121
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 5258 10112 5264 10124
rect 4295 10084 5264 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 7190 10112 7196 10124
rect 6196 10084 7196 10112
rect 6196 10053 6224 10084
rect 7190 10072 7196 10084
rect 7248 10112 7254 10124
rect 7668 10121 7696 10152
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 9674 10140 9680 10192
rect 9732 10140 9738 10192
rect 9766 10140 9772 10192
rect 9824 10140 9830 10192
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 10744 10152 11100 10180
rect 10744 10140 10750 10152
rect 7926 10121 7932 10124
rect 7653 10115 7711 10121
rect 7653 10112 7665 10115
rect 7248 10084 7665 10112
rect 7248 10072 7254 10084
rect 7653 10081 7665 10084
rect 7699 10081 7711 10115
rect 7920 10112 7932 10121
rect 7887 10084 7932 10112
rect 7653 10075 7711 10081
rect 7920 10075 7932 10084
rect 7926 10072 7932 10075
rect 7984 10072 7990 10124
rect 8478 10072 8484 10124
rect 8536 10112 8542 10124
rect 9214 10112 9220 10124
rect 8536 10084 9220 10112
rect 8536 10072 8542 10084
rect 9214 10072 9220 10084
rect 9272 10112 9278 10124
rect 9401 10115 9459 10121
rect 9401 10112 9413 10115
rect 9272 10084 9413 10112
rect 9272 10072 9278 10084
rect 9401 10081 9413 10084
rect 9447 10081 9459 10115
rect 9401 10075 9459 10081
rect 9494 10115 9552 10121
rect 9494 10081 9506 10115
rect 9540 10081 9552 10115
rect 9494 10075 9552 10081
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5552 10016 6193 10044
rect 5552 9908 5580 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 9508 10044 9536 10075
rect 9858 10072 9864 10124
rect 9916 10121 9922 10124
rect 9916 10112 9924 10121
rect 9916 10084 9961 10112
rect 9916 10075 9924 10084
rect 9916 10072 9922 10075
rect 10134 10072 10140 10124
rect 10192 10072 10198 10124
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 10284 10084 10333 10112
rect 10284 10072 10290 10084
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 10321 10075 10379 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 10594 10112 10600 10124
rect 10551 10084 10600 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 10428 10044 10456 10075
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 11072 10121 11100 10152
rect 12342 10140 12348 10192
rect 12400 10180 12406 10192
rect 12437 10183 12495 10189
rect 12437 10180 12449 10183
rect 12400 10152 12449 10180
rect 12400 10140 12406 10152
rect 12437 10149 12449 10152
rect 12483 10180 12495 10183
rect 12986 10180 12992 10192
rect 12483 10152 12992 10180
rect 12483 10149 12495 10152
rect 12437 10143 12495 10149
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 10965 10115 11023 10121
rect 10965 10112 10977 10115
rect 10796 10084 10977 10112
rect 6181 10007 6239 10013
rect 8956 10016 9536 10044
rect 9968 10016 10456 10044
rect 3252 9880 5580 9908
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 7561 9911 7619 9917
rect 7561 9877 7573 9911
rect 7607 9908 7619 9911
rect 8956 9908 8984 10016
rect 9968 9976 9996 10016
rect 9048 9948 9996 9976
rect 10045 9979 10103 9985
rect 9048 9917 9076 9948
rect 10045 9945 10057 9979
rect 10091 9976 10103 9979
rect 10796 9976 10824 10084
rect 10965 10081 10977 10084
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10081 11115 10115
rect 11057 10075 11115 10081
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 11572 10084 12081 10112
rect 11572 10072 11578 10084
rect 12069 10081 12081 10084
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10112 12679 10115
rect 13096 10112 13124 10220
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 14240 10220 14381 10248
rect 14240 10208 14246 10220
rect 14369 10217 14381 10220
rect 14415 10248 14427 10251
rect 14550 10248 14556 10260
rect 14415 10220 14556 10248
rect 14415 10217 14427 10220
rect 14369 10211 14427 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15197 10251 15255 10257
rect 15197 10217 15209 10251
rect 15243 10248 15255 10251
rect 15378 10248 15384 10260
rect 15243 10220 15384 10248
rect 15243 10217 15255 10220
rect 15197 10211 15255 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 15562 10208 15568 10260
rect 15620 10208 15626 10260
rect 16390 10208 16396 10260
rect 16448 10208 16454 10260
rect 17589 10251 17647 10257
rect 17589 10217 17601 10251
rect 17635 10248 17647 10251
rect 18049 10251 18107 10257
rect 18049 10248 18061 10251
rect 17635 10220 18061 10248
rect 17635 10217 17647 10220
rect 17589 10211 17647 10217
rect 18049 10217 18061 10220
rect 18095 10217 18107 10251
rect 18049 10211 18107 10217
rect 19429 10251 19487 10257
rect 19429 10217 19441 10251
rect 19475 10248 19487 10251
rect 20070 10248 20076 10260
rect 19475 10220 20076 10248
rect 19475 10217 19487 10220
rect 19429 10211 19487 10217
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20346 10208 20352 10260
rect 20404 10208 20410 10260
rect 20898 10208 20904 10260
rect 20956 10208 20962 10260
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21232 10220 21680 10248
rect 21232 10208 21238 10220
rect 13998 10140 14004 10192
rect 14056 10180 14062 10192
rect 14093 10183 14151 10189
rect 14093 10180 14105 10183
rect 14056 10152 14105 10180
rect 14056 10140 14062 10152
rect 14093 10149 14105 10152
rect 14139 10180 14151 10183
rect 15580 10180 15608 10208
rect 14139 10152 15608 10180
rect 14139 10149 14151 10152
rect 14093 10143 14151 10149
rect 14274 10112 14280 10124
rect 12667 10084 14280 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 12084 10044 12112 10075
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 14921 10115 14979 10121
rect 14921 10112 14933 10115
rect 14792 10084 14933 10112
rect 14792 10072 14798 10084
rect 14921 10081 14933 10084
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 16206 10072 16212 10124
rect 16264 10072 16270 10124
rect 16408 10112 16436 10208
rect 19638 10183 19696 10189
rect 19638 10180 19650 10183
rect 19444 10152 19650 10180
rect 19444 10124 19472 10152
rect 19638 10149 19650 10152
rect 19684 10149 19696 10183
rect 19638 10143 19696 10149
rect 16465 10115 16523 10121
rect 16465 10112 16477 10115
rect 16408 10084 16477 10112
rect 16465 10081 16477 10084
rect 16511 10081 16523 10115
rect 16465 10075 16523 10081
rect 19426 10072 19432 10124
rect 19484 10072 19490 10124
rect 14829 10047 14887 10053
rect 12084 10016 14320 10044
rect 10091 9948 10824 9976
rect 10091 9945 10103 9948
rect 10045 9939 10103 9945
rect 10870 9936 10876 9988
rect 10928 9976 10934 9988
rect 11333 9979 11391 9985
rect 11333 9976 11345 9979
rect 10928 9948 11345 9976
rect 10928 9936 10934 9948
rect 11333 9945 11345 9948
rect 11379 9945 11391 9979
rect 11333 9939 11391 9945
rect 7607 9880 8984 9908
rect 9033 9911 9091 9917
rect 7607 9877 7619 9880
rect 7561 9871 7619 9877
rect 9033 9877 9045 9911
rect 9079 9877 9091 9911
rect 9033 9871 9091 9877
rect 10689 9911 10747 9917
rect 10689 9877 10701 9911
rect 10735 9908 10747 9911
rect 10965 9911 11023 9917
rect 10965 9908 10977 9911
rect 10735 9880 10977 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 10965 9877 10977 9880
rect 11011 9877 11023 9911
rect 10965 9871 11023 9877
rect 12710 9868 12716 9920
rect 12768 9868 12774 9920
rect 14292 9908 14320 10016
rect 14829 10013 14841 10047
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 14844 9976 14872 10007
rect 15010 10004 15016 10056
rect 15068 10004 15074 10056
rect 18138 10004 18144 10056
rect 18196 10004 18202 10056
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 18966 10004 18972 10056
rect 19024 10004 19030 10056
rect 19150 10004 19156 10056
rect 19208 10004 19214 10056
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10013 19579 10047
rect 19521 10007 19579 10013
rect 16206 9976 16212 9988
rect 14844 9948 16212 9976
rect 16206 9936 16212 9948
rect 16264 9936 16270 9988
rect 18984 9976 19012 10004
rect 19536 9976 19564 10007
rect 18984 9948 19564 9976
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9976 19855 9979
rect 19978 9976 19984 9988
rect 19843 9948 19984 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 16390 9908 16396 9920
rect 14292 9880 16396 9908
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 17681 9911 17739 9917
rect 17681 9908 17693 9911
rect 16632 9880 17693 9908
rect 16632 9868 16638 9880
rect 17681 9877 17693 9880
rect 17727 9877 17739 9911
rect 20364 9908 20392 10208
rect 20916 10180 20944 10208
rect 21514 10183 21572 10189
rect 21514 10180 21526 10183
rect 20916 10152 21526 10180
rect 21514 10149 21526 10152
rect 21560 10149 21572 10183
rect 21514 10143 21572 10149
rect 20714 10072 20720 10124
rect 20772 10072 20778 10124
rect 20901 10115 20959 10121
rect 20901 10081 20913 10115
rect 20947 10112 20959 10115
rect 21358 10112 21364 10124
rect 20947 10084 21364 10112
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 21652 10112 21680 10220
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22649 10251 22707 10257
rect 22649 10248 22661 10251
rect 22244 10220 22661 10248
rect 22244 10208 22250 10220
rect 22649 10217 22661 10220
rect 22695 10217 22707 10251
rect 22649 10211 22707 10217
rect 23032 10220 23980 10248
rect 22278 10140 22284 10192
rect 22336 10180 22342 10192
rect 23032 10180 23060 10220
rect 22336 10152 23060 10180
rect 22336 10140 22342 10152
rect 22646 10112 22652 10124
rect 21652 10084 22652 10112
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 23106 10072 23112 10124
rect 23164 10072 23170 10124
rect 23382 10121 23388 10124
rect 23376 10075 23388 10121
rect 23382 10072 23388 10075
rect 23440 10072 23446 10124
rect 23952 10112 23980 10220
rect 25222 10180 25228 10192
rect 24688 10152 25228 10180
rect 24688 10121 24716 10152
rect 25222 10140 25228 10152
rect 25280 10140 25286 10192
rect 26620 10152 27752 10180
rect 24673 10115 24731 10121
rect 24673 10112 24685 10115
rect 23952 10084 24685 10112
rect 24673 10081 24685 10084
rect 24719 10081 24731 10115
rect 24673 10075 24731 10081
rect 24854 10072 24860 10124
rect 24912 10072 24918 10124
rect 25406 10072 25412 10124
rect 25464 10072 25470 10124
rect 25590 10072 25596 10124
rect 25648 10072 25654 10124
rect 26620 10121 26648 10152
rect 26878 10121 26884 10124
rect 26605 10115 26663 10121
rect 26605 10081 26617 10115
rect 26651 10081 26663 10115
rect 26605 10075 26663 10081
rect 26872 10075 26884 10121
rect 21174 10004 21180 10056
rect 21232 10044 21238 10056
rect 21269 10047 21327 10053
rect 21269 10044 21281 10047
rect 21232 10016 21281 10044
rect 21232 10004 21238 10016
rect 21269 10013 21281 10016
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 24394 10004 24400 10056
rect 24452 10004 24458 10056
rect 24412 9976 24440 10004
rect 26620 9976 26648 10075
rect 26878 10072 26884 10075
rect 26936 10072 26942 10124
rect 27724 10044 27752 10152
rect 27890 10072 27896 10124
rect 27948 10112 27954 10124
rect 28333 10115 28391 10121
rect 28333 10112 28345 10115
rect 27948 10084 28345 10112
rect 27948 10072 27954 10084
rect 28333 10081 28345 10084
rect 28379 10081 28391 10115
rect 28333 10075 28391 10081
rect 27982 10044 27988 10056
rect 27724 10016 27988 10044
rect 27982 10004 27988 10016
rect 28040 10044 28046 10056
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 28040 10016 28089 10044
rect 28040 10004 28046 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 24412 9948 26648 9976
rect 20717 9911 20775 9917
rect 20717 9908 20729 9911
rect 20364 9880 20729 9908
rect 17681 9871 17739 9877
rect 20717 9877 20729 9880
rect 20763 9877 20775 9911
rect 20717 9871 20775 9877
rect 21085 9911 21143 9917
rect 21085 9877 21097 9911
rect 21131 9908 21143 9911
rect 22278 9908 22284 9920
rect 21131 9880 22284 9908
rect 21131 9877 21143 9880
rect 21085 9871 21143 9877
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 24489 9911 24547 9917
rect 24489 9877 24501 9911
rect 24535 9908 24547 9911
rect 24670 9908 24676 9920
rect 24535 9880 24676 9908
rect 24535 9877 24547 9880
rect 24489 9871 24547 9877
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 25866 9868 25872 9920
rect 25924 9868 25930 9920
rect 27982 9868 27988 9920
rect 28040 9868 28046 9920
rect 29454 9868 29460 9920
rect 29512 9868 29518 9920
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 9766 9704 9772 9716
rect 6380 9676 6592 9704
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 3252 9568 3280 9596
rect 4893 9571 4951 9577
rect 3252 9540 3372 9568
rect 3234 9460 3240 9512
rect 3292 9460 3298 9512
rect 3344 9500 3372 9540
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5905 9571 5963 9577
rect 5905 9568 5917 9571
rect 4939 9540 5917 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 5905 9537 5917 9540
rect 5951 9568 5963 9571
rect 6380 9568 6408 9676
rect 6457 9639 6515 9645
rect 6457 9605 6469 9639
rect 6503 9605 6515 9639
rect 6564 9636 6592 9676
rect 9232 9676 9772 9704
rect 9232 9636 9260 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 13998 9704 14004 9716
rect 9916 9676 14004 9704
rect 9916 9664 9922 9676
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 18049 9707 18107 9713
rect 16684 9676 17632 9704
rect 6564 9608 9260 9636
rect 9309 9639 9367 9645
rect 6457 9599 6515 9605
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 10594 9636 10600 9648
rect 9355 9608 10600 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 5951 9540 6408 9568
rect 6472 9568 6500 9599
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 11330 9636 11336 9648
rect 10796 9608 11336 9636
rect 10796 9577 10824 9608
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 16209 9639 16267 9645
rect 16209 9636 16221 9639
rect 15712 9608 16221 9636
rect 15712 9596 15718 9608
rect 16209 9605 16221 9608
rect 16255 9605 16267 9639
rect 16209 9599 16267 9605
rect 10781 9571 10839 9577
rect 6472 9540 10732 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 3493 9503 3551 9509
rect 3493 9500 3505 9503
rect 3344 9472 3505 9500
rect 3493 9469 3505 9472
rect 3539 9469 3551 9503
rect 3493 9463 3551 9469
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5684 9472 6101 9500
rect 5684 9460 5690 9472
rect 6089 9469 6101 9472
rect 6135 9469 6147 9503
rect 6089 9463 6147 9469
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 9416 9472 9996 9500
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4632 9404 5089 9432
rect 4632 9373 4660 9404
rect 5077 9401 5089 9404
rect 5123 9401 5135 9435
rect 9416 9432 9444 9472
rect 5077 9395 5135 9401
rect 5460 9404 9444 9432
rect 9585 9435 9643 9441
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9333 4675 9367
rect 4617 9327 4675 9333
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5460 9373 5488 9404
rect 9585 9401 9597 9435
rect 9631 9401 9643 9435
rect 9968 9432 9996 9472
rect 10042 9460 10048 9512
rect 10100 9460 10106 9512
rect 10704 9509 10732 9540
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10870 9528 10876 9580
rect 10928 9568 10934 9580
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10928 9540 10977 9568
rect 10928 9528 10934 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 12952 9540 14013 9568
rect 12952 9528 12958 9540
rect 14001 9537 14013 9540
rect 14047 9568 14059 9571
rect 15749 9571 15807 9577
rect 15749 9568 15761 9571
rect 14047 9540 15761 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 15749 9537 15761 9540
rect 15795 9568 15807 9571
rect 16684 9568 16712 9676
rect 17604 9636 17632 9676
rect 18049 9673 18061 9707
rect 18095 9704 18107 9707
rect 18138 9704 18144 9716
rect 18095 9676 18144 9704
rect 18095 9673 18107 9676
rect 18049 9667 18107 9673
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 20456 9676 20668 9704
rect 20456 9636 20484 9676
rect 17604 9608 20484 9636
rect 20533 9639 20591 9645
rect 20533 9605 20545 9639
rect 20579 9605 20591 9639
rect 20640 9636 20668 9676
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 21453 9707 21511 9713
rect 21453 9704 21465 9707
rect 20772 9676 21465 9704
rect 20772 9664 20778 9676
rect 21453 9673 21465 9676
rect 21499 9673 21511 9707
rect 23293 9707 23351 9713
rect 21453 9667 21511 9673
rect 21652 9676 22692 9704
rect 20898 9636 20904 9648
rect 20640 9608 20904 9636
rect 20533 9599 20591 9605
rect 15795 9540 16712 9568
rect 18984 9540 20024 9568
rect 15795 9537 15807 9540
rect 15749 9531 15807 9537
rect 18984 9512 19012 9540
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9469 10747 9503
rect 10689 9463 10747 9469
rect 11054 9460 11060 9512
rect 11112 9460 11118 9512
rect 11514 9460 11520 9512
rect 11572 9500 11578 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11572 9472 11621 9500
rect 11572 9460 11578 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 11609 9463 11667 9469
rect 11716 9472 14197 9500
rect 11716 9432 11744 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14550 9460 14556 9512
rect 14608 9460 14614 9512
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 15378 9460 15384 9512
rect 15436 9460 15442 9512
rect 15470 9460 15476 9512
rect 15528 9460 15534 9512
rect 15841 9503 15899 9509
rect 15841 9469 15853 9503
rect 15887 9500 15899 9503
rect 16574 9500 16580 9512
rect 15887 9472 16580 9500
rect 15887 9469 15899 9472
rect 15841 9463 15899 9469
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9500 16727 9503
rect 17494 9500 17500 9512
rect 16715 9472 17500 9500
rect 16715 9469 16727 9472
rect 16669 9463 16727 9469
rect 17494 9460 17500 9472
rect 17552 9500 17558 9512
rect 18598 9500 18604 9512
rect 17552 9472 18604 9500
rect 17552 9460 17558 9472
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 18966 9460 18972 9512
rect 19024 9460 19030 9512
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9469 19947 9503
rect 19996 9500 20024 9540
rect 20162 9528 20168 9580
rect 20220 9568 20226 9580
rect 20374 9571 20432 9577
rect 20374 9568 20386 9571
rect 20220 9540 20386 9568
rect 20220 9528 20226 9540
rect 20374 9537 20386 9540
rect 20420 9537 20432 9571
rect 20548 9568 20576 9599
rect 20898 9596 20904 9608
rect 20956 9636 20962 9648
rect 21652 9636 21680 9676
rect 22664 9636 22692 9676
rect 23293 9673 23305 9707
rect 23339 9704 23351 9707
rect 23382 9704 23388 9716
rect 23339 9676 23388 9704
rect 23339 9673 23351 9676
rect 23293 9667 23351 9673
rect 23382 9664 23388 9676
rect 23440 9664 23446 9716
rect 24857 9707 24915 9713
rect 24857 9673 24869 9707
rect 24903 9704 24915 9707
rect 25406 9704 25412 9716
rect 24903 9676 25412 9704
rect 24903 9673 24915 9676
rect 24857 9667 24915 9673
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 26145 9707 26203 9713
rect 26145 9673 26157 9707
rect 26191 9673 26203 9707
rect 26145 9667 26203 9673
rect 26329 9707 26387 9713
rect 26329 9673 26341 9707
rect 26375 9704 26387 9707
rect 26694 9704 26700 9716
rect 26375 9676 26700 9704
rect 26375 9673 26387 9676
rect 26329 9667 26387 9673
rect 24578 9636 24584 9648
rect 20956 9608 21680 9636
rect 21836 9608 22600 9636
rect 22664 9608 24584 9636
rect 20956 9596 20962 9608
rect 21726 9568 21732 9580
rect 20548 9540 21732 9568
rect 20374 9531 20432 9537
rect 21726 9528 21732 9540
rect 21784 9528 21790 9580
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 19996 9472 20269 9500
rect 19889 9463 19947 9469
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 21637 9503 21695 9509
rect 21637 9469 21649 9503
rect 21683 9500 21695 9503
rect 21836 9500 21864 9608
rect 21910 9528 21916 9580
rect 21968 9528 21974 9580
rect 22186 9568 22192 9580
rect 22112 9540 22192 9568
rect 21683 9472 21864 9500
rect 21928 9500 21956 9528
rect 22112 9509 22140 9540
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 22572 9577 22600 9608
rect 24578 9596 24584 9608
rect 24636 9636 24642 9648
rect 25774 9636 25780 9648
rect 24636 9608 25780 9636
rect 24636 9596 24642 9608
rect 25774 9596 25780 9608
rect 25832 9596 25838 9648
rect 26160 9636 26188 9667
rect 26694 9664 26700 9676
rect 26752 9664 26758 9716
rect 26789 9707 26847 9713
rect 26789 9673 26801 9707
rect 26835 9704 26847 9707
rect 26878 9704 26884 9716
rect 26835 9676 26884 9704
rect 26835 9673 26847 9676
rect 26789 9667 26847 9673
rect 26878 9664 26884 9676
rect 26936 9664 26942 9716
rect 27062 9664 27068 9716
rect 27120 9704 27126 9716
rect 27249 9707 27307 9713
rect 27249 9704 27261 9707
rect 27120 9676 27261 9704
rect 27120 9664 27126 9676
rect 27249 9673 27261 9676
rect 27295 9673 27307 9707
rect 27249 9667 27307 9673
rect 27617 9707 27675 9713
rect 27617 9673 27629 9707
rect 27663 9704 27675 9707
rect 27890 9704 27896 9716
rect 27663 9676 27896 9704
rect 27663 9673 27675 9676
rect 27617 9667 27675 9673
rect 27890 9664 27896 9676
rect 27948 9664 27954 9716
rect 27982 9664 27988 9716
rect 28040 9704 28046 9716
rect 28040 9676 29592 9704
rect 28040 9664 28046 9676
rect 28997 9639 29055 9645
rect 28997 9636 29009 9639
rect 26160 9608 29009 9636
rect 28997 9605 29009 9608
rect 29043 9605 29055 9639
rect 28997 9599 29055 9605
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9537 22339 9571
rect 22281 9531 22339 9537
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9537 22615 9571
rect 22557 9531 22615 9537
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 24302 9568 24308 9580
rect 22787 9540 24308 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 21928 9472 22017 9500
rect 21683 9469 21695 9472
rect 21637 9463 21695 9469
rect 22005 9469 22017 9472
rect 22051 9469 22063 9503
rect 22005 9463 22063 9469
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 9968 9404 11744 9432
rect 11876 9435 11934 9441
rect 9585 9395 9643 9401
rect 11876 9401 11888 9435
rect 11922 9432 11934 9435
rect 12250 9432 12256 9444
rect 11922 9404 12256 9432
rect 11922 9401 11934 9404
rect 11876 9395 11934 9401
rect 4985 9367 5043 9373
rect 4985 9364 4997 9367
rect 4856 9336 4997 9364
rect 4856 9324 4862 9336
rect 4985 9333 4997 9336
rect 5031 9333 5043 9367
rect 4985 9327 5043 9333
rect 5445 9367 5503 9373
rect 5445 9333 5457 9367
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 5994 9324 6000 9376
rect 6052 9324 6058 9376
rect 7282 9324 7288 9376
rect 7340 9324 7346 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9600 9364 9628 9395
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 16936 9435 16994 9441
rect 16936 9401 16948 9435
rect 16982 9432 16994 9435
rect 17678 9432 17684 9444
rect 16982 9404 17684 9432
rect 16982 9401 16994 9404
rect 16936 9395 16994 9401
rect 17678 9392 17684 9404
rect 17736 9392 17742 9444
rect 18414 9392 18420 9444
rect 18472 9432 18478 9444
rect 19150 9432 19156 9444
rect 18472 9404 19156 9432
rect 18472 9392 18478 9404
rect 19150 9392 19156 9404
rect 19208 9432 19214 9444
rect 19904 9432 19932 9463
rect 19208 9404 19932 9432
rect 19208 9392 19214 9404
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 21652 9432 21680 9463
rect 20036 9404 21680 9432
rect 21731 9435 21789 9441
rect 20036 9392 20042 9404
rect 21731 9401 21743 9435
rect 21777 9401 21789 9435
rect 21731 9395 21789 9401
rect 9272 9336 9628 9364
rect 9272 9324 9278 9336
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 9824 9336 9873 9364
rect 9824 9324 9830 9336
rect 9861 9333 9873 9336
rect 9907 9364 9919 9367
rect 10962 9364 10968 9376
rect 9907 9336 10968 9364
rect 9907 9333 9919 9336
rect 9861 9327 9919 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 12894 9364 12900 9376
rect 11388 9336 12900 9364
rect 11388 9324 11394 9336
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 12989 9367 13047 9373
rect 12989 9333 13001 9367
rect 13035 9364 13047 9367
rect 13078 9364 13084 9376
rect 13035 9336 13084 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 13630 9324 13636 9376
rect 13688 9324 13694 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 16758 9364 16764 9376
rect 14792 9336 16764 9364
rect 14792 9324 14798 9336
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 19484 9336 20177 9364
rect 19484 9324 19490 9336
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20165 9327 20223 9333
rect 20622 9324 20628 9376
rect 20680 9364 20686 9376
rect 21749 9364 21777 9395
rect 21818 9392 21824 9444
rect 21876 9392 21882 9444
rect 22186 9392 22192 9444
rect 22244 9432 22250 9444
rect 22296 9432 22324 9531
rect 24302 9528 24308 9540
rect 24360 9528 24366 9580
rect 27338 9568 27344 9580
rect 27080 9540 27344 9568
rect 22370 9460 22376 9512
rect 22428 9460 22434 9512
rect 22462 9460 22468 9512
rect 22520 9460 22526 9512
rect 23014 9460 23020 9512
rect 23072 9500 23078 9512
rect 23109 9503 23167 9509
rect 23109 9500 23121 9503
rect 23072 9472 23121 9500
rect 23072 9460 23078 9472
rect 23109 9469 23121 9472
rect 23155 9469 23167 9503
rect 23109 9463 23167 9469
rect 24486 9460 24492 9512
rect 24544 9460 24550 9512
rect 24578 9460 24584 9512
rect 24636 9460 24642 9512
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9500 24915 9503
rect 25130 9500 25136 9512
rect 24903 9472 25136 9500
rect 24903 9469 24915 9472
rect 24857 9463 24915 9469
rect 22244 9404 24440 9432
rect 22244 9392 22250 9404
rect 22462 9364 22468 9376
rect 20680 9336 22468 9364
rect 20680 9324 20686 9336
rect 22462 9324 22468 9336
rect 22520 9324 22526 9376
rect 24118 9324 24124 9376
rect 24176 9364 24182 9376
rect 24305 9367 24363 9373
rect 24305 9364 24317 9367
rect 24176 9336 24317 9364
rect 24176 9324 24182 9336
rect 24305 9333 24317 9336
rect 24351 9333 24363 9367
rect 24412 9364 24440 9404
rect 24670 9392 24676 9444
rect 24728 9392 24734 9444
rect 24872 9364 24900 9463
rect 25130 9460 25136 9472
rect 25188 9460 25194 9512
rect 25958 9460 25964 9512
rect 26016 9460 26022 9512
rect 26050 9460 26056 9512
rect 26108 9460 26114 9512
rect 26878 9460 26884 9512
rect 26936 9500 26942 9512
rect 27080 9509 27108 9540
rect 27338 9528 27344 9540
rect 27396 9568 27402 9580
rect 27396 9540 27936 9568
rect 27396 9528 27402 9540
rect 26973 9503 27031 9509
rect 26973 9500 26985 9503
rect 26936 9472 26985 9500
rect 26936 9460 26942 9472
rect 26973 9469 26985 9472
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 27065 9503 27123 9509
rect 27065 9469 27077 9503
rect 27111 9469 27123 9503
rect 27249 9503 27307 9509
rect 27249 9500 27261 9503
rect 27065 9463 27123 9469
rect 27172 9472 27261 9500
rect 24412 9336 24900 9364
rect 24305 9327 24363 9333
rect 26970 9324 26976 9376
rect 27028 9364 27034 9376
rect 27172 9364 27200 9472
rect 27249 9469 27261 9472
rect 27295 9469 27307 9503
rect 27249 9463 27307 9469
rect 27430 9460 27436 9512
rect 27488 9460 27494 9512
rect 27798 9460 27804 9512
rect 27856 9460 27862 9512
rect 27908 9509 27936 9540
rect 27893 9503 27951 9509
rect 27893 9469 27905 9503
rect 27939 9469 27951 9503
rect 27893 9463 27951 9469
rect 28074 9460 28080 9512
rect 28132 9500 28138 9512
rect 29178 9500 29184 9512
rect 28132 9472 29184 9500
rect 28132 9460 28138 9472
rect 29178 9460 29184 9472
rect 29236 9460 29242 9512
rect 29273 9503 29331 9509
rect 29273 9469 29285 9503
rect 29319 9500 29331 9503
rect 29454 9500 29460 9512
rect 29319 9472 29460 9500
rect 29319 9469 29331 9472
rect 29273 9463 29331 9469
rect 29454 9460 29460 9472
rect 29512 9460 29518 9512
rect 29564 9509 29592 9676
rect 29549 9503 29607 9509
rect 29549 9469 29561 9503
rect 29595 9469 29607 9503
rect 29549 9463 29607 9469
rect 27816 9432 27844 9460
rect 29362 9432 29368 9444
rect 27816 9404 29368 9432
rect 29362 9392 29368 9404
rect 29420 9392 29426 9444
rect 27028 9336 27200 9364
rect 27028 9324 27034 9336
rect 28074 9324 28080 9376
rect 28132 9324 28138 9376
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 5994 9160 6000 9172
rect 5675 9132 6000 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7282 9160 7288 9172
rect 6963 9132 7288 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 8665 9163 8723 9169
rect 8665 9129 8677 9163
rect 8711 9160 8723 9163
rect 11330 9160 11336 9172
rect 8711 9132 11336 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 13909 9163 13967 9169
rect 11992 9132 13308 9160
rect 7098 9092 7104 9104
rect 6748 9064 7104 9092
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 3605 9027 3663 9033
rect 3605 9024 3617 9027
rect 3292 8996 3617 9024
rect 3292 8984 3298 8996
rect 3605 8993 3617 8996
rect 3651 8993 3663 9027
rect 3605 8987 3663 8993
rect 4516 9027 4574 9033
rect 4516 8993 4528 9027
rect 4562 9024 4574 9027
rect 4982 9024 4988 9036
rect 4562 8996 4988 9024
rect 4562 8993 4574 8996
rect 4516 8987 4574 8993
rect 3620 8956 3648 8987
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 6748 9033 6776 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 7190 9052 7196 9104
rect 7248 9052 7254 9104
rect 7300 9092 7328 9120
rect 7530 9095 7588 9101
rect 7530 9092 7542 9095
rect 7300 9064 7542 9092
rect 7530 9061 7542 9064
rect 7576 9061 7588 9095
rect 7530 9055 7588 9061
rect 10410 9052 10416 9104
rect 10468 9052 10474 9104
rect 11057 9095 11115 9101
rect 11057 9061 11069 9095
rect 11103 9092 11115 9095
rect 11146 9092 11152 9104
rect 11103 9064 11152 9092
rect 11103 9061 11115 9064
rect 11057 9055 11115 9061
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 11238 9052 11244 9104
rect 11296 9092 11302 9104
rect 11425 9095 11483 9101
rect 11425 9092 11437 9095
rect 11296 9064 11437 9092
rect 11296 9052 11302 9064
rect 11425 9061 11437 9064
rect 11471 9061 11483 9095
rect 11425 9055 11483 9061
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 11885 9095 11943 9101
rect 11885 9092 11897 9095
rect 11664 9064 11897 9092
rect 11664 9052 11670 9064
rect 11885 9061 11897 9064
rect 11931 9061 11943 9095
rect 11885 9055 11943 9061
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 8993 6791 9027
rect 7208 9024 7236 9052
rect 7285 9027 7343 9033
rect 7285 9024 7297 9027
rect 7208 8996 7297 9024
rect 6733 8987 6791 8993
rect 7285 8993 7297 8996
rect 7331 8993 7343 9027
rect 7285 8987 7343 8993
rect 9585 9027 9643 9033
rect 9585 8993 9597 9027
rect 9631 9024 9643 9027
rect 9950 9024 9956 9036
rect 9631 8996 9956 9024
rect 9631 8993 9643 8996
rect 9585 8987 9643 8993
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10134 9024 10140 9036
rect 10091 8996 10140 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 11164 9024 11192 9052
rect 11992 9024 12020 9132
rect 13078 9052 13084 9104
rect 13136 9052 13142 9104
rect 13280 9036 13308 9132
rect 13909 9129 13921 9163
rect 13955 9160 13967 9163
rect 14550 9160 14556 9172
rect 13955 9132 14556 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 14921 9163 14979 9169
rect 14921 9129 14933 9163
rect 14967 9160 14979 9163
rect 15102 9160 15108 9172
rect 14967 9132 15108 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 16482 9120 16488 9172
rect 16540 9120 16546 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 16945 9163 17003 9169
rect 16945 9129 16957 9163
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 14185 9095 14243 9101
rect 14185 9061 14197 9095
rect 14231 9092 14243 9095
rect 15838 9092 15844 9104
rect 14231 9064 15844 9092
rect 14231 9061 14243 9064
rect 14185 9055 14243 9061
rect 11164 8996 12020 9024
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 9024 12311 9027
rect 12342 9024 12348 9036
rect 12299 8996 12348 9024
rect 12299 8993 12311 8996
rect 12253 8987 12311 8993
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12526 8984 12532 9036
rect 12584 8984 12590 9036
rect 12802 8984 12808 9036
rect 12860 8984 12866 9036
rect 12986 8984 12992 9036
rect 13044 8984 13050 9036
rect 13262 9033 13268 9036
rect 13219 9027 13268 9033
rect 13219 8993 13231 9027
rect 13265 8993 13268 9027
rect 13219 8987 13268 8993
rect 13262 8984 13268 8987
rect 13320 8984 13326 9036
rect 13538 8984 13544 9036
rect 13596 8984 13602 9036
rect 13722 8984 13728 9036
rect 13780 8984 13786 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14366 9024 14372 9036
rect 13872 8996 14372 9024
rect 13872 8984 13878 8996
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14553 9027 14611 9033
rect 14734 9028 14740 9036
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 14660 9024 14740 9028
rect 14599 9000 14740 9024
rect 14599 8996 14688 9000
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 14734 8984 14740 9000
rect 14792 8984 14798 9036
rect 14936 9033 14964 9064
rect 15838 9052 15844 9064
rect 15896 9092 15902 9104
rect 16960 9092 16988 9123
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17494 9160 17500 9172
rect 17184 9132 17500 9160
rect 17184 9120 17190 9132
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 17678 9120 17684 9172
rect 17736 9120 17742 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19794 9160 19800 9172
rect 19392 9132 19800 9160
rect 19392 9120 19398 9132
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 19889 9163 19947 9169
rect 19889 9129 19901 9163
rect 19935 9160 19947 9163
rect 19978 9160 19984 9172
rect 19935 9132 19984 9160
rect 19935 9129 19947 9132
rect 19889 9123 19947 9129
rect 19978 9120 19984 9132
rect 20036 9160 20042 9172
rect 20622 9160 20628 9172
rect 20036 9132 20628 9160
rect 20036 9120 20042 9132
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22428 9132 22661 9160
rect 22428 9120 22434 9132
rect 22649 9129 22661 9132
rect 22695 9129 22707 9163
rect 22649 9123 22707 9129
rect 24029 9163 24087 9169
rect 24029 9129 24041 9163
rect 24075 9129 24087 9163
rect 24029 9123 24087 9129
rect 25501 9163 25559 9169
rect 25501 9129 25513 9163
rect 25547 9160 25559 9163
rect 25961 9163 26019 9169
rect 25961 9160 25973 9163
rect 25547 9132 25973 9160
rect 25547 9129 25559 9132
rect 25501 9123 25559 9129
rect 25961 9129 25973 9132
rect 26007 9129 26019 9163
rect 25961 9123 26019 9129
rect 15896 9064 16988 9092
rect 15896 9052 15902 9064
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 8993 14979 9027
rect 14921 8987 14979 8993
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 15470 9024 15476 9036
rect 15068 8996 15476 9024
rect 15068 8984 15074 8996
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 16132 9033 16160 9064
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16853 9027 16911 9033
rect 16853 9024 16865 9027
rect 16264 8996 16865 9024
rect 16264 8984 16270 8996
rect 16853 8993 16865 8996
rect 16899 8993 16911 9027
rect 16960 9024 16988 9064
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 24044 9092 24072 9123
rect 26326 9120 26332 9172
rect 26384 9160 26390 9172
rect 29917 9163 29975 9169
rect 29917 9160 29929 9163
rect 26384 9132 29929 9160
rect 26384 9120 26390 9132
rect 29917 9129 29929 9132
rect 29963 9129 29975 9163
rect 29917 9123 29975 9129
rect 24366 9095 24424 9101
rect 24366 9092 24378 9095
rect 17092 9064 23980 9092
rect 24044 9064 24378 9092
rect 17092 9052 17098 9064
rect 17313 9027 17371 9033
rect 16960 8996 17264 9024
rect 16853 8987 16911 8993
rect 4062 8956 4068 8968
rect 3620 8928 4068 8956
rect 4062 8916 4068 8928
rect 4120 8956 4126 8968
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 4120 8928 4261 8956
rect 4120 8916 4126 8928
rect 4249 8925 4261 8928
rect 4295 8925 4307 8959
rect 10152 8956 10180 8984
rect 17236 8956 17264 8996
rect 17313 8993 17325 9027
rect 17359 9024 17371 9027
rect 17586 9024 17592 9036
rect 17359 8996 17592 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 17865 9027 17923 9033
rect 17865 9024 17877 9027
rect 17828 8996 17877 9024
rect 17828 8984 17834 8996
rect 17865 8993 17877 8996
rect 17911 8993 17923 9027
rect 17865 8987 17923 8993
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 18509 9027 18567 9033
rect 18509 9024 18521 9027
rect 18380 8996 18521 9024
rect 18380 8984 18386 8996
rect 18509 8993 18521 8996
rect 18555 8993 18567 9027
rect 18509 8987 18567 8993
rect 18414 8956 18420 8968
rect 10152 8928 13768 8956
rect 4249 8919 4307 8925
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 5776 8860 7328 8888
rect 5776 8848 5782 8860
rect 7300 8832 7328 8860
rect 8220 8860 11928 8888
rect 7190 8780 7196 8832
rect 7248 8780 7254 8832
rect 7282 8780 7288 8832
rect 7340 8780 7346 8832
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 8220 8820 8248 8860
rect 7984 8792 8248 8820
rect 7984 8780 7990 8792
rect 9398 8780 9404 8832
rect 9456 8780 9462 8832
rect 11514 8780 11520 8832
rect 11572 8820 11578 8832
rect 11793 8823 11851 8829
rect 11793 8820 11805 8823
rect 11572 8792 11805 8820
rect 11572 8780 11578 8792
rect 11793 8789 11805 8792
rect 11839 8789 11851 8823
rect 11900 8820 11928 8860
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 12345 8891 12403 8897
rect 12345 8888 12357 8891
rect 12308 8860 12357 8888
rect 12308 8848 12314 8860
rect 12345 8857 12357 8860
rect 12391 8857 12403 8891
rect 13740 8888 13768 8928
rect 14108 8928 16988 8956
rect 17236 8928 18420 8956
rect 13814 8888 13820 8900
rect 12345 8851 12403 8857
rect 13280 8860 13676 8888
rect 13740 8860 13820 8888
rect 13280 8820 13308 8860
rect 11900 8792 13308 8820
rect 13357 8823 13415 8829
rect 11793 8783 11851 8789
rect 13357 8789 13369 8823
rect 13403 8820 13415 8823
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13403 8792 13553 8820
rect 13403 8789 13415 8792
rect 13357 8783 13415 8789
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13648 8820 13676 8860
rect 13814 8848 13820 8860
rect 13872 8888 13878 8900
rect 14001 8891 14059 8897
rect 14001 8888 14013 8891
rect 13872 8860 14013 8888
rect 13872 8848 13878 8860
rect 14001 8857 14013 8860
rect 14047 8857 14059 8891
rect 14001 8851 14059 8857
rect 14108 8820 14136 8928
rect 16960 8888 16988 8928
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 18524 8956 18552 8987
rect 18598 8984 18604 9036
rect 18656 9024 18662 9036
rect 18656 8996 19334 9024
rect 18656 8984 18662 8996
rect 18966 8956 18972 8968
rect 18524 8928 18972 8956
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 19306 8956 19334 8996
rect 19426 8984 19432 9036
rect 19484 8984 19490 9036
rect 20070 8984 20076 9036
rect 20128 8984 20134 9036
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 9024 20407 9027
rect 20898 9024 20904 9036
rect 20395 8996 20904 9024
rect 20395 8993 20407 8996
rect 20349 8987 20407 8993
rect 20898 8984 20904 8996
rect 20956 8984 20962 9036
rect 21174 8984 21180 9036
rect 21232 9024 21238 9036
rect 21525 9027 21583 9033
rect 21525 9024 21537 9027
rect 21232 8996 21537 9024
rect 21232 8984 21238 8996
rect 21525 8993 21537 8996
rect 21571 8993 21583 9027
rect 21525 8987 21583 8993
rect 23014 8984 23020 9036
rect 23072 8984 23078 9036
rect 23106 8984 23112 9036
rect 23164 8984 23170 9036
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 8993 23903 9027
rect 23952 9024 23980 9064
rect 24366 9061 24378 9064
rect 24412 9061 24424 9095
rect 24366 9055 24424 9061
rect 25590 9052 25596 9104
rect 25648 9052 25654 9104
rect 25700 9064 26556 9092
rect 25700 9024 25728 9064
rect 23952 8996 25728 9024
rect 26053 9027 26111 9033
rect 23845 8987 23903 8993
rect 26053 8993 26065 9027
rect 26099 9024 26111 9027
rect 26418 9024 26424 9036
rect 26099 8996 26424 9024
rect 26099 8993 26111 8996
rect 26053 8987 26111 8993
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 19306 8928 21281 8956
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 22830 8916 22836 8968
rect 22888 8916 22894 8968
rect 21082 8888 21088 8900
rect 16500 8860 16896 8888
rect 16960 8860 21088 8888
rect 13648 8792 14136 8820
rect 14185 8823 14243 8829
rect 13541 8783 13599 8789
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 15010 8820 15016 8832
rect 14231 8792 15016 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 16500 8829 16528 8860
rect 16868 8832 16896 8860
rect 21082 8848 21088 8860
rect 21140 8848 21146 8900
rect 23109 8891 23167 8897
rect 23109 8857 23121 8891
rect 23155 8888 23167 8891
rect 23198 8888 23204 8900
rect 23155 8860 23204 8888
rect 23155 8857 23167 8860
rect 23109 8851 23167 8857
rect 23198 8848 23204 8860
rect 23256 8888 23262 8900
rect 23860 8888 23888 8987
rect 26418 8984 26424 8996
rect 26476 8984 26482 9036
rect 26528 9033 26556 9064
rect 26602 9052 26608 9104
rect 26660 9092 26666 9104
rect 26881 9095 26939 9101
rect 26881 9092 26893 9095
rect 26660 9064 26893 9092
rect 26660 9052 26666 9064
rect 26881 9061 26893 9064
rect 26927 9061 26939 9095
rect 26881 9055 26939 9061
rect 27062 9052 27068 9104
rect 27120 9092 27126 9104
rect 27249 9095 27307 9101
rect 27249 9092 27261 9095
rect 27120 9064 27261 9092
rect 27120 9052 27126 9064
rect 27249 9061 27261 9064
rect 27295 9061 27307 9095
rect 27249 9055 27307 9061
rect 27356 9064 27660 9092
rect 26513 9027 26571 9033
rect 26513 8993 26525 9027
rect 26559 8993 26571 9027
rect 26513 8987 26571 8993
rect 26694 8984 26700 9036
rect 26752 9024 26758 9036
rect 26789 9027 26847 9033
rect 26789 9024 26801 9027
rect 26752 8996 26801 9024
rect 26752 8984 26758 8996
rect 26789 8993 26801 8996
rect 26835 9024 26847 9027
rect 27157 9027 27215 9033
rect 27157 9024 27169 9027
rect 26835 8996 27169 9024
rect 26835 8993 26847 8996
rect 26789 8987 26847 8993
rect 27157 8993 27169 8996
rect 27203 9024 27215 9027
rect 27356 9024 27384 9064
rect 27632 9033 27660 9064
rect 28074 9052 28080 9104
rect 28132 9092 28138 9104
rect 28690 9095 28748 9101
rect 28690 9092 28702 9095
rect 28132 9064 28702 9092
rect 28132 9052 28138 9064
rect 28690 9061 28702 9064
rect 28736 9061 28748 9095
rect 28690 9055 28748 9061
rect 29362 9052 29368 9104
rect 29420 9092 29426 9104
rect 30006 9092 30012 9104
rect 29420 9064 30012 9092
rect 29420 9052 29426 9064
rect 30006 9052 30012 9064
rect 30064 9092 30070 9104
rect 30285 9095 30343 9101
rect 30285 9092 30297 9095
rect 30064 9064 30297 9092
rect 30064 9052 30070 9064
rect 30285 9061 30297 9064
rect 30331 9061 30343 9095
rect 30285 9055 30343 9061
rect 27525 9030 27583 9033
rect 27203 8996 27384 9024
rect 27448 9027 27583 9030
rect 27448 9002 27537 9027
rect 27203 8993 27215 8996
rect 27157 8987 27215 8993
rect 24118 8916 24124 8968
rect 24176 8916 24182 8968
rect 25222 8916 25228 8968
rect 25280 8956 25286 8968
rect 25685 8959 25743 8965
rect 25685 8956 25697 8959
rect 25280 8928 25697 8956
rect 25280 8916 25286 8928
rect 25685 8925 25697 8928
rect 25731 8925 25743 8959
rect 25685 8919 25743 8925
rect 25777 8959 25835 8965
rect 25777 8925 25789 8959
rect 25823 8956 25835 8959
rect 26326 8956 26332 8968
rect 25823 8928 26332 8956
rect 25823 8925 25835 8928
rect 25777 8919 25835 8925
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 27448 8956 27476 9002
rect 27525 8993 27537 9002
rect 27571 8993 27583 9027
rect 27525 8987 27583 8993
rect 27617 9027 27675 9033
rect 27617 8993 27629 9027
rect 27663 9024 27675 9027
rect 27982 9024 27988 9036
rect 27663 8996 27988 9024
rect 27663 8993 27675 8996
rect 27617 8987 27675 8993
rect 27982 8984 27988 8996
rect 28040 8984 28046 9036
rect 29178 8984 29184 9036
rect 29236 9024 29242 9036
rect 29730 9024 29736 9036
rect 29236 8996 29736 9024
rect 29236 8984 29242 8996
rect 29730 8984 29736 8996
rect 29788 9024 29794 9036
rect 30101 9027 30159 9033
rect 30101 9024 30113 9027
rect 29788 8996 30113 9024
rect 29788 8984 29794 8996
rect 30101 8993 30113 8996
rect 30147 8993 30159 9027
rect 30101 8987 30159 8993
rect 30190 8984 30196 9036
rect 30248 8984 30254 9036
rect 30469 9027 30527 9033
rect 30469 8993 30481 9027
rect 30515 8993 30527 9027
rect 30469 8987 30527 8993
rect 26620 8928 27476 8956
rect 23256 8860 23888 8888
rect 23256 8848 23262 8860
rect 16476 8823 16534 8829
rect 16476 8789 16488 8823
rect 16522 8789 16534 8823
rect 16476 8783 16534 8789
rect 16850 8780 16856 8832
rect 16908 8780 16914 8832
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 19116 8792 19533 8820
rect 19116 8780 19122 8792
rect 19521 8789 19533 8792
rect 19567 8789 19579 8823
rect 19521 8783 19579 8789
rect 19610 8780 19616 8832
rect 19668 8820 19674 8832
rect 22186 8820 22192 8832
rect 19668 8792 22192 8820
rect 19668 8780 19674 8792
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 23658 8780 23664 8832
rect 23716 8820 23722 8832
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 23716 8792 23765 8820
rect 23716 8780 23722 8792
rect 23753 8789 23765 8792
rect 23799 8789 23811 8823
rect 23860 8820 23888 8860
rect 26142 8848 26148 8900
rect 26200 8888 26206 8900
rect 26620 8888 26648 8928
rect 27798 8916 27804 8968
rect 27856 8956 27862 8968
rect 27893 8959 27951 8965
rect 27893 8956 27905 8959
rect 27856 8928 27905 8956
rect 27856 8916 27862 8928
rect 27893 8925 27905 8928
rect 27939 8925 27951 8959
rect 27893 8919 27951 8925
rect 28074 8916 28080 8968
rect 28132 8956 28138 8968
rect 28445 8959 28503 8965
rect 28445 8956 28457 8959
rect 28132 8928 28457 8956
rect 28132 8916 28138 8928
rect 28445 8925 28457 8928
rect 28491 8925 28503 8959
rect 28445 8919 28503 8925
rect 26200 8860 26648 8888
rect 26697 8891 26755 8897
rect 26200 8848 26206 8860
rect 26697 8857 26709 8891
rect 26743 8857 26755 8891
rect 26697 8851 26755 8857
rect 26789 8891 26847 8897
rect 26789 8857 26801 8891
rect 26835 8888 26847 8891
rect 27062 8888 27068 8900
rect 26835 8860 27068 8888
rect 26835 8857 26847 8860
rect 26789 8851 26847 8857
rect 24394 8820 24400 8832
rect 23860 8792 24400 8820
rect 23753 8783 23811 8789
rect 24394 8780 24400 8792
rect 24452 8780 24458 8832
rect 24486 8780 24492 8832
rect 24544 8820 24550 8832
rect 26602 8820 26608 8832
rect 24544 8792 26608 8820
rect 24544 8780 24550 8792
rect 26602 8780 26608 8792
rect 26660 8780 26666 8832
rect 26712 8820 26740 8851
rect 27062 8848 27068 8860
rect 27120 8848 27126 8900
rect 27157 8891 27215 8897
rect 27157 8857 27169 8891
rect 27203 8888 27215 8891
rect 27338 8888 27344 8900
rect 27203 8860 27344 8888
rect 27203 8857 27215 8860
rect 27157 8851 27215 8857
rect 27172 8820 27200 8851
rect 27338 8848 27344 8860
rect 27396 8848 27402 8900
rect 27430 8848 27436 8900
rect 27488 8848 27494 8900
rect 27522 8848 27528 8900
rect 27580 8888 27586 8900
rect 27709 8891 27767 8897
rect 27709 8888 27721 8891
rect 27580 8860 27721 8888
rect 27580 8848 27586 8860
rect 27709 8857 27721 8860
rect 27755 8857 27767 8891
rect 27709 8851 27767 8857
rect 29825 8891 29883 8897
rect 29825 8857 29837 8891
rect 29871 8888 29883 8891
rect 30484 8888 30512 8987
rect 29871 8860 30512 8888
rect 29871 8857 29883 8860
rect 29825 8851 29883 8857
rect 26712 8792 27200 8820
rect 27246 8780 27252 8832
rect 27304 8820 27310 8832
rect 27448 8820 27476 8848
rect 27617 8823 27675 8829
rect 27617 8820 27629 8823
rect 27304 8792 27629 8820
rect 27304 8780 27310 8792
rect 27617 8789 27629 8792
rect 27663 8789 27675 8823
rect 27617 8783 27675 8789
rect 27890 8780 27896 8832
rect 27948 8820 27954 8832
rect 27985 8823 28043 8829
rect 27985 8820 27997 8823
rect 27948 8792 27997 8820
rect 27948 8780 27954 8792
rect 27985 8789 27997 8792
rect 28031 8789 28043 8823
rect 27985 8783 28043 8789
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 4798 8616 4804 8628
rect 4663 8588 4804 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 4982 8576 4988 8628
rect 5040 8576 5046 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 7190 8576 7196 8628
rect 7248 8576 7254 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 11146 8616 11152 8628
rect 9088 8588 11152 8616
rect 9088 8576 9094 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11793 8619 11851 8625
rect 11793 8585 11805 8619
rect 11839 8616 11851 8619
rect 11839 8588 12112 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 7006 8548 7012 8560
rect 6196 8520 7012 8548
rect 6196 8480 6224 8520
rect 7006 8508 7012 8520
rect 7064 8508 7070 8560
rect 5552 8452 6224 8480
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 4062 8412 4068 8424
rect 3283 8384 4068 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 5552 8421 5580 8452
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 3482 8347 3540 8353
rect 3482 8344 3494 8347
rect 3252 8316 3494 8344
rect 3252 8288 3280 8316
rect 3482 8313 3494 8316
rect 3528 8313 3540 8347
rect 5184 8344 5212 8375
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6196 8421 6224 8452
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 6457 8483 6515 8489
rect 6457 8449 6469 8483
rect 6503 8480 6515 8483
rect 7098 8480 7104 8492
rect 6503 8452 7104 8480
rect 6503 8449 6515 8452
rect 6457 8443 6515 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7208 8480 7236 8576
rect 12084 8560 12112 8588
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13780 8588 13829 8616
rect 13780 8576 13786 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 19702 8616 19708 8628
rect 13817 8579 13875 8585
rect 14476 8588 19708 8616
rect 10873 8551 10931 8557
rect 10873 8517 10885 8551
rect 10919 8548 10931 8551
rect 10919 8520 11928 8548
rect 10919 8517 10931 8520
rect 10873 8511 10931 8517
rect 7208 8452 7512 8480
rect 6181 8415 6239 8421
rect 5960 8384 6132 8412
rect 5960 8372 5966 8384
rect 6104 8344 6132 8384
rect 6181 8381 6193 8415
rect 6227 8381 6239 8415
rect 6181 8375 6239 8381
rect 6273 8415 6331 8421
rect 6273 8381 6285 8415
rect 6319 8412 6331 8415
rect 6380 8412 6408 8440
rect 6319 8384 6408 8412
rect 6549 8415 6607 8421
rect 6319 8381 6331 8384
rect 6273 8375 6331 8381
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6564 8344 6592 8375
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6696 8384 6837 8412
rect 6696 8372 6702 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8381 7067 8415
rect 7116 8412 7144 8440
rect 7484 8421 7512 8452
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8846 8480 8852 8492
rect 8536 8452 8852 8480
rect 8536 8440 8542 8452
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 10410 8480 10416 8492
rect 10284 8452 10416 8480
rect 10284 8440 10290 8452
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 11900 8489 11928 8520
rect 12066 8508 12072 8560
rect 12124 8508 12130 8560
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 14476 8557 14504 8588
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 19981 8619 20039 8625
rect 19981 8585 19993 8619
rect 20027 8616 20039 8619
rect 20070 8616 20076 8628
rect 20027 8588 20076 8616
rect 20027 8585 20039 8588
rect 19981 8579 20039 8585
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 21174 8576 21180 8628
rect 21232 8576 21238 8628
rect 23014 8576 23020 8628
rect 23072 8616 23078 8628
rect 23109 8619 23167 8625
rect 23109 8616 23121 8619
rect 23072 8588 23121 8616
rect 23072 8576 23078 8588
rect 23109 8585 23121 8588
rect 23155 8585 23167 8619
rect 24486 8616 24492 8628
rect 23109 8579 23167 8585
rect 23308 8588 24492 8616
rect 14461 8551 14519 8557
rect 12216 8520 12480 8548
rect 12216 8508 12222 8520
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 10888 8452 11253 8480
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 7116 8384 7205 8412
rect 7009 8375 7067 8381
rect 7193 8381 7205 8384
rect 7239 8412 7251 8415
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 7239 8384 7297 8412
rect 7239 8381 7251 8384
rect 7193 8375 7251 8381
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 9116 8415 9174 8421
rect 9116 8381 9128 8415
rect 9162 8412 9174 8415
rect 9398 8412 9404 8424
rect 9162 8384 9404 8412
rect 9162 8381 9174 8384
rect 9116 8375 9174 8381
rect 6730 8344 6736 8356
rect 5184 8316 5856 8344
rect 6104 8316 6736 8344
rect 3482 8307 3540 8313
rect 3234 8236 3240 8288
rect 3292 8236 3298 8288
rect 5828 8276 5856 8316
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7024 8344 7052 8375
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 10686 8412 10692 8424
rect 10008 8384 10692 8412
rect 10008 8372 10014 8384
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 10888 8421 10916 8452
rect 11241 8449 11253 8452
rect 11287 8449 11299 8483
rect 11885 8483 11943 8489
rect 11241 8443 11299 8449
rect 11348 8452 11836 8480
rect 11348 8424 11376 8452
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8381 11023 8415
rect 10965 8375 11023 8381
rect 6972 8316 7052 8344
rect 6972 8304 6978 8316
rect 7374 8304 7380 8356
rect 7432 8304 7438 8356
rect 10980 8344 11008 8375
rect 11146 8372 11152 8424
rect 11204 8372 11210 8424
rect 11330 8372 11336 8424
rect 11388 8372 11394 8424
rect 11808 8421 11836 8452
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 12342 8440 12348 8492
rect 12400 8440 12406 8492
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11839 8410 11931 8412
rect 11992 8410 12173 8412
rect 11839 8384 12173 8410
rect 11839 8381 11851 8384
rect 11903 8382 12020 8384
rect 11793 8375 11851 8381
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12360 8412 12388 8440
rect 12452 8421 12480 8520
rect 14461 8517 14473 8551
rect 14507 8517 14519 8551
rect 14461 8511 14519 8517
rect 15470 8508 15476 8560
rect 15528 8548 15534 8560
rect 16761 8551 16819 8557
rect 16761 8548 16773 8551
rect 15528 8520 16773 8548
rect 15528 8508 15534 8520
rect 12728 8452 14320 8480
rect 12299 8384 12388 8412
rect 12437 8415 12495 8421
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12526 8412 12532 8424
rect 12483 8384 12532 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 7484 8316 11008 8344
rect 7484 8276 7512 8316
rect 5828 8248 7512 8276
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10229 8279 10287 8285
rect 10229 8276 10241 8279
rect 10100 8248 10241 8276
rect 10100 8236 10106 8248
rect 10229 8245 10241 8248
rect 10275 8245 10287 8279
rect 10980 8276 11008 8316
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8344 11115 8347
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11103 8316 11529 8344
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 11146 8276 11152 8288
rect 10980 8248 11152 8276
rect 10229 8239 10287 8245
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 11716 8276 11744 8375
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 12728 8421 12756 8452
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 12728 8344 12756 8375
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 14292 8421 14320 8452
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13964 8384 14013 8412
rect 13964 8372 13970 8384
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 12124 8316 12756 8344
rect 12124 8304 12130 8316
rect 12802 8304 12808 8356
rect 12860 8344 12866 8356
rect 14108 8344 14136 8375
rect 14366 8372 14372 8424
rect 14424 8412 14430 8424
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 14424 8384 14473 8412
rect 14424 8372 14430 8384
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 15838 8372 15844 8424
rect 15896 8372 15902 8424
rect 16316 8421 16344 8520
rect 16761 8517 16773 8520
rect 16807 8548 16819 8551
rect 17034 8548 17040 8560
rect 16807 8520 17040 8548
rect 16807 8517 16819 8520
rect 16761 8511 16819 8517
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 19334 8548 19340 8560
rect 19306 8508 19340 8548
rect 19392 8548 19398 8560
rect 19392 8520 20116 8548
rect 19392 8508 19398 8520
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 19306 8480 19334 8508
rect 18800 8452 19334 8480
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 16482 8372 16488 8424
rect 16540 8372 16546 8424
rect 16577 8415 16635 8421
rect 16577 8381 16589 8415
rect 16623 8412 16635 8415
rect 16850 8412 16856 8424
rect 16623 8384 16856 8412
rect 16623 8381 16635 8384
rect 16577 8375 16635 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 18800 8406 18828 8452
rect 19518 8440 19524 8492
rect 19576 8440 19582 8492
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 19978 8480 19984 8492
rect 19659 8452 19984 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 18878 8409 18936 8415
rect 18878 8406 18890 8409
rect 18800 8378 18890 8406
rect 18878 8375 18890 8378
rect 18924 8375 18936 8409
rect 18878 8369 18936 8375
rect 19058 8372 19064 8424
rect 19116 8372 19122 8424
rect 19242 8372 19248 8424
rect 19300 8372 19306 8424
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 19536 8412 19564 8440
rect 19392 8384 19564 8412
rect 19392 8372 19398 8384
rect 12860 8316 14136 8344
rect 17396 8347 17454 8353
rect 12860 8304 12866 8316
rect 17396 8313 17408 8347
rect 17442 8344 17454 8347
rect 17678 8344 17684 8356
rect 17442 8316 17684 8344
rect 17442 8313 17454 8316
rect 17396 8307 17454 8313
rect 17678 8304 17684 8316
rect 17736 8304 17742 8356
rect 17788 8316 18828 8344
rect 12158 8276 12164 8288
rect 11716 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 12345 8279 12403 8285
rect 12345 8245 12357 8279
rect 12391 8276 12403 8279
rect 12434 8276 12440 8288
rect 12391 8248 12440 8276
rect 12391 8245 12403 8248
rect 12345 8239 12403 8245
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 12526 8236 12532 8288
rect 12584 8236 12590 8288
rect 16301 8279 16359 8285
rect 16301 8245 16313 8279
rect 16347 8276 16359 8279
rect 16390 8276 16396 8288
rect 16347 8248 16396 8276
rect 16347 8245 16359 8248
rect 16301 8239 16359 8245
rect 16390 8236 16396 8248
rect 16448 8276 16454 8288
rect 16574 8276 16580 8288
rect 16448 8248 16580 8276
rect 16448 8236 16454 8248
rect 16574 8236 16580 8248
rect 16632 8276 16638 8288
rect 17788 8276 17816 8316
rect 16632 8248 17816 8276
rect 16632 8236 16638 8248
rect 18506 8236 18512 8288
rect 18564 8236 18570 8288
rect 18690 8236 18696 8288
rect 18748 8236 18754 8288
rect 18800 8276 18828 8316
rect 18966 8304 18972 8356
rect 19024 8304 19030 8356
rect 19150 8304 19156 8356
rect 19208 8344 19214 8356
rect 19628 8344 19656 8443
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 19702 8372 19708 8424
rect 19760 8372 19766 8424
rect 19797 8415 19855 8421
rect 19797 8381 19809 8415
rect 19843 8412 19855 8415
rect 20088 8412 20116 8520
rect 22462 8508 22468 8560
rect 22520 8548 22526 8560
rect 23308 8548 23336 8588
rect 24486 8576 24492 8588
rect 24544 8576 24550 8628
rect 25314 8576 25320 8628
rect 25372 8616 25378 8628
rect 25409 8619 25467 8625
rect 25409 8616 25421 8619
rect 25372 8588 25421 8616
rect 25372 8576 25378 8588
rect 25409 8585 25421 8588
rect 25455 8585 25467 8619
rect 25409 8579 25467 8585
rect 25774 8576 25780 8628
rect 25832 8576 25838 8628
rect 27246 8616 27252 8628
rect 26436 8588 27252 8616
rect 22520 8520 23336 8548
rect 22520 8508 22526 8520
rect 23658 8508 23664 8560
rect 23716 8508 23722 8560
rect 23842 8508 23848 8560
rect 23900 8548 23906 8560
rect 23937 8551 23995 8557
rect 23937 8548 23949 8551
rect 23900 8520 23949 8548
rect 23900 8508 23906 8520
rect 23937 8517 23949 8520
rect 23983 8517 23995 8551
rect 23937 8511 23995 8517
rect 23017 8483 23075 8489
rect 21008 8452 22968 8480
rect 21008 8421 21036 8452
rect 19843 8384 20116 8412
rect 20993 8415 21051 8421
rect 19843 8381 19855 8384
rect 19797 8375 19855 8381
rect 20993 8381 21005 8415
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 21082 8372 21088 8424
rect 21140 8412 21146 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 21140 8384 22569 8412
rect 21140 8372 21146 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 22738 8372 22744 8424
rect 22796 8372 22802 8424
rect 19208 8316 19656 8344
rect 19720 8344 19748 8372
rect 22462 8344 22468 8356
rect 19720 8316 22468 8344
rect 19208 8304 19214 8316
rect 22462 8304 22468 8316
rect 22520 8304 22526 8356
rect 22649 8347 22707 8353
rect 22649 8313 22661 8347
rect 22695 8344 22707 8347
rect 22833 8347 22891 8353
rect 22833 8344 22845 8347
rect 22695 8316 22845 8344
rect 22695 8313 22707 8316
rect 22649 8307 22707 8313
rect 22833 8313 22845 8316
rect 22879 8313 22891 8347
rect 22940 8344 22968 8452
rect 23017 8449 23029 8483
rect 23063 8480 23075 8483
rect 23198 8480 23204 8492
rect 23063 8452 23204 8480
rect 23063 8449 23075 8452
rect 23017 8443 23075 8449
rect 23198 8440 23204 8452
rect 23256 8440 23262 8492
rect 23676 8480 23704 8508
rect 25792 8480 25820 8576
rect 23308 8452 23520 8480
rect 23676 8452 24256 8480
rect 23106 8372 23112 8424
rect 23164 8412 23170 8424
rect 23308 8412 23336 8452
rect 23492 8421 23520 8452
rect 24228 8421 24256 8452
rect 25608 8452 25820 8480
rect 23164 8384 23336 8412
rect 23385 8415 23443 8421
rect 23164 8372 23170 8384
rect 23385 8381 23397 8415
rect 23431 8381 23443 8415
rect 23385 8375 23443 8381
rect 23477 8415 23535 8421
rect 23477 8381 23489 8415
rect 23523 8412 23535 8415
rect 23845 8415 23903 8421
rect 23845 8412 23857 8415
rect 23523 8384 23857 8412
rect 23523 8381 23535 8384
rect 23477 8375 23535 8381
rect 23845 8381 23857 8384
rect 23891 8412 23903 8415
rect 24213 8415 24271 8421
rect 23891 8384 24072 8412
rect 23891 8381 23903 8384
rect 23845 8375 23903 8381
rect 22940 8316 23152 8344
rect 22833 8307 22891 8313
rect 21726 8276 21732 8288
rect 18800 8248 21732 8276
rect 21726 8236 21732 8248
rect 21784 8236 21790 8288
rect 23124 8276 23152 8316
rect 23198 8304 23204 8356
rect 23256 8304 23262 8356
rect 23400 8344 23428 8375
rect 23400 8316 23888 8344
rect 23477 8279 23535 8285
rect 23477 8276 23489 8279
rect 23124 8248 23489 8276
rect 23477 8245 23489 8248
rect 23523 8276 23535 8279
rect 23750 8276 23756 8288
rect 23523 8248 23756 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23750 8236 23756 8248
rect 23808 8236 23814 8288
rect 23860 8285 23888 8316
rect 23845 8279 23903 8285
rect 23845 8245 23857 8279
rect 23891 8276 23903 8279
rect 23934 8276 23940 8288
rect 23891 8248 23940 8276
rect 23891 8245 23903 8248
rect 23845 8239 23903 8245
rect 23934 8236 23940 8248
rect 23992 8236 23998 8288
rect 24044 8276 24072 8384
rect 24213 8381 24225 8415
rect 24259 8381 24271 8415
rect 24213 8375 24271 8381
rect 24394 8372 24400 8424
rect 24452 8372 24458 8424
rect 25608 8421 25636 8452
rect 25593 8415 25651 8421
rect 25593 8381 25605 8415
rect 25639 8381 25651 8415
rect 25593 8375 25651 8381
rect 25682 8372 25688 8424
rect 25740 8372 25746 8424
rect 25866 8372 25872 8424
rect 25924 8372 25930 8424
rect 25958 8372 25964 8424
rect 26016 8372 26022 8424
rect 26436 8421 26464 8588
rect 27246 8576 27252 8588
rect 27304 8576 27310 8628
rect 27798 8576 27804 8628
rect 27856 8616 27862 8628
rect 27893 8619 27951 8625
rect 27893 8616 27905 8619
rect 27856 8588 27905 8616
rect 27856 8576 27862 8588
rect 27893 8585 27905 8588
rect 27939 8585 27951 8619
rect 27893 8579 27951 8585
rect 30190 8576 30196 8628
rect 30248 8616 30254 8628
rect 30377 8619 30435 8625
rect 30377 8616 30389 8619
rect 30248 8588 30389 8616
rect 30248 8576 30254 8588
rect 30377 8585 30389 8588
rect 30423 8585 30435 8619
rect 30377 8579 30435 8585
rect 26605 8551 26663 8557
rect 26605 8517 26617 8551
rect 26651 8548 26663 8551
rect 27614 8548 27620 8560
rect 26651 8520 27620 8548
rect 26651 8517 26663 8520
rect 26605 8511 26663 8517
rect 27614 8508 27620 8520
rect 27672 8508 27678 8560
rect 27985 8483 28043 8489
rect 27985 8480 27997 8483
rect 26620 8452 27997 8480
rect 26620 8421 26648 8452
rect 27985 8449 27997 8452
rect 28031 8449 28043 8483
rect 27985 8443 28043 8449
rect 26421 8415 26479 8421
rect 26421 8381 26433 8415
rect 26467 8381 26479 8415
rect 26421 8375 26479 8381
rect 26605 8415 26663 8421
rect 26605 8381 26617 8415
rect 26651 8381 26663 8415
rect 26605 8375 26663 8381
rect 26697 8415 26755 8421
rect 26697 8381 26709 8415
rect 26743 8381 26755 8415
rect 26697 8375 26755 8381
rect 24121 8347 24179 8353
rect 24121 8313 24133 8347
rect 24167 8344 24179 8347
rect 24305 8347 24363 8353
rect 24305 8344 24317 8347
rect 24167 8316 24317 8344
rect 24167 8313 24179 8316
rect 24121 8307 24179 8313
rect 24305 8313 24317 8316
rect 24351 8313 24363 8347
rect 26712 8344 26740 8375
rect 26878 8372 26884 8424
rect 26936 8372 26942 8424
rect 26973 8415 27031 8421
rect 26973 8381 26985 8415
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 26712 8316 26924 8344
rect 24305 8307 24363 8313
rect 26896 8288 26924 8316
rect 26142 8276 26148 8288
rect 24044 8248 26148 8276
rect 26142 8236 26148 8248
rect 26200 8236 26206 8288
rect 26786 8236 26792 8288
rect 26844 8236 26850 8288
rect 26878 8236 26884 8288
rect 26936 8236 26942 8288
rect 26988 8276 27016 8375
rect 27062 8372 27068 8424
rect 27120 8372 27126 8424
rect 27154 8372 27160 8424
rect 27212 8412 27218 8424
rect 27341 8415 27399 8421
rect 27341 8412 27353 8415
rect 27212 8384 27353 8412
rect 27212 8372 27218 8384
rect 27341 8381 27353 8384
rect 27387 8381 27399 8415
rect 27341 8375 27399 8381
rect 27709 8415 27767 8421
rect 27709 8381 27721 8415
rect 27755 8381 27767 8415
rect 27709 8375 27767 8381
rect 27080 8344 27108 8372
rect 27724 8344 27752 8375
rect 27890 8372 27896 8424
rect 27948 8372 27954 8424
rect 28261 8415 28319 8421
rect 28261 8381 28273 8415
rect 28307 8381 28319 8415
rect 28261 8375 28319 8381
rect 28276 8344 28304 8375
rect 28994 8372 29000 8424
rect 29052 8372 29058 8424
rect 29242 8347 29300 8353
rect 29242 8344 29254 8347
rect 27080 8316 28304 8344
rect 28460 8316 29254 8344
rect 27062 8276 27068 8288
rect 26988 8248 27068 8276
rect 27062 8236 27068 8248
rect 27120 8236 27126 8288
rect 27154 8236 27160 8288
rect 27212 8236 27218 8288
rect 27246 8236 27252 8288
rect 27304 8276 27310 8288
rect 27525 8279 27583 8285
rect 27525 8276 27537 8279
rect 27304 8248 27537 8276
rect 27304 8236 27310 8248
rect 27525 8245 27537 8248
rect 27571 8245 27583 8279
rect 27525 8239 27583 8245
rect 27614 8236 27620 8288
rect 27672 8276 27678 8288
rect 27798 8276 27804 8288
rect 27672 8248 27804 8276
rect 27672 8236 27678 8248
rect 27798 8236 27804 8248
rect 27856 8236 27862 8288
rect 28460 8285 28488 8316
rect 29242 8313 29254 8316
rect 29288 8313 29300 8347
rect 29242 8307 29300 8313
rect 28445 8279 28503 8285
rect 28445 8245 28457 8279
rect 28491 8245 28503 8279
rect 28445 8239 28503 8245
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 5902 8072 5908 8084
rect 5307 8044 5908 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7064 8044 7297 8072
rect 7064 8032 7070 8044
rect 7285 8041 7297 8044
rect 7331 8072 7343 8075
rect 7926 8072 7932 8084
rect 7331 8044 7932 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 9033 8075 9091 8081
rect 9033 8041 9045 8075
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 7208 7976 8984 8004
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5997 7939 6055 7945
rect 5997 7936 6009 7939
rect 5399 7908 6009 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5997 7905 6009 7908
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 6638 7936 6644 7948
rect 6503 7908 6644 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 4816 7800 4844 7899
rect 5184 7868 5212 7899
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 6730 7896 6736 7948
rect 6788 7896 6794 7948
rect 7098 7896 7104 7948
rect 7156 7896 7162 7948
rect 7208 7945 7236 7976
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 7742 7896 7748 7948
rect 7800 7936 7806 7948
rect 7909 7939 7967 7945
rect 7909 7936 7921 7939
rect 7800 7908 7921 7936
rect 7800 7896 7806 7908
rect 7909 7905 7921 7908
rect 7955 7905 7967 7939
rect 7909 7899 7967 7905
rect 7006 7868 7012 7880
rect 5184 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7837 7711 7871
rect 8956 7868 8984 7976
rect 9048 7936 9076 8035
rect 9674 8032 9680 8084
rect 9732 8032 9738 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 11054 8072 11060 8084
rect 10643 8044 11060 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 9692 8004 9720 8032
rect 9769 8007 9827 8013
rect 9769 8004 9781 8007
rect 9692 7976 9781 8004
rect 9769 7973 9781 7976
rect 9815 7973 9827 8007
rect 9769 7967 9827 7973
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 10042 8004 10048 8016
rect 9907 7976 10048 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9048 7908 9597 7936
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 9950 7896 9956 7948
rect 10008 7896 10014 7948
rect 10152 7942 10180 8035
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8041 11207 8075
rect 11149 8035 11207 8041
rect 10686 7964 10692 8016
rect 10744 8004 10750 8016
rect 11164 8004 11192 8035
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 13357 8075 13415 8081
rect 11572 8044 11744 8072
rect 11572 8032 11578 8044
rect 10744 7976 11652 8004
rect 10744 7964 10750 7976
rect 10217 7945 10275 7951
rect 10217 7942 10229 7945
rect 10152 7914 10229 7942
rect 10217 7911 10229 7914
rect 10263 7911 10275 7945
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10217 7905 10275 7911
rect 11072 7908 11161 7936
rect 9674 7868 9680 7880
rect 8956 7840 9680 7868
rect 7653 7831 7711 7837
rect 4816 7772 5488 7800
rect 5460 7744 5488 7772
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 7668 7800 7696 7831
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10502 7868 10508 7880
rect 10367 7840 10508 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 6604 7772 7696 7800
rect 9692 7800 9720 7828
rect 11072 7800 11100 7908
rect 11149 7905 11161 7908
rect 11195 7936 11207 7939
rect 11330 7936 11336 7948
rect 11195 7908 11336 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 11330 7896 11336 7908
rect 11388 7936 11394 7948
rect 11624 7945 11652 7976
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 11388 7908 11529 7936
rect 11388 7896 11394 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11422 7828 11428 7880
rect 11480 7828 11486 7880
rect 11716 7868 11744 8044
rect 13357 8041 13369 8075
rect 13403 8041 13415 8075
rect 13357 8035 13415 8041
rect 13449 8075 13507 8081
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 13538 8072 13544 8084
rect 13495 8044 13544 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 12244 8007 12302 8013
rect 12244 7973 12256 8007
rect 12290 8004 12302 8007
rect 12526 8004 12532 8016
rect 12290 7976 12532 8004
rect 12290 7973 12302 7976
rect 12244 7967 12302 7973
rect 12526 7964 12532 7976
rect 12584 7964 12590 8016
rect 13372 8004 13400 8035
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 14274 8072 14280 8084
rect 13688 8044 14280 8072
rect 13688 8032 13694 8044
rect 14274 8032 14280 8044
rect 14332 8072 14338 8084
rect 14332 8044 15148 8072
rect 14332 8032 14338 8044
rect 15120 8016 15148 8044
rect 15378 8032 15384 8084
rect 15436 8032 15442 8084
rect 16482 8032 16488 8084
rect 16540 8032 16546 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16816 8044 16957 8072
rect 16816 8032 16822 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 16945 8035 17003 8041
rect 13725 8007 13783 8013
rect 13725 8004 13737 8007
rect 13372 7976 13737 8004
rect 13725 7973 13737 7976
rect 13771 7973 13783 8007
rect 13725 7967 13783 7973
rect 13814 7964 13820 8016
rect 13872 7964 13878 8016
rect 15102 7964 15108 8016
rect 15160 8004 15166 8016
rect 16500 8004 16528 8032
rect 16853 8007 16911 8013
rect 16853 8004 16865 8007
rect 15160 7976 15700 8004
rect 16500 7976 16865 8004
rect 15160 7964 15166 7976
rect 11790 7896 11796 7948
rect 11848 7896 11854 7948
rect 13630 7945 13636 7948
rect 13628 7936 13636 7945
rect 13591 7908 13636 7936
rect 13628 7899 13636 7908
rect 13630 7896 13636 7899
rect 13688 7896 13694 7948
rect 13945 7939 14003 7945
rect 13945 7936 13957 7939
rect 13740 7908 13957 7936
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11716 7840 11989 7868
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 13740 7868 13768 7908
rect 13945 7905 13957 7908
rect 13991 7905 14003 7939
rect 13945 7899 14003 7905
rect 14093 7939 14151 7945
rect 14093 7905 14105 7939
rect 14139 7905 14151 7939
rect 14093 7899 14151 7905
rect 14108 7868 14136 7899
rect 15010 7896 15016 7948
rect 15068 7896 15074 7948
rect 15672 7945 15700 7976
rect 16853 7973 16865 7976
rect 16899 7973 16911 8007
rect 16853 7967 16911 7973
rect 15197 7939 15255 7945
rect 15197 7905 15209 7939
rect 15243 7936 15255 7939
rect 15473 7939 15531 7945
rect 15473 7936 15485 7939
rect 15243 7908 15485 7936
rect 15243 7905 15255 7908
rect 15197 7899 15255 7905
rect 15473 7905 15485 7908
rect 15519 7905 15531 7939
rect 15473 7899 15531 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16298 7896 16304 7948
rect 16356 7896 16362 7948
rect 16390 7896 16396 7948
rect 16448 7896 16454 7948
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 16574 7936 16580 7948
rect 16531 7908 16580 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 16669 7899 16727 7905
rect 13228 7840 13768 7868
rect 13924 7840 14136 7868
rect 13228 7828 13234 7840
rect 9692 7772 11100 7800
rect 6604 7760 6610 7772
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 11241 7803 11299 7809
rect 11241 7800 11253 7803
rect 11204 7772 11253 7800
rect 11204 7760 11210 7772
rect 11241 7769 11253 7772
rect 11287 7800 11299 7803
rect 11517 7803 11575 7809
rect 11517 7800 11529 7803
rect 11287 7772 11529 7800
rect 11287 7769 11299 7772
rect 11241 7763 11299 7769
rect 11517 7769 11529 7772
rect 11563 7769 11575 7803
rect 11517 7763 11575 7769
rect 5442 7692 5448 7744
rect 5500 7692 5506 7744
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 6178 7732 6184 7744
rect 5675 7704 6184 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 13924 7732 13952 7840
rect 14108 7800 14136 7840
rect 15286 7828 15292 7880
rect 15344 7868 15350 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15344 7840 15853 7868
rect 15344 7828 15350 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16684 7868 16712 7899
rect 16172 7840 16712 7868
rect 16960 7868 16988 8035
rect 17678 8032 17684 8084
rect 17736 8032 17742 8084
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 18472 8044 18705 8072
rect 18472 8032 18478 8044
rect 18693 8041 18705 8044
rect 18739 8041 18751 8075
rect 18693 8035 18751 8041
rect 19061 8075 19119 8081
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19242 8072 19248 8084
rect 19107 8044 19248 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 19426 8072 19432 8084
rect 19352 8044 19432 8072
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 19352 8013 19380 8044
rect 19426 8032 19432 8044
rect 19484 8072 19490 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 19484 8044 20269 8072
rect 19484 8032 19490 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 20257 8035 20315 8041
rect 22738 8032 22744 8084
rect 22796 8032 22802 8084
rect 23017 8075 23075 8081
rect 23017 8041 23029 8075
rect 23063 8072 23075 8075
rect 23198 8072 23204 8084
rect 23063 8044 23204 8072
rect 23063 8041 23075 8044
rect 23017 8035 23075 8041
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 25682 8032 25688 8084
rect 25740 8032 25746 8084
rect 25958 8032 25964 8084
rect 26016 8072 26022 8084
rect 29549 8075 29607 8081
rect 29549 8072 29561 8075
rect 26016 8044 29561 8072
rect 26016 8032 26022 8044
rect 29549 8041 29561 8044
rect 29595 8041 29607 8075
rect 29549 8035 29607 8041
rect 18601 8007 18659 8013
rect 18601 8004 18613 8007
rect 17092 7976 18613 8004
rect 17092 7964 17098 7976
rect 18601 7973 18613 7976
rect 18647 8004 18659 8007
rect 19337 8007 19395 8013
rect 19337 8004 19349 8007
rect 18647 7976 19349 8004
rect 18647 7973 18659 7976
rect 18601 7967 18659 7973
rect 19337 7973 19349 7976
rect 19383 7973 19395 8007
rect 19337 7967 19395 7973
rect 19797 8007 19855 8013
rect 19797 7973 19809 8007
rect 19843 8004 19855 8007
rect 20349 8007 20407 8013
rect 20349 8004 20361 8007
rect 19843 7976 20361 8004
rect 19843 7973 19855 7976
rect 19797 7967 19855 7973
rect 20349 7973 20361 7976
rect 20395 7973 20407 8007
rect 22756 8004 22784 8032
rect 22756 7976 23152 8004
rect 20349 7967 20407 7973
rect 17126 7896 17132 7948
rect 17184 7936 17190 7948
rect 17497 7939 17555 7945
rect 17497 7936 17509 7939
rect 17184 7908 17509 7936
rect 17184 7896 17190 7908
rect 17497 7905 17509 7908
rect 17543 7936 17555 7939
rect 17678 7936 17684 7948
rect 17543 7908 17684 7936
rect 17543 7905 17555 7908
rect 17497 7899 17555 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17862 7896 17868 7948
rect 17920 7896 17926 7948
rect 18230 7896 18236 7948
rect 18288 7936 18294 7948
rect 18810 7939 18868 7945
rect 18810 7936 18822 7939
rect 18288 7908 18822 7936
rect 18288 7896 18294 7908
rect 18810 7905 18822 7908
rect 18856 7905 18868 7939
rect 18810 7899 18868 7905
rect 19245 7939 19303 7945
rect 19245 7905 19257 7939
rect 19291 7936 19303 7939
rect 19518 7936 19524 7948
rect 19291 7908 19524 7936
rect 19291 7905 19303 7908
rect 19245 7899 19303 7905
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 18322 7868 18328 7880
rect 16960 7840 18328 7868
rect 16172 7828 16178 7840
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 18414 7828 18420 7880
rect 18472 7868 18478 7880
rect 19812 7868 19840 7967
rect 20070 7896 20076 7948
rect 20128 7936 20134 7948
rect 20466 7939 20524 7945
rect 20466 7936 20478 7939
rect 20128 7908 20478 7936
rect 20128 7896 20134 7908
rect 20466 7905 20478 7908
rect 20512 7905 20524 7939
rect 20466 7899 20524 7905
rect 22393 7939 22451 7945
rect 22393 7905 22405 7939
rect 22439 7936 22451 7939
rect 22925 7939 22983 7945
rect 22439 7908 22876 7936
rect 22439 7905 22451 7908
rect 22393 7899 22451 7905
rect 18472 7840 19840 7868
rect 19981 7871 20039 7877
rect 18472 7828 18478 7840
rect 19981 7837 19993 7871
rect 20027 7837 20039 7871
rect 19981 7831 20039 7837
rect 18340 7800 18368 7828
rect 19797 7803 19855 7809
rect 19797 7800 19809 7803
rect 14108 7772 17540 7800
rect 18340 7772 19809 7800
rect 13596 7704 13952 7732
rect 15197 7735 15255 7741
rect 13596 7692 13602 7704
rect 15197 7701 15209 7735
rect 15243 7732 15255 7735
rect 16117 7735 16175 7741
rect 16117 7732 16129 7735
rect 15243 7704 16129 7732
rect 15243 7701 15255 7704
rect 15197 7695 15255 7701
rect 16117 7701 16129 7704
rect 16163 7701 16175 7735
rect 16117 7695 16175 7701
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 17405 7735 17463 7741
rect 17405 7732 17417 7735
rect 16264 7704 17417 7732
rect 16264 7692 16270 7704
rect 17405 7701 17417 7704
rect 17451 7701 17463 7735
rect 17512 7732 17540 7772
rect 19797 7769 19809 7772
rect 19843 7800 19855 7803
rect 19996 7800 20024 7831
rect 22646 7828 22652 7880
rect 22704 7828 22710 7880
rect 22848 7868 22876 7908
rect 22925 7905 22937 7939
rect 22971 7936 22983 7939
rect 23014 7936 23020 7948
rect 22971 7908 23020 7936
rect 22971 7905 22983 7908
rect 22925 7899 22983 7905
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 23124 7945 23152 7976
rect 23400 7976 24072 8004
rect 23400 7945 23428 7976
rect 24044 7948 24072 7976
rect 24136 7976 24348 8004
rect 24136 7948 24164 7976
rect 23109 7939 23167 7945
rect 23109 7905 23121 7939
rect 23155 7936 23167 7939
rect 23385 7939 23443 7945
rect 23155 7908 23336 7936
rect 23155 7905 23167 7908
rect 23109 7899 23167 7905
rect 23308 7880 23336 7908
rect 23385 7905 23397 7939
rect 23431 7905 23443 7939
rect 23753 7939 23811 7945
rect 23753 7936 23765 7939
rect 23385 7899 23443 7905
rect 23584 7908 23765 7936
rect 22848 7840 23244 7868
rect 23216 7809 23244 7840
rect 23290 7828 23296 7880
rect 23348 7868 23354 7880
rect 23584 7868 23612 7908
rect 23753 7905 23765 7908
rect 23799 7905 23811 7939
rect 23753 7899 23811 7905
rect 23842 7896 23848 7948
rect 23900 7936 23906 7948
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 23900 7908 23949 7936
rect 23900 7896 23906 7908
rect 23937 7905 23949 7908
rect 23983 7905 23995 7939
rect 23937 7899 23995 7905
rect 24026 7896 24032 7948
rect 24084 7896 24090 7948
rect 24118 7896 24124 7948
rect 24176 7896 24182 7948
rect 24320 7945 24348 7976
rect 26786 7964 26792 8016
rect 26844 8004 26850 8016
rect 27341 8007 27399 8013
rect 27341 8004 27353 8007
rect 26844 7976 27353 8004
rect 26844 7964 26850 7976
rect 27341 7973 27353 7976
rect 27387 7973 27399 8007
rect 27798 8004 27804 8016
rect 27341 7967 27399 7973
rect 27724 7976 27804 8004
rect 24213 7939 24271 7945
rect 24213 7905 24225 7939
rect 24259 7905 24271 7939
rect 24213 7899 24271 7905
rect 24305 7939 24363 7945
rect 24305 7905 24317 7939
rect 24351 7905 24363 7939
rect 24305 7899 24363 7905
rect 23348 7840 23612 7868
rect 23661 7871 23719 7877
rect 23348 7828 23354 7840
rect 23661 7837 23673 7871
rect 23707 7868 23719 7871
rect 24228 7868 24256 7899
rect 24394 7896 24400 7948
rect 24452 7936 24458 7948
rect 24561 7939 24619 7945
rect 24561 7936 24573 7939
rect 24452 7908 24573 7936
rect 24452 7896 24458 7908
rect 24561 7905 24573 7908
rect 24607 7905 24619 7939
rect 24561 7899 24619 7905
rect 26878 7896 26884 7948
rect 26936 7936 26942 7948
rect 27154 7936 27160 7948
rect 26936 7908 27160 7936
rect 26936 7896 26942 7908
rect 27154 7896 27160 7908
rect 27212 7896 27218 7948
rect 27246 7896 27252 7948
rect 27304 7896 27310 7948
rect 27448 7945 27660 7958
rect 27724 7945 27752 7976
rect 27798 7964 27804 7976
rect 27856 7964 27862 8016
rect 29825 8007 29883 8013
rect 29825 7973 29837 8007
rect 29871 8004 29883 8007
rect 30374 8004 30380 8016
rect 29871 7976 30380 8004
rect 29871 7973 29883 7976
rect 29825 7967 29883 7973
rect 30374 7964 30380 7976
rect 30432 7964 30438 8016
rect 27448 7939 27669 7945
rect 27448 7936 27623 7939
rect 27356 7930 27623 7936
rect 27356 7908 27476 7930
rect 23707 7840 24256 7868
rect 23707 7837 23719 7840
rect 23661 7831 23719 7837
rect 26142 7828 26148 7880
rect 26200 7868 26206 7880
rect 27356 7868 27384 7908
rect 27611 7905 27623 7930
rect 27657 7905 27669 7939
rect 27611 7899 27669 7905
rect 27709 7939 27767 7945
rect 27709 7905 27721 7939
rect 27755 7905 27767 7939
rect 27709 7899 27767 7905
rect 27982 7896 27988 7948
rect 28040 7896 28046 7948
rect 28074 7896 28080 7948
rect 28132 7896 28138 7948
rect 28166 7896 28172 7948
rect 28224 7936 28230 7948
rect 28333 7939 28391 7945
rect 28333 7936 28345 7939
rect 28224 7908 28345 7936
rect 28224 7896 28230 7908
rect 28333 7905 28345 7908
rect 28379 7905 28391 7939
rect 28333 7899 28391 7905
rect 29730 7896 29736 7948
rect 29788 7896 29794 7948
rect 29917 7939 29975 7945
rect 29917 7905 29929 7939
rect 29963 7936 29975 7939
rect 30006 7936 30012 7948
rect 29963 7908 30012 7936
rect 29963 7905 29975 7908
rect 29917 7899 29975 7905
rect 30006 7896 30012 7908
rect 30064 7896 30070 7948
rect 30101 7939 30159 7945
rect 30101 7905 30113 7939
rect 30147 7905 30159 7939
rect 30101 7899 30159 7905
rect 26200 7840 27384 7868
rect 26200 7828 26206 7840
rect 23201 7803 23259 7809
rect 19843 7772 20024 7800
rect 20548 7772 21404 7800
rect 19843 7769 19855 7772
rect 19797 7763 19855 7769
rect 18874 7732 18880 7744
rect 17512 7704 18880 7732
rect 17405 7695 17463 7701
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 18969 7735 19027 7741
rect 18969 7701 18981 7735
rect 19015 7732 19027 7735
rect 20548 7732 20576 7772
rect 19015 7704 20576 7732
rect 19015 7701 19027 7704
rect 18969 7695 19027 7701
rect 20622 7692 20628 7744
rect 20680 7692 20686 7744
rect 21266 7692 21272 7744
rect 21324 7692 21330 7744
rect 21376 7732 21404 7772
rect 23201 7769 23213 7803
rect 23247 7769 23259 7803
rect 23201 7763 23259 7769
rect 23492 7772 24348 7800
rect 23492 7732 23520 7772
rect 21376 7704 23520 7732
rect 23750 7692 23756 7744
rect 23808 7692 23814 7744
rect 24026 7692 24032 7744
rect 24084 7732 24090 7744
rect 24213 7735 24271 7741
rect 24213 7732 24225 7735
rect 24084 7704 24225 7732
rect 24084 7692 24090 7704
rect 24213 7701 24225 7704
rect 24259 7701 24271 7735
rect 24320 7732 24348 7772
rect 24946 7732 24952 7744
rect 24320 7704 24952 7732
rect 24213 7695 24271 7701
rect 24946 7692 24952 7704
rect 25004 7692 25010 7744
rect 26160 7732 26188 7828
rect 26234 7760 26240 7812
rect 26292 7800 26298 7812
rect 27522 7800 27528 7812
rect 26292 7772 27528 7800
rect 26292 7760 26298 7772
rect 27522 7760 27528 7772
rect 27580 7760 27586 7812
rect 27893 7803 27951 7809
rect 27893 7769 27905 7803
rect 27939 7769 27951 7803
rect 27893 7763 27951 7769
rect 27065 7735 27123 7741
rect 27065 7732 27077 7735
rect 26160 7704 27077 7732
rect 27065 7701 27077 7704
rect 27111 7701 27123 7735
rect 27065 7695 27123 7701
rect 27154 7692 27160 7744
rect 27212 7732 27218 7744
rect 27433 7735 27491 7741
rect 27433 7732 27445 7735
rect 27212 7704 27445 7732
rect 27212 7692 27218 7704
rect 27433 7701 27445 7704
rect 27479 7732 27491 7735
rect 27908 7732 27936 7763
rect 27982 7760 27988 7812
rect 28040 7760 28046 7812
rect 29457 7803 29515 7809
rect 29457 7769 29469 7803
rect 29503 7800 29515 7803
rect 30116 7800 30144 7899
rect 30742 7896 30748 7948
rect 30800 7896 30806 7948
rect 31018 7828 31024 7880
rect 31076 7828 31082 7880
rect 29503 7772 30144 7800
rect 29503 7769 29515 7772
rect 29457 7763 29515 7769
rect 27479 7704 27936 7732
rect 27479 7701 27491 7704
rect 27433 7695 27491 7701
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 6178 7488 6184 7540
rect 6236 7488 6242 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6730 7528 6736 7540
rect 6687 7500 6736 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 6917 7531 6975 7537
rect 6917 7528 6929 7531
rect 6880 7500 6929 7528
rect 6880 7488 6886 7500
rect 6917 7497 6929 7500
rect 6963 7497 6975 7531
rect 6917 7491 6975 7497
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 7650 7528 7656 7540
rect 7515 7500 7656 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 10410 7488 10416 7540
rect 10468 7488 10474 7540
rect 10502 7488 10508 7540
rect 10560 7488 10566 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11480 7500 11805 7528
rect 11480 7488 11486 7500
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 11793 7491 11851 7497
rect 14185 7531 14243 7537
rect 14185 7497 14197 7531
rect 14231 7528 14243 7531
rect 15010 7528 15016 7540
rect 14231 7500 15016 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 16114 7488 16120 7540
rect 16172 7528 16178 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 16172 7500 16221 7528
rect 16172 7488 16178 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 16209 7491 16267 7497
rect 16485 7531 16543 7537
rect 16485 7497 16497 7531
rect 16531 7528 16543 7531
rect 16574 7528 16580 7540
rect 16531 7500 16580 7528
rect 16531 7497 16543 7500
rect 16485 7491 16543 7497
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 16945 7531 17003 7537
rect 16945 7497 16957 7531
rect 16991 7528 17003 7531
rect 17310 7528 17316 7540
rect 16991 7500 17316 7528
rect 16991 7497 17003 7500
rect 16945 7491 17003 7497
rect 17310 7488 17316 7500
rect 17368 7528 17374 7540
rect 17862 7528 17868 7540
rect 17368 7500 17868 7528
rect 17368 7488 17374 7500
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 20622 7488 20628 7540
rect 20680 7488 20686 7540
rect 21266 7488 21272 7540
rect 21324 7488 21330 7540
rect 21913 7531 21971 7537
rect 21913 7497 21925 7531
rect 21959 7528 21971 7531
rect 21959 7500 24072 7528
rect 21959 7497 21971 7500
rect 21913 7491 21971 7497
rect 2774 7352 2780 7404
rect 2832 7352 2838 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 3099 7364 3525 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4120 7364 5120 7392
rect 4120 7352 4126 7364
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 2700 7188 2728 7287
rect 3234 7284 3240 7336
rect 3292 7284 3298 7336
rect 5092 7333 5120 7364
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 6196 7324 6224 7488
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7064 7432 7849 7460
rect 7064 7420 7070 7432
rect 7024 7392 7052 7420
rect 6748 7364 6960 7392
rect 7024 7364 7144 7392
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 5123 7296 5488 7324
rect 6196 7296 6653 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 4246 7216 4252 7268
rect 4304 7216 4310 7268
rect 5322 7259 5380 7265
rect 5322 7256 5334 7259
rect 5000 7228 5334 7256
rect 5000 7197 5028 7228
rect 5322 7225 5334 7228
rect 5368 7225 5380 7259
rect 5460 7256 5488 7296
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 6546 7256 6552 7268
rect 5460 7228 6552 7256
rect 5322 7219 5380 7225
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 2700 7160 4997 7188
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 6454 7148 6460 7200
rect 6512 7148 6518 7200
rect 6748 7188 6776 7364
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 6932 7333 6960 7364
rect 7116 7333 7144 7364
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 7331 7296 7420 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 7392 7268 7420 7296
rect 7484 7320 7512 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 17497 7463 17555 7469
rect 17497 7460 17509 7463
rect 9916 7432 10272 7460
rect 9916 7420 9922 7432
rect 8220 7364 8524 7392
rect 8220 7336 8248 7364
rect 7553 7323 7611 7329
rect 7553 7320 7565 7323
rect 7484 7292 7565 7320
rect 7553 7289 7565 7292
rect 7599 7289 7611 7323
rect 7553 7283 7611 7289
rect 7650 7284 7656 7336
rect 7708 7284 7714 7336
rect 8018 7284 8024 7336
rect 8076 7284 8082 7336
rect 8202 7284 8208 7336
rect 8260 7284 8266 7336
rect 8386 7284 8392 7336
rect 8444 7284 8450 7336
rect 8496 7324 8524 7364
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 8496 7296 9873 7324
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 9861 7287 9919 7293
rect 9950 7284 9956 7336
rect 10008 7324 10014 7336
rect 10244 7333 10272 7432
rect 16316 7432 17509 7460
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11664 7364 14504 7392
rect 11664 7352 11670 7364
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 10008 7296 10149 7324
rect 10008 7284 10014 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 10652 7296 10701 7324
rect 10652 7284 10658 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 7374 7216 7380 7268
rect 7432 7216 7438 7268
rect 7668 7256 7696 7284
rect 8634 7259 8692 7265
rect 8634 7256 8646 7259
rect 7668 7228 8646 7256
rect 8634 7225 8646 7228
rect 8680 7225 8692 7259
rect 8634 7219 8692 7225
rect 10042 7216 10048 7268
rect 10100 7216 10106 7268
rect 10704 7256 10732 7287
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11238 7324 11244 7336
rect 11020 7296 11244 7324
rect 11020 7284 11026 7296
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11992 7333 12020 7364
rect 14476 7336 14504 7364
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7324 11759 7327
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11747 7296 11805 7324
rect 11747 7293 11759 7296
rect 11701 7287 11759 7293
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 13538 7284 13544 7336
rect 13596 7284 13602 7336
rect 13630 7284 13636 7336
rect 13688 7284 13694 7336
rect 13814 7284 13820 7336
rect 13872 7284 13878 7336
rect 13998 7284 14004 7336
rect 14056 7333 14062 7336
rect 14056 7324 14064 7333
rect 14056 7296 14101 7324
rect 14056 7287 14064 7296
rect 14056 7284 14062 7287
rect 14458 7284 14464 7336
rect 14516 7284 14522 7336
rect 14826 7284 14832 7336
rect 14884 7284 14890 7336
rect 15096 7327 15154 7333
rect 15096 7293 15108 7327
rect 15142 7324 15154 7327
rect 16316 7324 16344 7432
rect 17497 7429 17509 7432
rect 17543 7429 17555 7463
rect 17497 7423 17555 7429
rect 17678 7420 17684 7472
rect 17736 7460 17742 7472
rect 20530 7460 20536 7472
rect 17736 7432 20536 7460
rect 17736 7420 17742 7432
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 17037 7395 17095 7401
rect 16684 7364 16988 7392
rect 16684 7333 16712 7364
rect 15142 7296 16344 7324
rect 16491 7327 16549 7333
rect 16491 7320 16503 7327
rect 15142 7293 15154 7296
rect 15096 7287 15154 7293
rect 16408 7293 16503 7320
rect 16537 7293 16549 7327
rect 16408 7292 16549 7293
rect 13556 7256 13584 7284
rect 10704 7228 13584 7256
rect 13909 7259 13967 7265
rect 13909 7225 13921 7259
rect 13955 7225 13967 7259
rect 16408 7256 16436 7292
rect 16491 7287 16549 7292
rect 16669 7327 16727 7333
rect 16669 7293 16681 7327
rect 16715 7293 16727 7327
rect 16669 7287 16727 7293
rect 16758 7284 16764 7336
rect 16816 7284 16822 7336
rect 16853 7327 16911 7333
rect 16853 7293 16865 7327
rect 16899 7293 16911 7327
rect 16960 7324 16988 7364
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17083 7364 17877 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 18782 7392 18788 7404
rect 17865 7355 17923 7361
rect 17972 7364 18788 7392
rect 17310 7324 17316 7336
rect 16960 7296 17316 7324
rect 16853 7287 16911 7293
rect 13909 7219 13967 7225
rect 16224 7228 16436 7256
rect 8478 7188 8484 7200
rect 6748 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7188 8542 7200
rect 9030 7188 9036 7200
rect 8536 7160 9036 7188
rect 8536 7148 8542 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 10873 7191 10931 7197
rect 10873 7188 10885 7191
rect 9815 7160 10885 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 10873 7157 10885 7160
rect 10919 7157 10931 7191
rect 10873 7151 10931 7157
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 13924 7188 13952 7219
rect 16224 7200 16252 7228
rect 13780 7160 13952 7188
rect 13780 7148 13786 7160
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14366 7188 14372 7200
rect 14056 7160 14372 7188
rect 14056 7148 14062 7160
rect 14366 7148 14372 7160
rect 14424 7188 14430 7200
rect 16206 7188 16212 7200
rect 14424 7160 16212 7188
rect 14424 7148 14430 7160
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 16868 7188 16896 7287
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 17451 7296 17632 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 17126 7216 17132 7268
rect 17184 7216 17190 7268
rect 17604 7200 17632 7296
rect 17678 7284 17684 7336
rect 17736 7284 17742 7336
rect 17770 7284 17776 7336
rect 17828 7284 17834 7336
rect 17972 7333 18000 7364
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 18046 7284 18052 7336
rect 18104 7284 18110 7336
rect 18708 7333 18736 7364
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7293 18751 7327
rect 18693 7287 18751 7293
rect 18877 7327 18935 7333
rect 18877 7293 18889 7327
rect 18923 7324 18935 7327
rect 19978 7324 19984 7336
rect 18923 7296 19984 7324
rect 18923 7293 18935 7296
rect 18877 7287 18935 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20640 7324 20668 7488
rect 21284 7392 21312 7488
rect 23293 7463 23351 7469
rect 23293 7429 23305 7463
rect 23339 7429 23351 7463
rect 23293 7423 23351 7429
rect 23385 7463 23443 7469
rect 23385 7429 23397 7463
rect 23431 7460 23443 7463
rect 23842 7460 23848 7472
rect 23431 7432 23848 7460
rect 23431 7429 23443 7432
rect 23385 7423 23443 7429
rect 23308 7392 23336 7423
rect 23842 7420 23848 7432
rect 23900 7420 23906 7472
rect 23937 7463 23995 7469
rect 23937 7429 23949 7463
rect 23983 7429 23995 7463
rect 24044 7460 24072 7500
rect 24394 7488 24400 7540
rect 24452 7488 24458 7540
rect 25593 7531 25651 7537
rect 25593 7497 25605 7531
rect 25639 7528 25651 7531
rect 25866 7528 25872 7540
rect 25639 7500 25872 7528
rect 25639 7497 25651 7500
rect 25593 7491 25651 7497
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 28077 7531 28135 7537
rect 28077 7497 28089 7531
rect 28123 7528 28135 7531
rect 28166 7528 28172 7540
rect 28123 7500 28172 7528
rect 28123 7497 28135 7500
rect 28077 7491 28135 7497
rect 28166 7488 28172 7500
rect 28224 7488 28230 7540
rect 30374 7488 30380 7540
rect 30432 7488 30438 7540
rect 26050 7460 26056 7472
rect 24044 7432 26056 7460
rect 23937 7423 23995 7429
rect 21284 7364 21680 7392
rect 21450 7333 21456 7336
rect 21269 7327 21327 7333
rect 21269 7324 21281 7327
rect 20640 7296 21281 7324
rect 21269 7293 21281 7296
rect 21315 7293 21327 7327
rect 21269 7287 21327 7293
rect 21417 7327 21456 7333
rect 21417 7293 21429 7327
rect 21417 7287 21456 7293
rect 21450 7284 21456 7287
rect 21508 7284 21514 7336
rect 21652 7333 21680 7364
rect 23032 7364 23336 7392
rect 23569 7395 23627 7401
rect 21637 7327 21695 7333
rect 21637 7293 21649 7327
rect 21683 7293 21695 7327
rect 21637 7287 21695 7293
rect 21726 7284 21732 7336
rect 21784 7333 21790 7336
rect 21784 7287 21792 7333
rect 21784 7284 21790 7287
rect 20714 7216 20720 7268
rect 20772 7256 20778 7268
rect 21545 7259 21603 7265
rect 21545 7256 21557 7259
rect 20772 7228 21557 7256
rect 20772 7216 20778 7228
rect 21545 7225 21557 7228
rect 21591 7225 21603 7259
rect 23032 7256 23060 7364
rect 23569 7361 23581 7395
rect 23615 7392 23627 7395
rect 23750 7392 23756 7404
rect 23615 7364 23756 7392
rect 23615 7361 23627 7364
rect 23569 7355 23627 7361
rect 23750 7352 23756 7364
rect 23808 7352 23814 7404
rect 23106 7284 23112 7336
rect 23164 7324 23170 7336
rect 23293 7327 23351 7333
rect 23293 7324 23305 7327
rect 23164 7296 23305 7324
rect 23164 7284 23170 7296
rect 23293 7293 23305 7296
rect 23339 7324 23351 7327
rect 23845 7327 23903 7333
rect 23845 7324 23857 7327
rect 23339 7296 23857 7324
rect 23339 7293 23351 7296
rect 23293 7287 23351 7293
rect 23845 7293 23857 7296
rect 23891 7293 23903 7327
rect 23952 7324 23980 7423
rect 26050 7420 26056 7432
rect 26108 7420 26114 7472
rect 24026 7352 24032 7404
rect 24084 7392 24090 7404
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 24084 7364 24133 7392
rect 24084 7352 24090 7364
rect 24121 7361 24133 7364
rect 24167 7361 24179 7395
rect 26329 7395 26387 7401
rect 26329 7392 26341 7395
rect 24121 7355 24179 7361
rect 26068 7364 26341 7392
rect 24213 7327 24271 7333
rect 24213 7324 24225 7327
rect 23952 7296 24225 7324
rect 23845 7287 23903 7293
rect 24213 7293 24225 7296
rect 24259 7293 24271 7327
rect 24213 7287 24271 7293
rect 23934 7256 23940 7268
rect 23032 7228 23940 7256
rect 21545 7219 21603 7225
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 16632 7160 17417 7188
rect 16632 7148 16638 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17405 7151 17463 7157
rect 17586 7148 17592 7200
rect 17644 7148 17650 7200
rect 18782 7148 18788 7200
rect 18840 7148 18846 7200
rect 21560 7188 21588 7219
rect 23934 7216 23940 7228
rect 23992 7256 23998 7268
rect 24228 7256 24256 7287
rect 24946 7284 24952 7336
rect 25004 7284 25010 7336
rect 25038 7284 25044 7336
rect 25096 7284 25102 7336
rect 26068 7333 26096 7364
rect 26329 7361 26341 7364
rect 26375 7361 26387 7395
rect 26329 7355 26387 7361
rect 28994 7352 29000 7404
rect 29052 7352 29058 7404
rect 25455 7327 25513 7333
rect 25455 7293 25467 7327
rect 25501 7324 25513 7327
rect 26053 7327 26111 7333
rect 25501 7296 26004 7324
rect 25501 7293 25513 7296
rect 25455 7287 25513 7293
rect 23992 7228 24256 7256
rect 25225 7259 25283 7265
rect 23992 7216 23998 7228
rect 25225 7225 25237 7259
rect 25271 7225 25283 7259
rect 25225 7219 25283 7225
rect 24854 7188 24860 7200
rect 21560 7160 24860 7188
rect 24854 7148 24860 7160
rect 24912 7188 24918 7200
rect 25240 7188 25268 7219
rect 25314 7216 25320 7268
rect 25372 7216 25378 7268
rect 25976 7256 26004 7296
rect 26053 7293 26065 7327
rect 26099 7293 26111 7327
rect 26053 7287 26111 7293
rect 26234 7284 26240 7336
rect 26292 7284 26298 7336
rect 26418 7284 26424 7336
rect 26476 7324 26482 7336
rect 26970 7324 26976 7336
rect 26476 7296 26976 7324
rect 26476 7284 26482 7296
rect 26970 7284 26976 7296
rect 27028 7284 27034 7336
rect 27154 7284 27160 7336
rect 27212 7324 27218 7336
rect 27893 7327 27951 7333
rect 27893 7324 27905 7327
rect 27212 7296 27905 7324
rect 27212 7284 27218 7296
rect 27893 7293 27905 7296
rect 27939 7293 27951 7327
rect 27893 7287 27951 7293
rect 27982 7284 27988 7336
rect 28040 7324 28046 7336
rect 28169 7327 28227 7333
rect 28169 7324 28181 7327
rect 28040 7296 28181 7324
rect 28040 7284 28046 7296
rect 28169 7293 28181 7296
rect 28215 7293 28227 7327
rect 28169 7287 28227 7293
rect 26436 7256 26464 7284
rect 25976 7228 26464 7256
rect 26602 7216 26608 7268
rect 26660 7256 26666 7268
rect 26697 7259 26755 7265
rect 26697 7256 26709 7259
rect 26660 7228 26709 7256
rect 26660 7216 26666 7228
rect 26697 7225 26709 7228
rect 26743 7256 26755 7259
rect 27246 7256 27252 7268
rect 26743 7228 27252 7256
rect 26743 7225 26755 7228
rect 26697 7219 26755 7225
rect 27246 7216 27252 7228
rect 27304 7256 27310 7268
rect 27341 7259 27399 7265
rect 27341 7256 27353 7259
rect 27304 7228 27353 7256
rect 27304 7216 27310 7228
rect 27341 7225 27353 7228
rect 27387 7225 27399 7259
rect 27341 7219 27399 7225
rect 27706 7216 27712 7268
rect 27764 7216 27770 7268
rect 29242 7259 29300 7265
rect 29242 7256 29254 7259
rect 28368 7228 29254 7256
rect 24912 7160 25268 7188
rect 24912 7148 24918 7160
rect 26142 7148 26148 7200
rect 26200 7148 26206 7200
rect 26786 7148 26792 7200
rect 26844 7148 26850 7200
rect 28368 7197 28396 7228
rect 29242 7225 29254 7228
rect 29288 7225 29300 7259
rect 29242 7219 29300 7225
rect 28353 7191 28411 7197
rect 28353 7157 28365 7191
rect 28399 7157 28411 7191
rect 28353 7151 28411 7157
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 4246 6944 4252 6996
rect 4304 6944 4310 6996
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 7374 6984 7380 6996
rect 6880 6956 7380 6984
rect 6880 6944 6886 6956
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 7469 6987 7527 6993
rect 7469 6953 7481 6987
rect 7515 6984 7527 6987
rect 7515 6956 7972 6984
rect 7515 6953 7527 6956
rect 7469 6947 7527 6953
rect 5442 6916 5448 6928
rect 4356 6888 5448 6916
rect 4356 6857 4384 6888
rect 5442 6876 5448 6888
rect 5500 6916 5506 6928
rect 5500 6888 6224 6916
rect 5500 6876 5506 6888
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 6069 6851 6127 6857
rect 6069 6848 6081 6851
rect 5960 6820 6081 6848
rect 5960 6808 5966 6820
rect 6069 6817 6081 6820
rect 6115 6817 6127 6851
rect 6196 6848 6224 6888
rect 6914 6848 6920 6860
rect 6196 6820 6920 6848
rect 6069 6811 6127 6817
rect 6914 6808 6920 6820
rect 6972 6848 6978 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 6972 6820 7481 6848
rect 6972 6808 6978 6820
rect 7469 6817 7481 6820
rect 7515 6848 7527 6851
rect 7834 6848 7840 6860
rect 7515 6820 7840 6848
rect 7515 6817 7527 6820
rect 7469 6811 7527 6817
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 7944 6857 7972 6956
rect 11330 6944 11336 6996
rect 11388 6944 11394 6996
rect 12713 6987 12771 6993
rect 12713 6953 12725 6987
rect 12759 6984 12771 6987
rect 12759 6956 13676 6984
rect 12759 6953 12771 6956
rect 12713 6947 12771 6953
rect 11348 6916 11376 6944
rect 8404 6888 8800 6916
rect 11348 6888 12848 6916
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6848 7987 6851
rect 8018 6848 8024 6860
rect 7975 6820 8024 6848
rect 7975 6817 7987 6820
rect 7929 6811 7987 6817
rect 8018 6808 8024 6820
rect 8076 6808 8082 6860
rect 8404 6857 8432 6888
rect 8389 6851 8447 6857
rect 8389 6817 8401 6851
rect 8435 6817 8447 6851
rect 8389 6811 8447 6817
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 8662 6808 8668 6860
rect 8720 6808 8726 6860
rect 8772 6857 8800 6888
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6817 8815 6851
rect 8757 6811 8815 6817
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 11425 6851 11483 6857
rect 8987 6820 9904 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9876 6792 9904 6820
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11606 6848 11612 6860
rect 11471 6820 11612 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 11698 6808 11704 6860
rect 11756 6808 11762 6860
rect 12820 6857 12848 6888
rect 13538 6857 13544 6860
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6848 12587 6851
rect 12805 6851 12863 6857
rect 12575 6820 12609 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 12805 6817 12817 6851
rect 12851 6848 12863 6851
rect 13265 6851 13323 6857
rect 12851 6820 13216 6848
rect 12851 6817 12863 6820
rect 12805 6811 12863 6817
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8113 6783 8171 6789
rect 7791 6752 8064 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 5828 6644 5856 6743
rect 7374 6672 7380 6724
rect 7432 6712 7438 6724
rect 7561 6715 7619 6721
rect 7561 6712 7573 6715
rect 7432 6684 7573 6712
rect 7432 6672 7438 6684
rect 7561 6681 7573 6684
rect 7607 6712 7619 6715
rect 7837 6715 7895 6721
rect 7837 6712 7849 6715
rect 7607 6684 7849 6712
rect 7607 6681 7619 6684
rect 7561 6675 7619 6681
rect 7837 6681 7849 6684
rect 7883 6681 7895 6715
rect 8036 6712 8064 6752
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8849 6783 8907 6789
rect 8849 6780 8861 6783
rect 8159 6752 8861 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8849 6749 8861 6752
rect 8895 6749 8907 6783
rect 8849 6743 8907 6749
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 11790 6740 11796 6792
rect 11848 6740 11854 6792
rect 12544 6780 12572 6811
rect 12897 6783 12955 6789
rect 12406 6752 12848 6780
rect 8481 6715 8539 6721
rect 8481 6712 8493 6715
rect 8036 6684 8493 6712
rect 7837 6675 7895 6681
rect 8481 6681 8493 6684
rect 8527 6681 8539 6715
rect 8481 6675 8539 6681
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 12406 6712 12434 6752
rect 12820 6721 12848 6752
rect 12897 6749 12909 6783
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 8720 6684 12434 6712
rect 12805 6715 12863 6721
rect 8720 6672 8726 6684
rect 12805 6681 12817 6715
rect 12851 6681 12863 6715
rect 12805 6675 12863 6681
rect 12912 6656 12940 6743
rect 13078 6740 13084 6792
rect 13136 6740 13142 6792
rect 6546 6644 6552 6656
rect 5828 6616 6552 6644
rect 6546 6604 6552 6616
rect 6604 6644 6610 6656
rect 6822 6644 6828 6656
rect 6604 6616 6828 6644
rect 6604 6604 6610 6616
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 10318 6644 10324 6656
rect 7239 6616 10324 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 11241 6647 11299 6653
rect 11241 6644 11253 6647
rect 11112 6616 11253 6644
rect 11112 6604 11118 6616
rect 11241 6613 11253 6616
rect 11287 6613 11299 6647
rect 11241 6607 11299 6613
rect 11698 6604 11704 6656
rect 11756 6604 11762 6656
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 11940 6616 12081 6644
rect 11940 6604 11946 6616
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12894 6604 12900 6656
rect 12952 6604 12958 6656
rect 13188 6644 13216 6820
rect 13265 6817 13277 6851
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13532 6811 13544 6857
rect 13280 6724 13308 6811
rect 13538 6808 13544 6811
rect 13596 6808 13602 6860
rect 13648 6848 13676 6956
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 16574 6984 16580 6996
rect 14516 6956 16580 6984
rect 14516 6944 14522 6956
rect 16574 6944 16580 6956
rect 16632 6944 16638 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17221 6987 17279 6993
rect 17221 6984 17233 6987
rect 17184 6956 17233 6984
rect 17184 6944 17190 6956
rect 17221 6953 17233 6956
rect 17267 6953 17279 6987
rect 17221 6947 17279 6953
rect 17405 6987 17463 6993
rect 17405 6953 17417 6987
rect 17451 6984 17463 6987
rect 17678 6984 17684 6996
rect 17451 6956 17684 6984
rect 17451 6953 17463 6956
rect 17405 6947 17463 6953
rect 17420 6916 17448 6947
rect 17678 6944 17684 6956
rect 17736 6944 17742 6996
rect 17770 6944 17776 6996
rect 17828 6944 17834 6996
rect 19334 6944 19340 6996
rect 19392 6944 19398 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19797 6987 19855 6993
rect 19797 6984 19809 6987
rect 19576 6956 19809 6984
rect 19576 6944 19582 6956
rect 19797 6953 19809 6956
rect 19843 6953 19855 6987
rect 22833 6987 22891 6993
rect 22833 6984 22845 6987
rect 19797 6947 19855 6953
rect 22756 6956 22845 6984
rect 17328 6888 17448 6916
rect 17696 6916 17724 6944
rect 18049 6919 18107 6925
rect 17696 6888 17908 6916
rect 14642 6848 14648 6860
rect 13648 6820 14648 6848
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 15010 6808 15016 6860
rect 15068 6808 15074 6860
rect 17328 6857 17356 6888
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17313 6851 17371 6857
rect 17313 6817 17325 6851
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 17405 6851 17463 6857
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 17586 6848 17592 6860
rect 17451 6820 17592 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 15286 6780 15292 6792
rect 14660 6752 15292 6780
rect 13262 6672 13268 6724
rect 13320 6672 13326 6724
rect 14660 6721 14688 6752
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 17144 6780 17172 6811
rect 17586 6808 17592 6820
rect 17644 6848 17650 6860
rect 17880 6857 17908 6888
rect 18049 6885 18061 6919
rect 18095 6916 18107 6919
rect 18782 6916 18788 6928
rect 18095 6888 18788 6916
rect 18095 6885 18107 6888
rect 18049 6879 18107 6885
rect 18782 6876 18788 6888
rect 18840 6876 18846 6928
rect 19352 6916 19380 6944
rect 22756 6916 22784 6956
rect 22833 6953 22845 6956
rect 22879 6953 22891 6987
rect 22833 6947 22891 6953
rect 23290 6944 23296 6996
rect 23348 6984 23354 6996
rect 23348 6956 23612 6984
rect 23348 6944 23354 6956
rect 23584 6916 23612 6956
rect 25314 6944 25320 6996
rect 25372 6984 25378 6996
rect 25409 6987 25467 6993
rect 25409 6984 25421 6987
rect 25372 6956 25421 6984
rect 25372 6944 25378 6956
rect 25409 6953 25421 6956
rect 25455 6953 25467 6987
rect 26878 6984 26884 6996
rect 25409 6947 25467 6953
rect 25700 6956 26884 6984
rect 25700 6916 25728 6956
rect 26878 6944 26884 6956
rect 26936 6984 26942 6996
rect 28629 6987 28687 6993
rect 26936 6956 27016 6984
rect 26936 6944 26942 6956
rect 19352 6888 20484 6916
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 17644 6820 17785 6848
rect 17644 6808 17650 6820
rect 17773 6817 17785 6820
rect 17819 6817 17831 6851
rect 17773 6811 17831 6817
rect 17865 6851 17923 6857
rect 17865 6817 17877 6851
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 18138 6808 18144 6860
rect 18196 6808 18202 6860
rect 18673 6851 18731 6857
rect 18673 6848 18685 6851
rect 18340 6820 18685 6848
rect 17144 6752 17632 6780
rect 14645 6715 14703 6721
rect 14645 6681 14657 6715
rect 14691 6681 14703 6715
rect 14645 6675 14703 6681
rect 17497 6715 17555 6721
rect 17497 6681 17509 6715
rect 17543 6681 17555 6715
rect 17604 6712 17632 6752
rect 17678 6740 17684 6792
rect 17736 6740 17742 6792
rect 18046 6780 18052 6792
rect 17788 6752 18052 6780
rect 17788 6712 17816 6752
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 18340 6721 18368 6820
rect 18673 6817 18685 6820
rect 18719 6817 18731 6851
rect 18673 6811 18731 6817
rect 19978 6808 19984 6860
rect 20036 6848 20042 6860
rect 20456 6857 20484 6888
rect 21836 6888 22048 6916
rect 20622 6857 20628 6860
rect 20073 6851 20131 6857
rect 20073 6848 20085 6851
rect 20036 6820 20085 6848
rect 20036 6808 20042 6820
rect 20073 6817 20085 6820
rect 20119 6817 20131 6851
rect 20073 6811 20131 6817
rect 20441 6851 20499 6857
rect 20441 6817 20453 6851
rect 20487 6817 20499 6851
rect 20441 6811 20499 6817
rect 20589 6851 20628 6857
rect 20589 6817 20601 6851
rect 20589 6811 20628 6817
rect 18417 6783 18475 6789
rect 18417 6749 18429 6783
rect 18463 6749 18475 6783
rect 20088 6780 20116 6811
rect 20622 6808 20628 6811
rect 20680 6808 20686 6860
rect 20714 6808 20720 6860
rect 20772 6808 20778 6860
rect 20806 6808 20812 6860
rect 20864 6808 20870 6860
rect 20898 6808 20904 6860
rect 20956 6857 20962 6860
rect 20956 6811 20964 6857
rect 21836 6848 21864 6888
rect 21100 6820 21864 6848
rect 21913 6851 21971 6857
rect 20956 6808 20962 6811
rect 21100 6780 21128 6820
rect 21913 6817 21925 6851
rect 21959 6817 21971 6851
rect 22020 6848 22048 6888
rect 22756 6888 23336 6916
rect 22756 6848 22784 6888
rect 22020 6820 22784 6848
rect 22833 6851 22891 6857
rect 21913 6811 21971 6817
rect 22833 6817 22845 6851
rect 22879 6848 22891 6851
rect 23198 6848 23204 6860
rect 22879 6820 23204 6848
rect 22879 6817 22891 6820
rect 22833 6811 22891 6817
rect 20088 6752 21128 6780
rect 18417 6743 18475 6749
rect 17604 6684 17816 6712
rect 18325 6715 18383 6721
rect 17497 6675 17555 6681
rect 18325 6681 18337 6715
rect 18371 6681 18383 6715
rect 18325 6675 18383 6681
rect 14734 6644 14740 6656
rect 13188 6616 14740 6644
rect 14734 6604 14740 6616
rect 14792 6644 14798 6656
rect 14829 6647 14887 6653
rect 14829 6644 14841 6647
rect 14792 6616 14841 6644
rect 14792 6604 14798 6616
rect 14829 6613 14841 6616
rect 14875 6613 14887 6647
rect 14829 6607 14887 6613
rect 15102 6604 15108 6656
rect 15160 6604 15166 6656
rect 17512 6644 17540 6675
rect 17770 6644 17776 6656
rect 17512 6616 17776 6644
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18432 6644 18460 6743
rect 21726 6740 21732 6792
rect 21784 6740 21790 6792
rect 21085 6715 21143 6721
rect 19352 6684 20484 6712
rect 18598 6644 18604 6656
rect 18432 6616 18604 6644
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 19058 6604 19064 6656
rect 19116 6644 19122 6656
rect 19352 6644 19380 6684
rect 19116 6616 19380 6644
rect 20257 6647 20315 6653
rect 19116 6604 19122 6616
rect 20257 6613 20269 6647
rect 20303 6644 20315 6647
rect 20346 6644 20352 6656
rect 20303 6616 20352 6644
rect 20303 6613 20315 6616
rect 20257 6607 20315 6613
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 20456 6644 20484 6684
rect 21085 6681 21097 6715
rect 21131 6712 21143 6715
rect 21928 6712 21956 6811
rect 23198 6808 23204 6820
rect 23256 6808 23262 6860
rect 23308 6857 23336 6888
rect 23584 6888 25728 6916
rect 23584 6857 23612 6888
rect 23293 6851 23351 6857
rect 23293 6817 23305 6851
rect 23339 6817 23351 6851
rect 23293 6811 23351 6817
rect 23569 6851 23627 6857
rect 23569 6817 23581 6851
rect 23615 6817 23627 6851
rect 23569 6811 23627 6817
rect 23753 6851 23811 6857
rect 23753 6817 23765 6851
rect 23799 6848 23811 6851
rect 23934 6848 23940 6860
rect 23799 6820 23940 6848
rect 23799 6817 23811 6820
rect 23753 6811 23811 6817
rect 23934 6808 23940 6820
rect 23992 6808 23998 6860
rect 24026 6808 24032 6860
rect 24084 6808 24090 6860
rect 24118 6808 24124 6860
rect 24176 6848 24182 6860
rect 25700 6857 25728 6888
rect 25961 6919 26019 6925
rect 25961 6885 25973 6919
rect 26007 6916 26019 6919
rect 26142 6916 26148 6928
rect 26007 6888 26148 6916
rect 26007 6885 26019 6888
rect 25961 6879 26019 6885
rect 26142 6876 26148 6888
rect 26200 6876 26206 6928
rect 24285 6851 24343 6857
rect 24285 6848 24297 6851
rect 24176 6820 24297 6848
rect 24176 6808 24182 6820
rect 24285 6817 24297 6820
rect 24331 6817 24343 6851
rect 24285 6811 24343 6817
rect 25685 6851 25743 6857
rect 25685 6817 25697 6851
rect 25731 6817 25743 6851
rect 25685 6811 25743 6817
rect 25869 6851 25927 6857
rect 25869 6817 25881 6851
rect 25915 6848 25927 6851
rect 26237 6851 26295 6857
rect 25915 6820 26188 6848
rect 25915 6817 25927 6820
rect 25869 6811 25927 6817
rect 22189 6783 22247 6789
rect 22189 6749 22201 6783
rect 22235 6780 22247 6783
rect 22278 6780 22284 6792
rect 22235 6752 22284 6780
rect 22235 6749 22247 6752
rect 22189 6743 22247 6749
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 22738 6740 22744 6792
rect 22796 6740 22802 6792
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6780 23167 6783
rect 23155 6752 23428 6780
rect 23155 6749 23167 6752
rect 23109 6743 23167 6749
rect 21131 6684 21956 6712
rect 22066 6684 22876 6712
rect 21131 6681 21143 6684
rect 21085 6675 21143 6681
rect 22066 6644 22094 6684
rect 20456 6616 22094 6644
rect 22848 6644 22876 6684
rect 22922 6672 22928 6724
rect 22980 6712 22986 6724
rect 23201 6715 23259 6721
rect 23201 6712 23213 6715
rect 22980 6684 23213 6712
rect 22980 6672 22986 6684
rect 23201 6681 23213 6684
rect 23247 6681 23259 6715
rect 23400 6712 23428 6752
rect 23474 6740 23480 6792
rect 23532 6740 23538 6792
rect 26160 6721 26188 6820
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26605 6851 26663 6857
rect 26605 6848 26617 6851
rect 26283 6820 26617 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26605 6817 26617 6820
rect 26651 6848 26663 6851
rect 26786 6848 26792 6860
rect 26651 6820 26792 6848
rect 26651 6817 26663 6820
rect 26605 6811 26663 6817
rect 26786 6808 26792 6820
rect 26844 6808 26850 6860
rect 26988 6857 27016 6956
rect 28629 6953 28641 6987
rect 28675 6953 28687 6987
rect 28629 6947 28687 6953
rect 27246 6876 27252 6928
rect 27304 6916 27310 6928
rect 27494 6919 27552 6925
rect 27494 6916 27506 6919
rect 27304 6888 27506 6916
rect 27304 6876 27310 6888
rect 27494 6885 27506 6888
rect 27540 6885 27552 6919
rect 28644 6916 28672 6947
rect 28997 6919 29055 6925
rect 28644 6888 28856 6916
rect 27494 6879 27552 6885
rect 26973 6851 27031 6857
rect 26973 6817 26985 6851
rect 27019 6817 27031 6851
rect 26973 6811 27031 6817
rect 27154 6808 27160 6860
rect 27212 6808 27218 6860
rect 28074 6848 28080 6860
rect 27264 6820 28080 6848
rect 26418 6740 26424 6792
rect 26476 6780 26482 6792
rect 27264 6789 27292 6820
rect 28074 6808 28080 6820
rect 28132 6808 28138 6860
rect 28718 6808 28724 6860
rect 28776 6808 28782 6860
rect 28828 6857 28856 6888
rect 28997 6885 29009 6919
rect 29043 6916 29055 6919
rect 30006 6916 30012 6928
rect 29043 6888 30012 6916
rect 29043 6885 29055 6888
rect 28997 6879 29055 6885
rect 30006 6876 30012 6888
rect 30064 6876 30070 6928
rect 28814 6851 28872 6857
rect 28814 6817 28826 6851
rect 28860 6817 28872 6851
rect 28814 6811 28872 6817
rect 29086 6808 29092 6860
rect 29144 6808 29150 6860
rect 29227 6851 29285 6857
rect 29227 6817 29239 6851
rect 29273 6848 29285 6851
rect 29730 6848 29736 6860
rect 29273 6820 29736 6848
rect 29273 6817 29285 6820
rect 29227 6811 29285 6817
rect 29730 6808 29736 6820
rect 29788 6808 29794 6860
rect 26881 6783 26939 6789
rect 26476 6752 26832 6780
rect 26476 6740 26482 6752
rect 23569 6715 23627 6721
rect 23569 6712 23581 6715
rect 23400 6684 23581 6712
rect 23201 6675 23259 6681
rect 23569 6681 23581 6684
rect 23615 6681 23627 6715
rect 23569 6675 23627 6681
rect 26145 6715 26203 6721
rect 26145 6681 26157 6715
rect 26191 6681 26203 6715
rect 26145 6675 26203 6681
rect 26237 6715 26295 6721
rect 26237 6681 26249 6715
rect 26283 6712 26295 6715
rect 26694 6712 26700 6724
rect 26283 6684 26700 6712
rect 26283 6681 26295 6684
rect 26237 6675 26295 6681
rect 25685 6647 25743 6653
rect 25685 6644 25697 6647
rect 22848 6616 25697 6644
rect 25685 6613 25697 6616
rect 25731 6613 25743 6647
rect 26160 6644 26188 6675
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 26804 6712 26832 6752
rect 26881 6749 26893 6783
rect 26927 6780 26939 6783
rect 27065 6783 27123 6789
rect 27065 6780 27077 6783
rect 26927 6752 27077 6780
rect 26927 6749 26939 6752
rect 26881 6743 26939 6749
rect 27065 6749 27077 6752
rect 27111 6749 27123 6783
rect 27065 6743 27123 6749
rect 27249 6783 27307 6789
rect 27249 6749 27261 6783
rect 27295 6749 27307 6783
rect 27249 6743 27307 6749
rect 27264 6712 27292 6743
rect 26804 6684 27292 6712
rect 29362 6672 29368 6724
rect 29420 6672 29426 6724
rect 26789 6647 26847 6653
rect 26789 6644 26801 6647
rect 26160 6616 26801 6644
rect 25685 6607 25743 6613
rect 26789 6613 26801 6616
rect 26835 6644 26847 6647
rect 27154 6644 27160 6656
rect 26835 6616 27160 6644
rect 26835 6613 26847 6616
rect 26789 6607 26847 6613
rect 27154 6604 27160 6616
rect 27212 6604 27218 6656
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 9858 6440 9864 6452
rect 8680 6412 9864 6440
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5123 6276 5764 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 3326 6196 3332 6248
rect 3384 6196 3390 6248
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6236 5411 6239
rect 5442 6236 5448 6248
rect 5399 6208 5448 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5736 6245 5764 6276
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 5810 6236 5816 6248
rect 5767 6208 5816 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 5810 6196 5816 6208
rect 5868 6236 5874 6248
rect 5868 6208 6132 6236
rect 5868 6196 5874 6208
rect 3602 6128 3608 6180
rect 3660 6128 3666 6180
rect 5261 6171 5319 6177
rect 5261 6168 5273 6171
rect 4830 6140 5273 6168
rect 5261 6137 5273 6140
rect 5307 6137 5319 6171
rect 5261 6131 5319 6137
rect 5902 6128 5908 6180
rect 5960 6128 5966 6180
rect 5994 6128 6000 6180
rect 6052 6128 6058 6180
rect 6104 6168 6132 6208
rect 6822 6196 6828 6248
rect 6880 6196 6886 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8680 6236 8708 6412
rect 9858 6400 9864 6412
rect 9916 6440 9922 6452
rect 9916 6412 11744 6440
rect 9916 6400 9922 6412
rect 11716 6372 11744 6412
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 11848 6412 12265 6440
rect 11848 6400 11854 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 12253 6403 12311 6409
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 13136 6412 13185 6440
rect 13136 6400 13142 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 13538 6400 13544 6452
rect 13596 6400 13602 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 13648 6412 14565 6440
rect 12894 6372 12900 6384
rect 11716 6344 12900 6372
rect 12894 6332 12900 6344
rect 12952 6372 12958 6384
rect 13648 6372 13676 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 14660 6412 16252 6440
rect 14660 6372 14688 6412
rect 12952 6344 13676 6372
rect 14108 6344 14688 6372
rect 12952 6332 12958 6344
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 12986 6304 12992 6316
rect 12452 6276 12992 6304
rect 11054 6245 11060 6248
rect 8527 6208 8708 6236
rect 10781 6239 10839 6245
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 10781 6205 10793 6239
rect 10827 6205 10839 6239
rect 11048 6236 11060 6245
rect 11015 6208 11060 6236
rect 10781 6199 10839 6205
rect 11048 6199 11060 6208
rect 7070 6171 7128 6177
rect 7070 6168 7082 6171
rect 6104 6140 7082 6168
rect 7070 6137 7082 6140
rect 7116 6137 7128 6171
rect 9002 6171 9060 6177
rect 9002 6168 9014 6171
rect 7070 6131 7128 6137
rect 8680 6140 9014 6168
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 3568 6072 5457 6100
rect 3568 6060 3574 6072
rect 5445 6069 5457 6072
rect 5491 6069 5503 6103
rect 5445 6063 5503 6069
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 5718 6100 5724 6112
rect 5675 6072 5724 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5813 6103 5871 6109
rect 5813 6069 5825 6103
rect 5859 6100 5871 6103
rect 5920 6100 5948 6128
rect 5859 6072 5948 6100
rect 8205 6103 8263 6109
rect 5859 6069 5871 6072
rect 5813 6063 5871 6069
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8570 6100 8576 6112
rect 8251 6072 8576 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 8680 6109 8708 6140
rect 9002 6137 9014 6140
rect 9048 6137 9060 6171
rect 10796 6168 10824 6199
rect 11054 6196 11060 6199
rect 11112 6196 11118 6248
rect 11514 6196 11520 6248
rect 11572 6196 11578 6248
rect 12452 6245 12480 6276
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13998 6304 14004 6316
rect 13188 6276 14004 6304
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 13188 6245 13216 6276
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12768 6208 12817 6236
rect 12768 6196 12774 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13403 6208 13737 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 13725 6205 13737 6208
rect 13771 6236 13783 6239
rect 14108 6236 14136 6344
rect 15194 6332 15200 6384
rect 15252 6332 15258 6384
rect 16224 6372 16252 6412
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 16448 6412 16681 6440
rect 16448 6400 16454 6412
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 16669 6403 16727 6409
rect 16758 6400 16764 6452
rect 16816 6440 16822 6452
rect 17586 6440 17592 6452
rect 16816 6412 17592 6440
rect 16816 6400 16822 6412
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 18656 6412 19334 6440
rect 18656 6400 18662 6412
rect 18693 6375 18751 6381
rect 18693 6372 18705 6375
rect 16224 6344 18705 6372
rect 18693 6341 18705 6344
rect 18739 6372 18751 6375
rect 19153 6375 19211 6381
rect 19153 6372 19165 6375
rect 18739 6344 19165 6372
rect 18739 6341 18751 6344
rect 18693 6335 18751 6341
rect 19153 6341 19165 6344
rect 19199 6341 19211 6375
rect 19306 6372 19334 6412
rect 20806 6400 20812 6452
rect 20864 6440 20870 6452
rect 21453 6443 21511 6449
rect 21453 6440 21465 6443
rect 20864 6412 21465 6440
rect 20864 6400 20870 6412
rect 21453 6409 21465 6412
rect 21499 6409 21511 6443
rect 21453 6403 21511 6409
rect 23474 6400 23480 6452
rect 23532 6400 23538 6452
rect 24029 6443 24087 6449
rect 24029 6409 24041 6443
rect 24075 6440 24087 6443
rect 24118 6440 24124 6452
rect 24075 6412 24124 6440
rect 24075 6409 24087 6412
rect 24029 6403 24087 6409
rect 24118 6400 24124 6412
rect 24176 6400 24182 6452
rect 24673 6443 24731 6449
rect 24673 6409 24685 6443
rect 24719 6440 24731 6443
rect 25222 6440 25228 6452
rect 24719 6412 25228 6440
rect 24719 6409 24731 6412
rect 24673 6403 24731 6409
rect 25222 6400 25228 6412
rect 25280 6400 25286 6452
rect 25958 6400 25964 6452
rect 26016 6440 26022 6452
rect 26881 6443 26939 6449
rect 26881 6440 26893 6443
rect 26016 6412 26893 6440
rect 26016 6400 26022 6412
rect 26881 6409 26893 6412
rect 26927 6409 26939 6443
rect 26881 6403 26939 6409
rect 27246 6400 27252 6452
rect 27304 6440 27310 6452
rect 27341 6443 27399 6449
rect 27341 6440 27353 6443
rect 27304 6412 27353 6440
rect 27304 6400 27310 6412
rect 27341 6409 27353 6412
rect 27387 6409 27399 6443
rect 27341 6403 27399 6409
rect 28718 6400 28724 6452
rect 28776 6400 28782 6452
rect 26789 6375 26847 6381
rect 19306 6344 20116 6372
rect 19153 6335 19211 6341
rect 15102 6304 15108 6316
rect 14384 6276 15108 6304
rect 14384 6245 14412 6276
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15212 6276 15424 6304
rect 13771 6208 14136 6236
rect 14185 6239 14243 6245
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 11532 6168 11560 6196
rect 12529 6171 12587 6177
rect 12529 6168 12541 6171
rect 10796 6140 11560 6168
rect 12176 6140 12541 6168
rect 9002 6131 9060 6137
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6069 8723 6103
rect 8665 6063 8723 6069
rect 10134 6060 10140 6112
rect 10192 6060 10198 6112
rect 12176 6109 12204 6140
rect 12529 6137 12541 6140
rect 12575 6137 12587 6171
rect 12529 6131 12587 6137
rect 12621 6171 12679 6177
rect 12621 6137 12633 6171
rect 12667 6168 12679 6171
rect 14090 6168 14096 6180
rect 12667 6140 14096 6168
rect 12667 6137 12679 6140
rect 12621 6131 12679 6137
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 12161 6103 12219 6109
rect 12161 6069 12173 6103
rect 12207 6069 12219 6103
rect 14200 6100 14228 6199
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 14734 6196 14740 6248
rect 14792 6196 14798 6248
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6236 15071 6239
rect 15212 6236 15240 6276
rect 15059 6208 15240 6236
rect 15059 6205 15071 6208
rect 15013 6199 15071 6205
rect 14277 6171 14335 6177
rect 14277 6137 14289 6171
rect 14323 6168 14335 6171
rect 14461 6171 14519 6177
rect 14461 6168 14473 6171
rect 14323 6140 14473 6168
rect 14323 6137 14335 6140
rect 14277 6131 14335 6137
rect 14461 6137 14473 6140
rect 14507 6137 14519 6171
rect 15028 6168 15056 6199
rect 15286 6196 15292 6248
rect 15344 6196 15350 6248
rect 15396 6236 15424 6276
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 20088 6313 20116 6344
rect 26789 6341 26801 6375
rect 26835 6372 26847 6375
rect 28736 6372 28764 6400
rect 26835 6344 28764 6372
rect 26835 6341 26847 6344
rect 26789 6335 26847 6341
rect 20073 6307 20131 6313
rect 17736 6276 19288 6304
rect 17736 6264 17742 6276
rect 15396 6208 16804 6236
rect 14461 6131 14519 6137
rect 14568 6140 15056 6168
rect 14568 6100 14596 6140
rect 15194 6128 15200 6180
rect 15252 6168 15258 6180
rect 15534 6171 15592 6177
rect 15534 6168 15546 6171
rect 15252 6140 15546 6168
rect 15252 6128 15258 6140
rect 15534 6137 15546 6140
rect 15580 6137 15592 6171
rect 16776 6168 16804 6208
rect 18690 6196 18696 6248
rect 18748 6196 18754 6248
rect 18785 6239 18843 6245
rect 18785 6205 18797 6239
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 18800 6168 18828 6199
rect 18966 6196 18972 6248
rect 19024 6196 19030 6248
rect 19061 6239 19119 6245
rect 19061 6205 19073 6239
rect 19107 6236 19119 6239
rect 19107 6208 19196 6236
rect 19107 6205 19119 6208
rect 19061 6199 19119 6205
rect 16776 6140 19104 6168
rect 15534 6131 15592 6137
rect 14200 6072 14596 6100
rect 12161 6063 12219 6069
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 18138 6100 18144 6112
rect 14700 6072 18144 6100
rect 14700 6060 14706 6072
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 19076 6109 19104 6140
rect 19168 6112 19196 6208
rect 19061 6103 19119 6109
rect 19061 6069 19073 6103
rect 19107 6069 19119 6103
rect 19061 6063 19119 6069
rect 19150 6060 19156 6112
rect 19208 6060 19214 6112
rect 19260 6100 19288 6276
rect 20073 6273 20085 6307
rect 20119 6273 20131 6307
rect 24854 6304 24860 6316
rect 20073 6267 20131 6273
rect 22066 6276 24348 6304
rect 20346 6245 20352 6248
rect 20340 6236 20352 6245
rect 20307 6208 20352 6236
rect 20340 6199 20352 6208
rect 20346 6196 20352 6199
rect 20404 6196 20410 6248
rect 20714 6196 20720 6248
rect 20772 6236 20778 6248
rect 22066 6236 22094 6276
rect 20772 6208 22094 6236
rect 22557 6239 22615 6245
rect 20772 6196 20778 6208
rect 22557 6205 22569 6239
rect 22603 6236 22615 6239
rect 22649 6239 22707 6245
rect 22649 6236 22661 6239
rect 22603 6208 22661 6236
rect 22603 6205 22615 6208
rect 22557 6199 22615 6205
rect 22649 6205 22661 6208
rect 22695 6205 22707 6239
rect 22649 6199 22707 6205
rect 22833 6239 22891 6245
rect 22833 6205 22845 6239
rect 22879 6236 22891 6239
rect 22922 6236 22928 6248
rect 22879 6208 22928 6236
rect 22879 6205 22891 6208
rect 22833 6199 22891 6205
rect 22922 6196 22928 6208
rect 22980 6196 22986 6248
rect 23385 6239 23443 6245
rect 23385 6205 23397 6239
rect 23431 6236 23443 6239
rect 23477 6239 23535 6245
rect 23477 6236 23489 6239
rect 23431 6208 23489 6236
rect 23431 6205 23443 6208
rect 23385 6199 23443 6205
rect 23477 6205 23489 6208
rect 23523 6205 23535 6239
rect 23477 6199 23535 6205
rect 23661 6239 23719 6245
rect 23661 6205 23673 6239
rect 23707 6236 23719 6239
rect 23842 6236 23848 6248
rect 23707 6208 23848 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 23842 6196 23848 6208
rect 23900 6196 23906 6248
rect 24118 6196 24124 6248
rect 24176 6196 24182 6248
rect 24320 6245 24348 6276
rect 24826 6264 24860 6304
rect 24912 6304 24918 6316
rect 24912 6276 26464 6304
rect 24912 6264 24918 6276
rect 24305 6239 24363 6245
rect 24305 6205 24317 6239
rect 24351 6205 24363 6239
rect 24305 6199 24363 6205
rect 24489 6239 24547 6245
rect 24489 6205 24501 6239
rect 24535 6236 24547 6239
rect 24826 6236 24854 6264
rect 24535 6208 24854 6236
rect 24535 6205 24547 6208
rect 24489 6199 24547 6205
rect 25958 6196 25964 6248
rect 26016 6196 26022 6248
rect 26145 6239 26203 6245
rect 26145 6205 26157 6239
rect 26191 6205 26203 6239
rect 26145 6199 26203 6205
rect 19337 6171 19395 6177
rect 19337 6137 19349 6171
rect 19383 6168 19395 6171
rect 19383 6140 24072 6168
rect 19383 6137 19395 6140
rect 19337 6131 19395 6137
rect 22741 6103 22799 6109
rect 22741 6100 22753 6103
rect 19260 6072 22753 6100
rect 22741 6069 22753 6072
rect 22787 6069 22799 6103
rect 22741 6063 22799 6069
rect 23106 6060 23112 6112
rect 23164 6060 23170 6112
rect 24044 6100 24072 6140
rect 24394 6128 24400 6180
rect 24452 6128 24458 6180
rect 26053 6171 26111 6177
rect 26053 6168 26065 6171
rect 24504 6140 26065 6168
rect 24504 6100 24532 6140
rect 26053 6137 26065 6140
rect 26099 6137 26111 6171
rect 26053 6131 26111 6137
rect 24044 6072 24532 6100
rect 26160 6100 26188 6199
rect 26234 6196 26240 6248
rect 26292 6196 26298 6248
rect 26436 6245 26464 6276
rect 26421 6239 26479 6245
rect 26421 6205 26433 6239
rect 26467 6205 26479 6239
rect 26421 6199 26479 6205
rect 26605 6239 26663 6245
rect 26605 6205 26617 6239
rect 26651 6236 26663 6239
rect 26970 6236 26976 6248
rect 26651 6208 26976 6236
rect 26651 6205 26663 6208
rect 26605 6199 26663 6205
rect 26970 6196 26976 6208
rect 27028 6196 27034 6248
rect 27154 6196 27160 6248
rect 27212 6196 27218 6248
rect 26510 6128 26516 6180
rect 26568 6128 26574 6180
rect 26694 6100 26700 6112
rect 26160 6072 26700 6100
rect 26694 6060 26700 6072
rect 26752 6060 26758 6112
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 3602 5856 3608 5908
rect 3660 5856 3666 5908
rect 5810 5856 5816 5908
rect 5868 5856 5874 5908
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 5960 5868 6101 5896
rect 5960 5856 5966 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10192 5868 10272 5896
rect 10192 5856 10198 5868
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 3510 5760 3516 5772
rect 2832 5732 3516 5760
rect 2832 5720 2838 5732
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 5828 5769 5856 5856
rect 3697 5763 3755 5769
rect 3697 5729 3709 5763
rect 3743 5729 3755 5763
rect 3697 5723 3755 5729
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5729 5871 5763
rect 5813 5723 5871 5729
rect 6181 5763 6239 5769
rect 6181 5729 6193 5763
rect 6227 5760 6239 5763
rect 8588 5760 8616 5856
rect 10244 5837 10272 5868
rect 10318 5856 10324 5908
rect 10376 5856 10382 5908
rect 10505 5899 10563 5905
rect 10505 5865 10517 5899
rect 10551 5896 10563 5899
rect 11698 5896 11704 5908
rect 10551 5868 11704 5896
rect 10551 5865 10563 5868
rect 10505 5859 10563 5865
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 12802 5856 12808 5908
rect 12860 5856 12866 5908
rect 17586 5896 17592 5908
rect 16316 5868 17592 5896
rect 10229 5831 10287 5837
rect 10229 5797 10241 5831
rect 10275 5797 10287 5831
rect 10336 5828 10364 5856
rect 13940 5831 13998 5837
rect 10336 5800 12434 5828
rect 10229 5791 10287 5797
rect 9953 5763 10011 5769
rect 9953 5760 9965 5763
rect 6227 5732 6684 5760
rect 8588 5732 9965 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 3712 5692 3740 5723
rect 3712 5664 5856 5692
rect 5828 5633 5856 5664
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 5813 5627 5871 5633
rect 5813 5593 5825 5627
rect 5859 5593 5871 5627
rect 5813 5587 5871 5593
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 6196 5556 6224 5723
rect 6656 5704 6684 5732
rect 9953 5729 9965 5732
rect 9999 5729 10011 5763
rect 9953 5723 10011 5729
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 10321 5763 10379 5769
rect 10183 5732 10272 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 10244 5704 10272 5732
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10962 5760 10968 5772
rect 10367 5732 10968 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 12406 5760 12434 5800
rect 13940 5797 13952 5831
rect 13986 5828 13998 5831
rect 13986 5800 16252 5828
rect 13986 5797 13998 5800
rect 13940 5791 13998 5797
rect 13630 5760 13636 5772
rect 12406 5732 13636 5760
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 14090 5720 14096 5772
rect 14148 5760 14154 5772
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14148 5732 14749 5760
rect 14148 5720 14154 5732
rect 14737 5729 14749 5732
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 15102 5720 15108 5772
rect 15160 5720 15166 5772
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 14185 5695 14243 5701
rect 14185 5661 14197 5695
rect 14231 5661 14243 5695
rect 14185 5655 14243 5661
rect 14200 5624 14228 5655
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 14332 5664 14473 5692
rect 14332 5652 14338 5664
rect 14461 5661 14473 5664
rect 14507 5692 14519 5695
rect 16224 5692 16252 5800
rect 16316 5769 16344 5868
rect 17586 5856 17592 5868
rect 17644 5896 17650 5908
rect 17862 5896 17868 5908
rect 17644 5868 17868 5896
rect 17644 5856 17650 5868
rect 17862 5856 17868 5868
rect 17920 5896 17926 5908
rect 17920 5868 18092 5896
rect 17920 5856 17926 5868
rect 18064 5828 18092 5868
rect 18230 5856 18236 5908
rect 18288 5856 18294 5908
rect 20622 5856 20628 5908
rect 20680 5896 20686 5908
rect 20809 5899 20867 5905
rect 20809 5896 20821 5899
rect 20680 5868 20821 5896
rect 20680 5856 20686 5868
rect 20809 5865 20821 5868
rect 20855 5865 20867 5899
rect 20809 5859 20867 5865
rect 23106 5856 23112 5908
rect 23164 5856 23170 5908
rect 23201 5899 23259 5905
rect 23201 5865 23213 5899
rect 23247 5896 23259 5899
rect 24118 5896 24124 5908
rect 23247 5868 24124 5896
rect 23247 5865 23259 5868
rect 23201 5859 23259 5865
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 24394 5856 24400 5908
rect 24452 5896 24458 5908
rect 24673 5899 24731 5905
rect 24673 5896 24685 5899
rect 24452 5868 24685 5896
rect 24452 5856 24458 5868
rect 24673 5865 24685 5868
rect 24719 5865 24731 5899
rect 24673 5859 24731 5865
rect 26145 5899 26203 5905
rect 26145 5865 26157 5899
rect 26191 5896 26203 5899
rect 26510 5896 26516 5908
rect 26191 5868 26516 5896
rect 26191 5865 26203 5868
rect 26145 5859 26203 5865
rect 26510 5856 26516 5868
rect 26568 5856 26574 5908
rect 27249 5899 27307 5905
rect 27249 5865 27261 5899
rect 27295 5865 27307 5899
rect 27249 5859 27307 5865
rect 28721 5899 28779 5905
rect 28721 5865 28733 5899
rect 28767 5896 28779 5899
rect 29086 5896 29092 5908
rect 28767 5868 29092 5896
rect 28767 5865 28779 5868
rect 28721 5859 28779 5865
rect 18690 5828 18696 5840
rect 16868 5800 17264 5828
rect 18064 5800 18696 5828
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5729 16359 5763
rect 16758 5760 16764 5772
rect 16301 5723 16359 5729
rect 16408 5732 16764 5760
rect 16408 5692 16436 5732
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 16868 5769 16896 5800
rect 16853 5763 16911 5769
rect 16853 5729 16865 5763
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17109 5763 17167 5769
rect 17109 5760 17121 5763
rect 17000 5732 17121 5760
rect 17000 5720 17006 5732
rect 17109 5729 17121 5732
rect 17155 5729 17167 5763
rect 17236 5760 17264 5800
rect 18690 5788 18696 5800
rect 18748 5828 18754 5840
rect 19150 5828 19156 5840
rect 18748 5800 19156 5828
rect 18748 5788 18754 5800
rect 19150 5788 19156 5800
rect 19208 5828 19214 5840
rect 23124 5828 23152 5856
rect 25010 5831 25068 5837
rect 25010 5828 25022 5831
rect 19208 5800 23060 5828
rect 23124 5800 25022 5828
rect 19208 5788 19214 5800
rect 18598 5760 18604 5772
rect 17236 5732 18604 5760
rect 17109 5723 17167 5729
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 22094 5769 22100 5772
rect 19685 5763 19743 5769
rect 19685 5760 19697 5763
rect 19392 5732 19697 5760
rect 19392 5720 19398 5732
rect 19685 5729 19697 5732
rect 19731 5729 19743 5763
rect 19685 5723 19743 5729
rect 22077 5763 22100 5769
rect 22077 5729 22089 5763
rect 22077 5723 22100 5729
rect 22094 5720 22100 5723
rect 22152 5720 22158 5772
rect 14507 5664 15608 5692
rect 16224 5664 16436 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 14826 5624 14832 5636
rect 14200 5596 14832 5624
rect 5776 5528 6224 5556
rect 5776 5516 5782 5528
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 13262 5556 13268 5568
rect 11572 5528 13268 5556
rect 11572 5516 11578 5528
rect 13262 5516 13268 5528
rect 13320 5556 13326 5568
rect 14200 5556 14228 5596
rect 14826 5584 14832 5596
rect 14884 5624 14890 5636
rect 15286 5624 15292 5636
rect 14884 5596 15292 5624
rect 14884 5584 14890 5596
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 15580 5624 15608 5664
rect 16482 5652 16488 5704
rect 16540 5652 16546 5704
rect 18616 5692 18644 5720
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 18616 5664 19441 5692
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 19429 5655 19487 5661
rect 20456 5664 21833 5692
rect 16500 5624 16528 5652
rect 15580 5596 16528 5624
rect 13320 5528 14228 5556
rect 13320 5516 13326 5528
rect 14550 5516 14556 5568
rect 14608 5516 14614 5568
rect 14921 5559 14979 5565
rect 14921 5525 14933 5559
rect 14967 5556 14979 5559
rect 15010 5556 15016 5568
rect 14967 5528 15016 5556
rect 14967 5525 14979 5528
rect 14921 5519 14979 5525
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 15197 5559 15255 5565
rect 15197 5525 15209 5559
rect 15243 5556 15255 5559
rect 15654 5556 15660 5568
rect 15243 5528 15660 5556
rect 15243 5525 15255 5528
rect 15197 5519 15255 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16206 5516 16212 5568
rect 16264 5516 16270 5568
rect 19444 5556 19472 5655
rect 20456 5556 20484 5664
rect 21821 5661 21833 5664
rect 21867 5661 21879 5695
rect 21821 5655 21879 5661
rect 19444 5528 20484 5556
rect 23032 5556 23060 5800
rect 25010 5797 25022 5800
rect 25056 5797 25068 5831
rect 27264 5828 27292 5859
rect 29086 5856 29092 5868
rect 29144 5856 29150 5908
rect 27586 5831 27644 5837
rect 27586 5828 27598 5831
rect 27264 5800 27598 5828
rect 25010 5791 25068 5797
rect 27586 5797 27598 5800
rect 27632 5797 27644 5831
rect 27586 5791 27644 5797
rect 23293 5763 23351 5769
rect 23293 5729 23305 5763
rect 23339 5760 23351 5763
rect 23382 5760 23388 5772
rect 23339 5732 23388 5760
rect 23339 5729 23351 5732
rect 23293 5723 23351 5729
rect 23382 5720 23388 5732
rect 23440 5720 23446 5772
rect 23560 5763 23618 5769
rect 23560 5729 23572 5763
rect 23606 5760 23618 5763
rect 23934 5760 23940 5772
rect 23606 5732 23940 5760
rect 23606 5729 23618 5732
rect 23560 5723 23618 5729
rect 23934 5720 23940 5732
rect 23992 5720 23998 5772
rect 24026 5720 24032 5772
rect 24084 5760 24090 5772
rect 24765 5763 24823 5769
rect 24765 5760 24777 5763
rect 24084 5732 24777 5760
rect 24084 5720 24090 5732
rect 24765 5729 24777 5732
rect 24811 5760 24823 5763
rect 26418 5760 26424 5772
rect 24811 5732 26424 5760
rect 24811 5729 24823 5732
rect 24765 5723 24823 5729
rect 26418 5720 26424 5732
rect 26476 5720 26482 5772
rect 26694 5720 26700 5772
rect 26752 5760 26758 5772
rect 27065 5763 27123 5769
rect 27065 5760 27077 5763
rect 26752 5732 27077 5760
rect 26752 5720 26758 5732
rect 27065 5729 27077 5732
rect 27111 5729 27123 5763
rect 27065 5723 27123 5729
rect 27338 5720 27344 5772
rect 27396 5760 27402 5772
rect 28994 5760 29000 5772
rect 27396 5732 29000 5760
rect 27396 5720 27402 5732
rect 28994 5720 29000 5732
rect 29052 5720 29058 5772
rect 26602 5556 26608 5568
rect 23032 5528 26608 5556
rect 26602 5516 26608 5528
rect 26660 5516 26666 5568
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 5902 5312 5908 5364
rect 5960 5312 5966 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 6880 5324 7420 5352
rect 6880 5312 6886 5324
rect 5920 5284 5948 5312
rect 6086 5284 6092 5296
rect 5920 5256 6092 5284
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 4062 5216 4068 5228
rect 3384 5188 4068 5216
rect 3384 5176 3390 5188
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5920 5216 5948 5256
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 6638 5284 6644 5296
rect 6564 5256 6644 5284
rect 6564 5225 6592 5256
rect 6638 5244 6644 5256
rect 6696 5284 6702 5296
rect 6696 5256 7328 5284
rect 6696 5244 6702 5256
rect 7300 5228 7328 5256
rect 5123 5188 5948 5216
rect 6549 5219 6607 5225
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5552 5157 5580 5188
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5776 5120 5825 5148
rect 5776 5108 5782 5120
rect 5813 5117 5825 5120
rect 5859 5117 5871 5151
rect 5813 5111 5871 5117
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 5960 5120 6040 5148
rect 5960 5108 5966 5120
rect 3602 5040 3608 5092
rect 3660 5040 3666 5092
rect 4338 5040 4344 5092
rect 4396 5040 4402 5092
rect 6012 5080 6040 5120
rect 6086 5108 6092 5160
rect 6144 5108 6150 5160
rect 6454 5108 6460 5160
rect 6512 5108 6518 5160
rect 7190 5108 7196 5160
rect 7248 5108 7254 5160
rect 6472 5080 6500 5108
rect 6012 5052 6500 5080
rect 7392 5080 7420 5324
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8938 5352 8944 5364
rect 7892 5324 8944 5352
rect 7892 5312 7898 5324
rect 7944 5157 7972 5324
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9950 5312 9956 5364
rect 10008 5312 10014 5364
rect 11425 5355 11483 5361
rect 11425 5321 11437 5355
rect 11471 5352 11483 5355
rect 12710 5352 12716 5364
rect 11471 5324 12716 5352
rect 11471 5321 11483 5324
rect 11425 5315 11483 5321
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 13170 5312 13176 5364
rect 13228 5312 13234 5364
rect 14200 5324 16436 5352
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 11572 5188 11805 5216
rect 11572 5176 11578 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5117 8631 5151
rect 8829 5151 8887 5157
rect 8829 5148 8841 5151
rect 8573 5111 8631 5117
rect 8772 5120 8841 5148
rect 8588 5080 8616 5111
rect 7392 5052 8616 5080
rect 8772 5024 8800 5120
rect 8829 5117 8841 5120
rect 8875 5117 8887 5151
rect 8829 5111 8887 5117
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 11532 5148 11560 5176
rect 14200 5148 14228 5324
rect 16206 5244 16212 5296
rect 16264 5244 16270 5296
rect 16408 5284 16436 5324
rect 16482 5312 16488 5364
rect 16540 5352 16546 5364
rect 16942 5352 16948 5364
rect 16540 5324 16948 5352
rect 16540 5312 16546 5324
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 19334 5352 19340 5364
rect 17052 5324 19340 5352
rect 17052 5284 17080 5324
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 20070 5312 20076 5364
rect 20128 5312 20134 5364
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 21729 5355 21787 5361
rect 21729 5352 21741 5355
rect 21508 5324 21741 5352
rect 21508 5312 21514 5324
rect 21729 5321 21741 5324
rect 21775 5321 21787 5355
rect 27246 5352 27252 5364
rect 21729 5315 21787 5321
rect 26620 5324 27252 5352
rect 16408 5256 17080 5284
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 10091 5120 11560 5148
rect 11624 5120 14228 5148
rect 14292 5188 14657 5216
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 9858 5040 9864 5092
rect 9916 5080 9922 5092
rect 10290 5083 10348 5089
rect 10290 5080 10302 5083
rect 9916 5052 10302 5080
rect 9916 5040 9922 5052
rect 10290 5049 10302 5052
rect 10336 5049 10348 5083
rect 10290 5043 10348 5049
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 11624 5080 11652 5120
rect 10744 5052 11652 5080
rect 12060 5083 12118 5089
rect 10744 5040 10750 5052
rect 12060 5049 12072 5083
rect 12106 5080 12118 5083
rect 13906 5080 13912 5092
rect 12106 5052 13912 5080
rect 12106 5049 12118 5052
rect 12060 5043 12118 5049
rect 13906 5040 13912 5052
rect 13964 5080 13970 5092
rect 14292 5080 14320 5188
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 15010 5176 15016 5228
rect 15068 5176 15074 5228
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 16224 5148 16252 5244
rect 16146 5120 16252 5148
rect 14737 5111 14795 5117
rect 13964 5052 14320 5080
rect 14369 5083 14427 5089
rect 13964 5040 13970 5052
rect 14369 5049 14381 5083
rect 14415 5080 14427 5083
rect 14752 5080 14780 5111
rect 17954 5108 17960 5160
rect 18012 5108 18018 5160
rect 18690 5108 18696 5160
rect 18748 5148 18754 5160
rect 26620 5157 26648 5324
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 27706 5312 27712 5364
rect 27764 5312 27770 5364
rect 27065 5287 27123 5293
rect 27065 5253 27077 5287
rect 27111 5253 27123 5287
rect 27065 5247 27123 5253
rect 27341 5287 27399 5293
rect 27341 5253 27353 5287
rect 27387 5284 27399 5287
rect 27387 5256 27936 5284
rect 27387 5253 27399 5256
rect 27341 5247 27399 5253
rect 27080 5216 27108 5247
rect 27080 5188 27660 5216
rect 27632 5157 27660 5188
rect 27908 5157 27936 5256
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 18748 5120 20361 5148
rect 18748 5108 18754 5120
rect 20349 5117 20361 5120
rect 20395 5117 20407 5151
rect 20605 5151 20663 5157
rect 20605 5148 20617 5151
rect 20349 5111 20407 5117
rect 20548 5120 20617 5148
rect 14415 5052 14596 5080
rect 14752 5052 14872 5080
rect 14415 5049 14427 5052
rect 14369 5043 14427 5049
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 5810 5012 5816 5024
rect 5767 4984 5816 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 5902 4972 5908 5024
rect 5960 4972 5966 5024
rect 7009 5015 7067 5021
rect 7009 4981 7021 5015
rect 7055 5012 7067 5015
rect 7098 5012 7104 5024
rect 7055 4984 7104 5012
rect 7055 4981 7067 4984
rect 7009 4975 7067 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7984 4984 8033 5012
rect 7984 4972 7990 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 8021 4975 8079 4981
rect 8754 4972 8760 5024
rect 8812 4972 8818 5024
rect 9398 4972 9404 5024
rect 9456 5012 9462 5024
rect 9674 5012 9680 5024
rect 9456 4984 9680 5012
rect 9456 4972 9462 4984
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 13262 4972 13268 5024
rect 13320 5012 13326 5024
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 13320 4984 14105 5012
rect 13320 4972 13326 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 14093 4975 14151 4981
rect 14274 4972 14280 5024
rect 14332 4972 14338 5024
rect 14458 4972 14464 5024
rect 14516 4972 14522 5024
rect 14568 5012 14596 5052
rect 14734 5012 14740 5024
rect 14568 4984 14740 5012
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 14844 5012 14872 5052
rect 18414 5040 18420 5092
rect 18472 5080 18478 5092
rect 18938 5083 18996 5089
rect 18938 5080 18950 5083
rect 18472 5052 18950 5080
rect 18472 5040 18478 5052
rect 18938 5049 18950 5052
rect 18984 5049 18996 5083
rect 18938 5043 18996 5049
rect 20548 5024 20576 5120
rect 20605 5117 20617 5120
rect 20651 5117 20663 5151
rect 20605 5111 20663 5117
rect 26605 5151 26663 5157
rect 26605 5117 26617 5151
rect 26651 5117 26663 5151
rect 26881 5151 26939 5157
rect 26881 5148 26893 5151
rect 26605 5111 26663 5117
rect 26804 5120 26893 5148
rect 15654 5012 15660 5024
rect 14844 4984 15660 5012
rect 15654 4972 15660 4984
rect 15712 5012 15718 5024
rect 16574 5012 16580 5024
rect 15712 4984 16580 5012
rect 15712 4972 15718 4984
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 17865 5015 17923 5021
rect 17865 4981 17877 5015
rect 17911 5012 17923 5015
rect 17954 5012 17960 5024
rect 17911 4984 17960 5012
rect 17911 4981 17923 4984
rect 17865 4975 17923 4981
rect 17954 4972 17960 4984
rect 18012 4972 18018 5024
rect 20530 4972 20536 5024
rect 20588 4972 20594 5024
rect 26804 5021 26832 5120
rect 26881 5117 26893 5120
rect 26927 5117 26939 5151
rect 26881 5111 26939 5117
rect 27157 5151 27215 5157
rect 27157 5117 27169 5151
rect 27203 5148 27215 5151
rect 27617 5151 27675 5157
rect 27203 5120 27476 5148
rect 27203 5117 27215 5120
rect 27157 5111 27215 5117
rect 27448 5021 27476 5120
rect 27617 5117 27629 5151
rect 27663 5117 27675 5151
rect 27617 5111 27675 5117
rect 27893 5151 27951 5157
rect 27893 5117 27905 5151
rect 27939 5117 27951 5151
rect 27893 5111 27951 5117
rect 26789 5015 26847 5021
rect 26789 4981 26801 5015
rect 26835 4981 26847 5015
rect 26789 4975 26847 4981
rect 27433 5015 27491 5021
rect 27433 4981 27445 5015
rect 27479 4981 27491 5015
rect 27433 4975 27491 4981
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 3602 4768 3608 4820
rect 3660 4768 3666 4820
rect 4338 4768 4344 4820
rect 4396 4808 4402 4820
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 4396 4780 4445 4808
rect 4396 4768 4402 4780
rect 4433 4777 4445 4780
rect 4479 4777 4491 4811
rect 4433 4771 4491 4777
rect 5350 4768 5356 4820
rect 5408 4768 5414 4820
rect 5902 4768 5908 4820
rect 5960 4768 5966 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 6880 4780 7236 4808
rect 6880 4768 6886 4780
rect 3620 4740 3648 4768
rect 5169 4743 5227 4749
rect 5169 4740 5181 4743
rect 3620 4712 5181 4740
rect 5169 4709 5181 4712
rect 5215 4709 5227 4743
rect 5169 4703 5227 4709
rect 5368 4681 5396 4768
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 5353 4675 5411 4681
rect 5353 4641 5365 4675
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5920 4672 5948 4768
rect 7098 4740 7104 4752
rect 6932 4712 7104 4740
rect 6932 4681 6960 4712
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 7208 4749 7236 4780
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 7340 4780 10241 4808
rect 7340 4768 7346 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 10413 4811 10471 4817
rect 10413 4777 10425 4811
rect 10459 4808 10471 4811
rect 12710 4808 12716 4820
rect 10459 4780 12716 4808
rect 10459 4777 10471 4780
rect 10413 4771 10471 4777
rect 12710 4768 12716 4780
rect 12768 4808 12774 4820
rect 13262 4808 13268 4820
rect 12768 4780 13268 4808
rect 12768 4768 12774 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13722 4808 13728 4820
rect 13587 4780 13728 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14109 4811 14167 4817
rect 14109 4808 14121 4811
rect 13832 4780 14121 4808
rect 7193 4743 7251 4749
rect 7193 4709 7205 4743
rect 7239 4709 7251 4743
rect 7193 4703 7251 4709
rect 7926 4700 7932 4752
rect 7984 4700 7990 4752
rect 8941 4743 8999 4749
rect 8941 4709 8953 4743
rect 8987 4740 8999 4743
rect 10686 4740 10692 4752
rect 8987 4712 10692 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 5583 4644 5948 4672
rect 6917 4675 6975 4681
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 4356 4604 4384 4635
rect 5442 4604 5448 4616
rect 4356 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5644 4468 5672 4567
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 8956 4604 8984 4703
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 13832 4740 13860 4780
rect 14109 4777 14121 4780
rect 14155 4777 14167 4811
rect 14109 4771 14167 4777
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 14550 4808 14556 4820
rect 14415 4780 14556 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 14734 4808 14740 4820
rect 14691 4780 14740 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 14734 4768 14740 4780
rect 14792 4808 14798 4820
rect 18414 4808 18420 4820
rect 14792 4780 18420 4808
rect 14792 4768 14798 4780
rect 12400 4712 13860 4740
rect 12400 4700 12406 4712
rect 9030 4632 9036 4684
rect 9088 4632 9094 4684
rect 9398 4632 9404 4684
rect 9456 4632 9462 4684
rect 9950 4632 9956 4684
rect 10008 4632 10014 4684
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4672 10195 4675
rect 10502 4672 10508 4684
rect 10183 4644 10508 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 11054 4672 11060 4684
rect 10643 4644 11060 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11146 4632 11152 4684
rect 11204 4632 11210 4684
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 12434 4681 12440 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 11572 4644 12173 4672
rect 11572 4632 11578 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 12428 4635 12440 4681
rect 12492 4672 12498 4684
rect 13832 4672 13860 4712
rect 13906 4700 13912 4752
rect 13964 4740 13970 4752
rect 14921 4743 14979 4749
rect 14921 4740 14933 4743
rect 13964 4712 14933 4740
rect 13964 4700 13970 4712
rect 14921 4709 14933 4712
rect 14967 4709 14979 4743
rect 14921 4703 14979 4709
rect 14550 4672 14556 4684
rect 12492 4644 12528 4672
rect 13832 4644 14556 4672
rect 12434 4632 12440 4635
rect 12492 4632 12498 4644
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 15102 4672 15108 4684
rect 14783 4644 15108 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 15580 4681 15608 4780
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20530 4808 20536 4820
rect 20395 4780 20536 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 20530 4768 20536 4780
rect 20588 4808 20594 4820
rect 24857 4811 24915 4817
rect 20588 4780 20760 4808
rect 20588 4768 20594 4780
rect 16945 4743 17003 4749
rect 16945 4740 16957 4743
rect 16500 4712 16957 4740
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 6512 4576 8984 4604
rect 9769 4607 9827 4613
rect 6512 4564 6518 4576
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 9858 4604 9864 4616
rect 9815 4576 9864 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 10704 4576 11376 4604
rect 10704 4536 10732 4576
rect 9048 4508 10732 4536
rect 9048 4468 9076 4508
rect 10778 4496 10784 4548
rect 10836 4496 10842 4548
rect 5644 4440 9076 4468
rect 11238 4428 11244 4480
rect 11296 4428 11302 4480
rect 11348 4468 11376 4576
rect 14292 4576 15485 4604
rect 14292 4545 14320 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 14277 4539 14335 4545
rect 14277 4505 14289 4539
rect 14323 4505 14335 4539
rect 14277 4499 14335 4505
rect 14458 4496 14464 4548
rect 14516 4536 14522 4548
rect 15102 4536 15108 4548
rect 14516 4508 15108 4536
rect 14516 4496 14522 4508
rect 15102 4496 15108 4508
rect 15160 4496 15166 4548
rect 15933 4539 15991 4545
rect 15933 4505 15945 4539
rect 15979 4536 15991 4539
rect 16500 4536 16528 4712
rect 16945 4709 16957 4712
rect 16991 4709 17003 4743
rect 16945 4703 17003 4709
rect 17954 4700 17960 4752
rect 18012 4700 18018 4752
rect 19518 4700 19524 4752
rect 19576 4700 19582 4752
rect 20438 4700 20444 4752
rect 20496 4740 20502 4752
rect 20625 4743 20683 4749
rect 20625 4740 20637 4743
rect 20496 4712 20637 4740
rect 20496 4700 20502 4712
rect 20625 4709 20637 4712
rect 20671 4709 20683 4743
rect 20732 4740 20760 4780
rect 21652 4780 22508 4808
rect 21652 4749 21680 4780
rect 20841 4743 20899 4749
rect 20841 4740 20853 4743
rect 20732 4712 20853 4740
rect 20625 4703 20683 4709
rect 20841 4709 20853 4712
rect 20887 4740 20899 4743
rect 21545 4743 21603 4749
rect 21545 4740 21557 4743
rect 20887 4712 21557 4740
rect 20887 4709 20899 4712
rect 20841 4703 20899 4709
rect 21545 4709 21557 4712
rect 21591 4709 21603 4743
rect 21545 4703 21603 4709
rect 21637 4743 21695 4749
rect 21637 4709 21649 4743
rect 21683 4709 21695 4743
rect 21637 4703 21695 4709
rect 22480 4740 22508 4780
rect 24857 4777 24869 4811
rect 24903 4808 24915 4811
rect 25038 4808 25044 4820
rect 24903 4780 25044 4808
rect 24903 4777 24915 4780
rect 24857 4771 24915 4777
rect 25038 4768 25044 4780
rect 25096 4768 25102 4820
rect 23382 4740 23388 4752
rect 22480 4712 23388 4740
rect 18598 4632 18604 4684
rect 18656 4632 18662 4684
rect 20640 4672 20668 4703
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 20640 4644 21281 4672
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 21450 4632 21456 4684
rect 21508 4632 21514 4684
rect 22480 4681 22508 4712
rect 23382 4700 23388 4712
rect 23440 4740 23446 4752
rect 23722 4743 23780 4749
rect 23722 4740 23734 4743
rect 23440 4712 23734 4740
rect 23440 4700 23446 4712
rect 23722 4709 23734 4712
rect 23768 4709 23780 4743
rect 23722 4703 23780 4709
rect 21821 4675 21879 4681
rect 21821 4641 21833 4675
rect 21867 4672 21879 4675
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21867 4644 22017 4672
rect 21867 4641 21879 4644
rect 21821 4635 21879 4641
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22269 4675 22327 4681
rect 22269 4672 22281 4675
rect 22005 4635 22063 4641
rect 22092 4644 22281 4672
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 16669 4607 16727 4613
rect 16669 4604 16681 4607
rect 16632 4576 16681 4604
rect 16632 4564 16638 4576
rect 16669 4573 16681 4576
rect 16715 4604 16727 4607
rect 18616 4604 18644 4632
rect 16715 4576 18644 4604
rect 18877 4607 18935 4613
rect 16715 4573 16727 4576
rect 16669 4567 16727 4573
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 20806 4604 20812 4616
rect 18923 4576 20812 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 15979 4508 16528 4536
rect 15979 4505 15991 4508
rect 15933 4499 15991 4505
rect 20990 4496 20996 4548
rect 21048 4536 21054 4548
rect 22092 4536 22120 4644
rect 22269 4641 22281 4644
rect 22315 4641 22327 4675
rect 22269 4635 22327 4641
rect 22465 4675 22523 4681
rect 22465 4641 22477 4675
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 22557 4675 22615 4681
rect 22557 4641 22569 4675
rect 22603 4641 22615 4675
rect 22557 4635 22615 4641
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4604 22431 4607
rect 22572 4604 22600 4635
rect 22646 4632 22652 4684
rect 22704 4672 22710 4684
rect 22741 4675 22799 4681
rect 22741 4672 22753 4675
rect 22704 4644 22753 4672
rect 22704 4632 22710 4644
rect 22741 4641 22753 4644
rect 22787 4641 22799 4675
rect 22741 4635 22799 4641
rect 22833 4675 22891 4681
rect 22833 4641 22845 4675
rect 22879 4641 22891 4675
rect 22833 4635 22891 4641
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4672 23535 4675
rect 23566 4672 23572 4684
rect 23523 4644 23572 4672
rect 23523 4641 23535 4644
rect 23477 4635 23535 4641
rect 22419 4576 22600 4604
rect 22419 4573 22431 4576
rect 22373 4567 22431 4573
rect 21048 4508 22120 4536
rect 21048 4496 21054 4508
rect 22186 4496 22192 4548
rect 22244 4536 22250 4548
rect 22848 4536 22876 4635
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 22244 4508 22876 4536
rect 22244 4496 22250 4508
rect 12526 4468 12532 4480
rect 11348 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4468 14151 4471
rect 14476 4468 14504 4496
rect 14139 4440 14504 4468
rect 14139 4437 14151 4440
rect 14093 4431 14151 4437
rect 20622 4428 20628 4480
rect 20680 4468 20686 4480
rect 20809 4471 20867 4477
rect 20809 4468 20821 4471
rect 20680 4440 20821 4468
rect 20680 4428 20686 4440
rect 20809 4437 20821 4440
rect 20855 4468 20867 4471
rect 21450 4468 21456 4480
rect 20855 4440 21456 4468
rect 20855 4437 20867 4440
rect 20809 4431 20867 4437
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 21910 4428 21916 4480
rect 21968 4468 21974 4480
rect 22097 4471 22155 4477
rect 22097 4468 22109 4471
rect 21968 4440 22109 4468
rect 21968 4428 21974 4440
rect 22097 4437 22109 4440
rect 22143 4468 22155 4471
rect 22462 4468 22468 4480
rect 22143 4440 22468 4468
rect 22143 4437 22155 4440
rect 22097 4431 22155 4437
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 22554 4428 22560 4480
rect 22612 4428 22618 4480
rect 22922 4428 22928 4480
rect 22980 4428 22986 4480
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 8205 4267 8263 4273
rect 8205 4233 8217 4267
rect 8251 4264 8263 4267
rect 8754 4264 8760 4276
rect 8251 4236 8760 4264
rect 8251 4233 8263 4236
rect 8205 4227 8263 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 10781 4267 10839 4273
rect 10781 4233 10793 4267
rect 10827 4233 10839 4267
rect 10781 4227 10839 4233
rect 10965 4267 11023 4273
rect 10965 4233 10977 4267
rect 11011 4264 11023 4267
rect 11146 4264 11152 4276
rect 11011 4236 11152 4264
rect 11011 4233 11023 4236
rect 10965 4227 11023 4233
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 8772 4196 8800 4224
rect 10796 4196 10824 4227
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11330 4264 11336 4276
rect 11287 4236 11336 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11054 4196 11060 4208
rect 4120 4168 6500 4196
rect 8772 4168 9996 4196
rect 10796 4168 11060 4196
rect 4120 4156 4126 4168
rect 6472 4137 6500 4168
rect 6457 4131 6515 4137
rect 6457 4097 6469 4131
rect 6503 4128 6515 4131
rect 7098 4128 7104 4140
rect 6503 4100 7104 4128
rect 6503 4097 6515 4100
rect 6457 4091 6515 4097
rect 7098 4088 7104 4100
rect 7156 4128 7162 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 7156 4100 7788 4128
rect 7156 4088 7162 4100
rect 7760 4072 7788 4100
rect 7852 4100 9045 4128
rect 7742 4020 7748 4072
rect 7800 4020 7806 4072
rect 7852 4046 7880 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 9968 4072 9996 4168
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 10778 4128 10784 4140
rect 10428 4100 10784 4128
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 8938 4060 8944 4072
rect 8435 4032 8944 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 9674 4060 9680 4072
rect 9539 4032 9680 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 6733 3995 6791 4001
rect 6733 3961 6745 3995
rect 6779 3992 6791 3995
rect 8665 3995 8723 4001
rect 6779 3964 7144 3992
rect 6779 3961 6791 3964
rect 6733 3955 6791 3961
rect 7116 3924 7144 3964
rect 8036 3964 8340 3992
rect 8036 3924 8064 3964
rect 7116 3896 8064 3924
rect 8312 3924 8340 3964
rect 8665 3961 8677 3995
rect 8711 3992 8723 3995
rect 9030 3992 9036 4004
rect 8711 3964 9036 3992
rect 8711 3961 8723 3964
rect 8665 3955 8723 3961
rect 9030 3952 9036 3964
rect 9088 3992 9094 4004
rect 9140 3992 9168 4023
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 9088 3964 9168 3992
rect 9088 3952 9094 3964
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 8312 3896 9321 3924
rect 9309 3893 9321 3896
rect 9355 3893 9367 3927
rect 9784 3924 9812 4023
rect 9950 4020 9956 4072
rect 10008 4020 10014 4072
rect 10428 3992 10456 4100
rect 10778 4088 10784 4100
rect 10836 4128 10842 4140
rect 11256 4128 11284 4227
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 12621 4267 12679 4273
rect 12621 4264 12633 4267
rect 12584 4236 12633 4264
rect 12584 4224 12590 4236
rect 12621 4233 12633 4236
rect 12667 4264 12679 4267
rect 14090 4264 14096 4276
rect 12667 4236 14096 4264
rect 12667 4233 12679 4236
rect 12621 4227 12679 4233
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 14550 4224 14556 4276
rect 14608 4224 14614 4276
rect 15166 4236 18276 4264
rect 11606 4128 11612 4140
rect 10836 4100 11284 4128
rect 11348 4100 11612 4128
rect 10836 4088 10842 4100
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 10560 4032 10732 4060
rect 10560 4020 10566 4032
rect 10597 3995 10655 4001
rect 10597 3992 10609 3995
rect 10428 3964 10609 3992
rect 10597 3961 10609 3964
rect 10643 3961 10655 3995
rect 10704 3992 10732 4032
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11348 4060 11376 4100
rect 11606 4088 11612 4100
rect 11664 4128 11670 4140
rect 11664 4100 12572 4128
rect 11664 4088 11670 4100
rect 12360 4072 12388 4100
rect 11296 4032 11376 4060
rect 12253 4063 12311 4069
rect 11296 4020 11302 4032
rect 12253 4029 12265 4063
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 10797 3995 10855 4001
rect 10797 3992 10809 3995
rect 10704 3964 10809 3992
rect 10597 3955 10655 3961
rect 10797 3961 10809 3964
rect 10843 3961 10855 3995
rect 10797 3955 10855 3961
rect 11330 3952 11336 4004
rect 11388 3992 11394 4004
rect 11425 3995 11483 4001
rect 11425 3992 11437 3995
rect 11388 3964 11437 3992
rect 11388 3952 11394 3964
rect 11425 3961 11437 3964
rect 11471 3961 11483 3995
rect 12268 3992 12296 4023
rect 12342 4020 12348 4072
rect 12400 4020 12406 4072
rect 12434 4020 12440 4072
rect 12492 4020 12498 4072
rect 12544 4069 12572 4100
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4029 12587 4063
rect 12529 4023 12587 4029
rect 12710 4020 12716 4072
rect 12768 4020 12774 4072
rect 14568 3992 14596 4224
rect 15166 4208 15194 4236
rect 18248 4208 18276 4236
rect 19518 4224 19524 4276
rect 19576 4264 19582 4276
rect 19613 4267 19671 4273
rect 19613 4264 19625 4267
rect 19576 4236 19625 4264
rect 19576 4224 19582 4236
rect 19613 4233 19625 4236
rect 19659 4233 19671 4267
rect 19613 4227 19671 4233
rect 19700 4236 20484 4264
rect 15102 4156 15108 4208
rect 15160 4168 15194 4208
rect 15657 4199 15715 4205
rect 15657 4196 15669 4199
rect 15396 4168 15669 4196
rect 15160 4156 15166 4168
rect 15120 4069 15148 4156
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 15396 4128 15424 4168
rect 15657 4165 15669 4168
rect 15703 4165 15715 4199
rect 15657 4159 15715 4165
rect 16224 4168 16620 4196
rect 15243 4100 15424 4128
rect 15488 4100 15792 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4029 15163 4063
rect 15488 4060 15516 4100
rect 15105 4023 15163 4029
rect 15212 4032 15516 4060
rect 15212 3992 15240 4032
rect 15562 4020 15568 4072
rect 15620 4020 15626 4072
rect 15764 4069 15792 4100
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 16224 4128 16252 4168
rect 15896 4100 16252 4128
rect 16592 4128 16620 4168
rect 18230 4156 18236 4208
rect 18288 4156 18294 4208
rect 18598 4156 18604 4208
rect 18656 4196 18662 4208
rect 19700 4196 19728 4236
rect 18656 4168 19728 4196
rect 20349 4199 20407 4205
rect 18656 4156 18662 4168
rect 20349 4165 20361 4199
rect 20395 4165 20407 4199
rect 20456 4196 20484 4236
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 20901 4227 20959 4233
rect 23382 4224 23388 4276
rect 23440 4264 23446 4276
rect 23661 4267 23719 4273
rect 23661 4264 23673 4267
rect 23440 4236 23673 4264
rect 23440 4224 23446 4236
rect 23661 4233 23673 4236
rect 23707 4233 23719 4267
rect 23661 4227 23719 4233
rect 20456 4168 21956 4196
rect 20349 4159 20407 4165
rect 20364 4128 20392 4159
rect 21928 4137 21956 4168
rect 21913 4131 21971 4137
rect 16592 4100 18920 4128
rect 20364 4100 20760 4128
rect 15896 4088 15902 4100
rect 15749 4063 15807 4069
rect 15749 4029 15761 4063
rect 15795 4029 15807 4063
rect 15749 4023 15807 4029
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 16482 4060 16488 4072
rect 16264 4032 16488 4060
rect 16264 4020 16270 4032
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 18892 4069 18920 4100
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4060 18935 4063
rect 19334 4060 19340 4072
rect 18923 4032 19340 4060
rect 18923 4029 18935 4032
rect 18877 4023 18935 4029
rect 19334 4020 19340 4032
rect 19392 4060 19398 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19392 4032 19533 4060
rect 19392 4020 19398 4032
rect 19521 4029 19533 4032
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 20349 4063 20407 4069
rect 20349 4029 20361 4063
rect 20395 4060 20407 4063
rect 20530 4060 20536 4072
rect 20395 4032 20536 4060
rect 20395 4029 20407 4032
rect 20349 4023 20407 4029
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20622 4020 20628 4072
rect 20680 4020 20686 4072
rect 20732 4069 20760 4100
rect 21913 4097 21925 4131
rect 21959 4097 21971 4131
rect 21913 4091 21971 4097
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4128 22247 4131
rect 22554 4128 22560 4140
rect 22235 4100 22560 4128
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22554 4088 22560 4100
rect 22612 4088 22618 4140
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 24857 4131 24915 4137
rect 24857 4128 24869 4131
rect 23624 4100 24869 4128
rect 23624 4088 23630 4100
rect 24857 4097 24869 4100
rect 24903 4097 24915 4131
rect 24857 4091 24915 4097
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 20901 4063 20959 4069
rect 20901 4029 20913 4063
rect 20947 4060 20959 4063
rect 20990 4060 20996 4072
rect 20947 4032 20996 4060
rect 20947 4029 20959 4032
rect 20901 4023 20959 4029
rect 20990 4020 20996 4032
rect 21048 4020 21054 4072
rect 16761 3995 16819 4001
rect 16761 3992 16773 3995
rect 12268 3964 12572 3992
rect 14568 3964 15240 3992
rect 15488 3964 16773 3992
rect 11425 3955 11483 3961
rect 12544 3936 12572 3964
rect 11054 3924 11060 3936
rect 9784 3896 11060 3924
rect 9309 3887 9367 3893
rect 11054 3884 11060 3896
rect 11112 3924 11118 3936
rect 11238 3933 11244 3936
rect 11225 3927 11244 3933
rect 11112 3896 11157 3924
rect 11112 3884 11118 3896
rect 11225 3893 11237 3927
rect 11296 3924 11302 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11296 3896 12081 3924
rect 11225 3887 11244 3893
rect 11238 3884 11244 3887
rect 11296 3884 11302 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 12526 3884 12532 3936
rect 12584 3884 12590 3936
rect 15488 3933 15516 3964
rect 16761 3961 16773 3964
rect 16807 3961 16819 3995
rect 18785 3995 18843 4001
rect 18785 3992 18797 3995
rect 17986 3964 18797 3992
rect 16761 3955 16819 3961
rect 18785 3961 18797 3964
rect 18831 3961 18843 3995
rect 22094 3992 22100 4004
rect 18785 3955 18843 3961
rect 18892 3964 22100 3992
rect 15473 3927 15531 3933
rect 15473 3893 15485 3927
rect 15519 3893 15531 3927
rect 15473 3887 15531 3893
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 18892 3924 18920 3964
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 22922 3952 22928 4004
rect 22980 3952 22986 4004
rect 23842 3952 23848 4004
rect 23900 3992 23906 4004
rect 25102 3995 25160 4001
rect 25102 3992 25114 3995
rect 23900 3964 25114 3992
rect 23900 3952 23906 3964
rect 25102 3961 25114 3964
rect 25148 3961 25160 3995
rect 25102 3955 25160 3961
rect 18288 3896 18920 3924
rect 18288 3884 18294 3896
rect 18966 3884 18972 3936
rect 19024 3924 19030 3936
rect 20438 3924 20444 3936
rect 19024 3896 20444 3924
rect 19024 3884 19030 3896
rect 20438 3884 20444 3896
rect 20496 3924 20502 3936
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 20496 3896 20545 3924
rect 20496 3884 20502 3896
rect 20533 3893 20545 3896
rect 20579 3924 20591 3927
rect 21082 3924 21088 3936
rect 20579 3896 21088 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 26234 3884 26240 3936
rect 26292 3884 26298 3936
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 11606 3720 11612 3732
rect 9732 3692 11612 3720
rect 9732 3680 9738 3692
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11977 3723 12035 3729
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 12434 3720 12440 3732
rect 12023 3692 12440 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12434 3680 12440 3692
rect 12492 3720 12498 3732
rect 13722 3720 13728 3732
rect 12492 3692 13728 3720
rect 12492 3680 12498 3692
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 13924 3692 15117 3720
rect 13924 3664 13952 3692
rect 15105 3689 15117 3692
rect 15151 3720 15163 3723
rect 15562 3720 15568 3732
rect 15151 3692 15568 3720
rect 15151 3689 15163 3692
rect 15105 3683 15163 3689
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 21450 3680 21456 3732
rect 21508 3720 21514 3732
rect 23293 3723 23351 3729
rect 23293 3720 23305 3723
rect 21508 3692 23305 3720
rect 21508 3680 21514 3692
rect 23293 3689 23305 3692
rect 23339 3720 23351 3723
rect 23934 3720 23940 3732
rect 23339 3692 23940 3720
rect 23339 3689 23351 3692
rect 23293 3683 23351 3689
rect 23934 3680 23940 3692
rect 23992 3680 23998 3732
rect 9122 3612 9128 3664
rect 9180 3612 9186 3664
rect 10965 3655 11023 3661
rect 10965 3652 10977 3655
rect 10336 3624 10977 3652
rect 7742 3544 7748 3596
rect 7800 3584 7806 3596
rect 8110 3584 8116 3596
rect 7800 3556 8116 3584
rect 7800 3544 7806 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 10134 3544 10140 3596
rect 10192 3544 10198 3596
rect 10336 3593 10364 3624
rect 10965 3621 10977 3624
rect 11011 3652 11023 3655
rect 11011 3624 11468 3652
rect 11011 3621 11023 3624
rect 10965 3615 11023 3621
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3584 10655 3587
rect 11054 3584 11060 3596
rect 10643 3556 11060 3584
rect 10643 3553 10655 3556
rect 10597 3547 10655 3553
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 10229 3519 10287 3525
rect 8435 3488 9444 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 9416 3448 9444 3488
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10428 3516 10456 3547
rect 11054 3544 11060 3556
rect 11112 3544 11118 3596
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11238 3584 11244 3596
rect 11195 3556 11244 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11440 3593 11468 3624
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 12250 3652 12256 3664
rect 11572 3624 12256 3652
rect 11572 3612 11578 3624
rect 11425 3587 11483 3593
rect 11425 3553 11437 3587
rect 11471 3553 11483 3587
rect 11425 3547 11483 3553
rect 10275 3488 10456 3516
rect 11333 3519 11391 3525
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11532 3516 11560 3612
rect 11900 3593 11928 3624
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 13906 3652 13912 3664
rect 12912 3624 13912 3652
rect 11609 3587 11667 3593
rect 11609 3553 11621 3587
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 11885 3587 11943 3593
rect 11885 3553 11897 3587
rect 11931 3553 11943 3587
rect 11885 3547 11943 3553
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3584 12219 3587
rect 12526 3584 12532 3596
rect 12207 3556 12532 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 11379 3488 11560 3516
rect 11624 3516 11652 3547
rect 12526 3544 12532 3556
rect 12584 3584 12590 3596
rect 12710 3584 12716 3596
rect 12584 3556 12716 3584
rect 12584 3544 12590 3556
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 12912 3593 12940 3624
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 15381 3655 15439 3661
rect 15381 3652 15393 3655
rect 14858 3624 15393 3652
rect 15381 3621 15393 3624
rect 15427 3621 15439 3655
rect 15381 3615 15439 3621
rect 16758 3612 16764 3664
rect 16816 3652 16822 3664
rect 18877 3655 18935 3661
rect 16816 3624 18828 3652
rect 16816 3612 16822 3624
rect 12897 3587 12955 3593
rect 12897 3553 12909 3587
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 14976 3556 15485 3584
rect 14976 3544 14982 3556
rect 15473 3553 15485 3556
rect 15519 3584 15531 3587
rect 15654 3584 15660 3596
rect 15519 3556 15660 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 16301 3587 16359 3593
rect 16301 3553 16313 3587
rect 16347 3584 16359 3587
rect 18414 3584 18420 3596
rect 16347 3556 18420 3584
rect 16347 3553 16359 3556
rect 16301 3547 16359 3553
rect 11624 3488 12204 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 12176 3457 12204 3488
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 12400 3488 12817 3516
rect 12400 3476 12406 3488
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 12805 3479 12863 3485
rect 13188 3488 13369 3516
rect 10413 3451 10471 3457
rect 10413 3448 10425 3451
rect 9416 3420 10425 3448
rect 10413 3417 10425 3420
rect 10459 3417 10471 3451
rect 10413 3411 10471 3417
rect 12161 3451 12219 3457
rect 12161 3417 12173 3451
rect 12207 3417 12219 3451
rect 12161 3411 12219 3417
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10134 3380 10140 3392
rect 9916 3352 10140 3380
rect 9916 3340 9922 3352
rect 10134 3340 10140 3352
rect 10192 3380 10198 3392
rect 11330 3380 11336 3392
rect 10192 3352 11336 3380
rect 10192 3340 10198 3352
rect 11330 3340 11336 3352
rect 11388 3340 11394 3392
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 13188 3380 13216 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13357 3479 13415 3485
rect 13464 3488 13645 3516
rect 13265 3451 13323 3457
rect 13265 3417 13277 3451
rect 13311 3448 13323 3451
rect 13464 3448 13492 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 16316 3516 16344 3547
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 18800 3593 18828 3624
rect 18877 3621 18889 3655
rect 18923 3652 18935 3655
rect 19337 3655 19395 3661
rect 19337 3652 19349 3655
rect 18923 3624 19349 3652
rect 18923 3621 18935 3624
rect 18877 3615 18935 3621
rect 19337 3621 19349 3624
rect 19383 3621 19395 3655
rect 19337 3615 19395 3621
rect 20070 3612 20076 3664
rect 20128 3612 20134 3664
rect 21082 3612 21088 3664
rect 21140 3612 21146 3664
rect 23569 3655 23627 3661
rect 23569 3652 23581 3655
rect 23046 3624 23581 3652
rect 23569 3621 23581 3624
rect 23615 3621 23627 3655
rect 23569 3615 23627 3621
rect 18785 3587 18843 3593
rect 18785 3553 18797 3587
rect 18831 3584 18843 3587
rect 18966 3584 18972 3596
rect 18831 3556 18972 3584
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 21545 3587 21603 3593
rect 21545 3584 21557 3587
rect 20548 3556 21557 3584
rect 13780 3488 16344 3516
rect 16393 3519 16451 3525
rect 13780 3476 13786 3488
rect 16393 3485 16405 3519
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 13311 3420 13492 3448
rect 13311 3417 13323 3420
rect 13265 3411 13323 3417
rect 14642 3408 14648 3460
rect 14700 3448 14706 3460
rect 16408 3448 16436 3479
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 19061 3519 19119 3525
rect 19061 3516 19073 3519
rect 16540 3488 19073 3516
rect 16540 3476 16546 3488
rect 19061 3485 19073 3488
rect 19107 3516 19119 3519
rect 20548 3516 20576 3556
rect 21545 3553 21557 3556
rect 21591 3553 21603 3587
rect 21545 3547 21603 3553
rect 23477 3587 23535 3593
rect 23477 3553 23489 3587
rect 23523 3553 23535 3587
rect 23477 3547 23535 3553
rect 19107 3488 20576 3516
rect 19107 3485 19119 3488
rect 19061 3479 19119 3485
rect 21818 3476 21824 3528
rect 21876 3476 21882 3528
rect 22186 3476 22192 3528
rect 22244 3516 22250 3528
rect 23492 3516 23520 3547
rect 22244 3488 23520 3516
rect 22244 3476 22250 3488
rect 14700 3420 19196 3448
rect 14700 3408 14706 3420
rect 16206 3380 16212 3392
rect 13188 3352 16212 3380
rect 16206 3340 16212 3352
rect 16264 3340 16270 3392
rect 16669 3383 16727 3389
rect 16669 3349 16681 3383
rect 16715 3380 16727 3383
rect 16942 3380 16948 3392
rect 16715 3352 16948 3380
rect 16715 3349 16727 3352
rect 16669 3343 16727 3349
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 19168 3380 19196 3420
rect 21910 3380 21916 3392
rect 19168 3352 21916 3380
rect 21910 3340 21916 3352
rect 21968 3340 21974 3392
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 9122 3136 9128 3188
rect 9180 3136 9186 3188
rect 10980 3148 12664 3176
rect 8110 3068 8116 3120
rect 8168 3108 8174 3120
rect 10980 3108 11008 3148
rect 8168 3080 11008 3108
rect 12636 3108 12664 3148
rect 12710 3136 12716 3188
rect 12768 3136 12774 3188
rect 16482 3136 16488 3188
rect 16540 3136 16546 3188
rect 20070 3136 20076 3188
rect 20128 3176 20134 3188
rect 20165 3179 20223 3185
rect 20165 3176 20177 3179
rect 20128 3148 20177 3176
rect 20128 3136 20134 3148
rect 20165 3145 20177 3148
rect 20211 3145 20223 3179
rect 20165 3139 20223 3145
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 21818 3176 21824 3188
rect 21315 3148 21824 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 23842 3136 23848 3188
rect 23900 3136 23906 3188
rect 16500 3108 16528 3136
rect 12636 3080 16528 3108
rect 8168 3068 8174 3080
rect 10980 3049 11008 3080
rect 18414 3068 18420 3120
rect 18472 3108 18478 3120
rect 23860 3108 23888 3136
rect 18472 3080 23888 3108
rect 18472 3068 18478 3080
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11241 3043 11299 3049
rect 11241 3009 11253 3043
rect 11287 3040 11299 3043
rect 11606 3040 11612 3052
rect 11287 3012 11612 3040
rect 11287 3009 11299 3012
rect 11241 3003 11299 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 16206 3000 16212 3052
rect 16264 3040 16270 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16264 3012 16681 3040
rect 16264 3000 16270 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 20993 3043 21051 3049
rect 20993 3009 21005 3043
rect 21039 3040 21051 3043
rect 21450 3040 21456 3052
rect 21039 3012 21456 3040
rect 21039 3009 21051 3012
rect 20993 3003 21051 3009
rect 21450 3000 21456 3012
rect 21508 3000 21514 3052
rect 9030 2932 9036 2984
rect 9088 2932 9094 2984
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 14918 2972 14924 2984
rect 13035 2944 14924 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 9048 2836 9076 2932
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 12466 2876 12909 2904
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 13004 2836 13032 2935
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2972 18935 2975
rect 19334 2972 19340 2984
rect 18923 2944 19340 2972
rect 18923 2941 18935 2944
rect 18877 2935 18935 2941
rect 19334 2932 19340 2944
rect 19392 2972 19398 2984
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19392 2944 20085 2972
rect 19392 2932 19398 2944
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 20901 2975 20959 2981
rect 20901 2941 20913 2975
rect 20947 2972 20959 2975
rect 21082 2972 21088 2984
rect 20947 2944 21088 2972
rect 20947 2941 20959 2944
rect 20901 2935 20959 2941
rect 16942 2864 16948 2916
rect 17000 2864 17006 2916
rect 18785 2907 18843 2913
rect 18785 2904 18797 2907
rect 18170 2876 18797 2904
rect 18785 2873 18797 2876
rect 18831 2873 18843 2907
rect 20088 2904 20116 2935
rect 21082 2932 21088 2944
rect 21140 2932 21146 2984
rect 22186 2904 22192 2916
rect 20088 2876 22192 2904
rect 18785 2867 18843 2873
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 9048 2808 13032 2836
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 15749 1003 15807 1009
rect 15749 969 15761 1003
rect 15795 1000 15807 1003
rect 16298 1000 16304 1012
rect 15795 972 16304 1000
rect 15795 969 15807 972
rect 15749 963 15807 969
rect 16298 960 16304 972
rect 16356 960 16362 1012
rect 16390 960 16396 1012
rect 16448 960 16454 1012
rect 16850 960 16856 1012
rect 16908 960 16914 1012
rect 6546 756 6552 808
rect 6604 756 6610 808
rect 14274 756 14280 808
rect 14332 756 14338 808
rect 15562 756 15568 808
rect 15620 756 15626 808
rect 16206 756 16212 808
rect 16264 756 16270 808
rect 16758 756 16764 808
rect 16816 796 16822 808
rect 17037 799 17095 805
rect 17037 796 17049 799
rect 16816 768 17049 796
rect 16816 756 16822 768
rect 17037 765 17049 768
rect 17083 765 17095 799
rect 17037 759 17095 765
rect 18782 756 18788 808
rect 18840 756 18846 808
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 10324 18776 10376 18828
rect 10968 18776 11020 18828
rect 12256 18776 12308 18828
rect 12900 18776 12952 18828
rect 16212 18819 16264 18828
rect 16212 18785 16221 18819
rect 16221 18785 16255 18819
rect 16255 18785 16264 18819
rect 16212 18776 16264 18785
rect 18052 18776 18104 18828
rect 18696 18776 18748 18828
rect 19340 18776 19392 18828
rect 19984 18776 20036 18828
rect 20628 18776 20680 18828
rect 21272 18776 21324 18828
rect 21916 18776 21968 18828
rect 31024 18615 31076 18624
rect 31024 18581 31033 18615
rect 31033 18581 31067 18615
rect 31067 18581 31076 18615
rect 31024 18572 31076 18581
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 18236 16779 18288 16788
rect 18236 16745 18245 16779
rect 18245 16745 18279 16779
rect 18279 16745 18288 16779
rect 18236 16736 18288 16745
rect 8944 16600 8996 16652
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 10324 16600 10376 16652
rect 11520 16668 11572 16720
rect 12624 16668 12676 16720
rect 15108 16600 15160 16652
rect 11612 16575 11664 16584
rect 11612 16541 11621 16575
rect 11621 16541 11655 16575
rect 11655 16541 11664 16575
rect 11612 16532 11664 16541
rect 19156 16532 19208 16584
rect 22468 16532 22520 16584
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 9772 16439 9824 16448
rect 9772 16405 9781 16439
rect 9781 16405 9815 16439
rect 9815 16405 9824 16439
rect 9772 16396 9824 16405
rect 11428 16396 11480 16448
rect 21548 16439 21600 16448
rect 21548 16405 21557 16439
rect 21557 16405 21591 16439
rect 21591 16405 21600 16439
rect 21548 16396 21600 16405
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 6644 16192 6696 16244
rect 10324 16192 10376 16244
rect 11612 16192 11664 16244
rect 12624 16192 12676 16244
rect 15384 16235 15436 16244
rect 9772 16056 9824 16108
rect 11520 16124 11572 16176
rect 10876 16056 10928 16108
rect 12716 16056 12768 16108
rect 9128 15920 9180 15972
rect 9036 15852 9088 15904
rect 10416 16031 10468 16040
rect 10416 15997 10425 16031
rect 10425 15997 10459 16031
rect 10459 15997 10468 16031
rect 10416 15988 10468 15997
rect 11428 15988 11480 16040
rect 12808 15988 12860 16040
rect 11060 15920 11112 15972
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 15016 16124 15068 16176
rect 15660 16056 15712 16108
rect 17224 16056 17276 16108
rect 18236 16056 18288 16108
rect 21456 16056 21508 16108
rect 22468 16056 22520 16108
rect 13544 15920 13596 15972
rect 14648 15920 14700 15972
rect 14924 15852 14976 15904
rect 17960 15988 18012 16040
rect 18328 15852 18380 15904
rect 18972 15963 19024 15972
rect 18972 15929 18981 15963
rect 18981 15929 19015 15963
rect 19015 15929 19024 15963
rect 18972 15920 19024 15929
rect 19432 15920 19484 15972
rect 20904 15963 20956 15972
rect 20904 15929 20913 15963
rect 20913 15929 20947 15963
rect 20947 15929 20956 15963
rect 20904 15920 20956 15929
rect 21548 15920 21600 15972
rect 19156 15852 19208 15904
rect 20260 15852 20312 15904
rect 20536 15852 20588 15904
rect 22836 15895 22888 15904
rect 22836 15861 22845 15895
rect 22845 15861 22879 15895
rect 22879 15861 22888 15895
rect 22836 15852 22888 15861
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 7932 15580 7984 15632
rect 6092 15444 6144 15496
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 9036 15648 9088 15700
rect 10416 15648 10468 15700
rect 9128 15555 9180 15564
rect 9128 15521 9137 15555
rect 9137 15521 9171 15555
rect 9171 15521 9180 15555
rect 9128 15512 9180 15521
rect 11428 15691 11480 15700
rect 11428 15657 11437 15691
rect 11437 15657 11471 15691
rect 11471 15657 11480 15691
rect 11428 15648 11480 15657
rect 11704 15648 11756 15700
rect 12624 15648 12676 15700
rect 12716 15648 12768 15700
rect 14648 15648 14700 15700
rect 15660 15648 15712 15700
rect 18972 15648 19024 15700
rect 19432 15648 19484 15700
rect 10508 15555 10560 15564
rect 10508 15521 10517 15555
rect 10517 15521 10551 15555
rect 10551 15521 10560 15555
rect 10508 15512 10560 15521
rect 10876 15512 10928 15564
rect 11612 15555 11664 15564
rect 11612 15521 11621 15555
rect 11621 15521 11655 15555
rect 11655 15521 11664 15555
rect 11612 15512 11664 15521
rect 9588 15444 9640 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 11060 15444 11112 15496
rect 12808 15376 12860 15428
rect 13728 15376 13780 15428
rect 15384 15580 15436 15632
rect 15660 15555 15712 15564
rect 15660 15521 15669 15555
rect 15669 15521 15703 15555
rect 15703 15521 15712 15555
rect 15660 15512 15712 15521
rect 17960 15376 18012 15428
rect 19156 15512 19208 15564
rect 20076 15512 20128 15564
rect 20260 15512 20312 15564
rect 20628 15555 20680 15564
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 20812 15555 20864 15564
rect 20812 15521 20821 15555
rect 20821 15521 20855 15555
rect 20855 15521 20864 15555
rect 20812 15512 20864 15521
rect 20996 15555 21048 15564
rect 20996 15521 21005 15555
rect 21005 15521 21039 15555
rect 21039 15521 21048 15555
rect 20996 15512 21048 15521
rect 22836 15580 22888 15632
rect 20536 15444 20588 15496
rect 20904 15444 20956 15496
rect 23664 15555 23716 15564
rect 23664 15521 23673 15555
rect 23673 15521 23707 15555
rect 23707 15521 23716 15555
rect 23664 15512 23716 15521
rect 21456 15376 21508 15428
rect 23296 15376 23348 15428
rect 9588 15308 9640 15360
rect 10324 15308 10376 15360
rect 11796 15308 11848 15360
rect 18144 15308 18196 15360
rect 20352 15308 20404 15360
rect 20812 15308 20864 15360
rect 24124 15308 24176 15360
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 3240 14900 3292 14952
rect 6092 14968 6144 15020
rect 9128 15036 9180 15088
rect 9036 14968 9088 15020
rect 10508 15104 10560 15156
rect 10140 15036 10192 15088
rect 14924 15011 14976 15020
rect 6276 14943 6328 14952
rect 6276 14909 6285 14943
rect 6285 14909 6319 14943
rect 6319 14909 6328 14943
rect 6276 14900 6328 14909
rect 6460 14943 6512 14952
rect 6460 14909 6469 14943
rect 6469 14909 6503 14943
rect 6503 14909 6512 14943
rect 6460 14900 6512 14909
rect 8944 14900 8996 14952
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 10508 14900 10560 14952
rect 11060 14900 11112 14952
rect 4068 14875 4120 14884
rect 4068 14841 4077 14875
rect 4077 14841 4111 14875
rect 4111 14841 4120 14875
rect 4068 14832 4120 14841
rect 4804 14832 4856 14884
rect 4712 14764 4764 14816
rect 6368 14764 6420 14816
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 7012 14764 7064 14816
rect 9956 14764 10008 14816
rect 10324 14832 10376 14884
rect 11428 14943 11480 14952
rect 11428 14909 11437 14943
rect 11437 14909 11471 14943
rect 11471 14909 11480 14943
rect 11428 14900 11480 14909
rect 11520 14900 11572 14952
rect 13728 14943 13780 14952
rect 13728 14909 13737 14943
rect 13737 14909 13771 14943
rect 13771 14909 13780 14943
rect 13728 14900 13780 14909
rect 15936 15104 15988 15156
rect 15384 15036 15436 15088
rect 16304 14968 16356 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 20444 15104 20496 15156
rect 20536 15104 20588 15156
rect 20628 15147 20680 15156
rect 20628 15113 20637 15147
rect 20637 15113 20671 15147
rect 20671 15113 20680 15147
rect 20628 15104 20680 15113
rect 11796 14832 11848 14884
rect 11612 14764 11664 14816
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 13544 14764 13596 14816
rect 16212 14900 16264 14952
rect 16764 14943 16816 14952
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 17500 14900 17552 14952
rect 18144 14900 18196 14952
rect 15200 14832 15252 14884
rect 15660 14832 15712 14884
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 15936 14807 15988 14816
rect 15936 14773 15945 14807
rect 15945 14773 15979 14807
rect 15979 14773 15988 14807
rect 15936 14764 15988 14773
rect 16580 14764 16632 14816
rect 17592 14764 17644 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 18788 14900 18840 14952
rect 19156 14832 19208 14884
rect 19892 14900 19944 14952
rect 20076 15079 20128 15088
rect 20076 15045 20085 15079
rect 20085 15045 20119 15079
rect 20119 15045 20128 15079
rect 20076 15036 20128 15045
rect 20260 15036 20312 15088
rect 20996 15104 21048 15156
rect 21456 14968 21508 15020
rect 23940 14900 23992 14952
rect 24124 14943 24176 14952
rect 24124 14909 24158 14943
rect 24158 14909 24176 14943
rect 24124 14900 24176 14909
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 20260 14807 20312 14816
rect 20260 14773 20269 14807
rect 20269 14773 20303 14807
rect 20303 14773 20312 14807
rect 20260 14764 20312 14773
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 20720 14875 20772 14884
rect 20720 14841 20729 14875
rect 20729 14841 20763 14875
rect 20763 14841 20772 14875
rect 20720 14832 20772 14841
rect 22652 14832 22704 14884
rect 23848 14764 23900 14816
rect 25044 14764 25096 14816
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 4804 14560 4856 14612
rect 6276 14560 6328 14612
rect 6368 14560 6420 14612
rect 848 14467 900 14476
rect 848 14433 857 14467
rect 857 14433 891 14467
rect 891 14433 900 14467
rect 848 14424 900 14433
rect 3424 14492 3476 14544
rect 6644 14560 6696 14612
rect 6736 14560 6788 14612
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 3700 14399 3752 14408
rect 3700 14365 3709 14399
rect 3709 14365 3743 14399
rect 3743 14365 3752 14399
rect 3700 14356 3752 14365
rect 2412 14288 2464 14340
rect 4068 14424 4120 14476
rect 4896 14424 4948 14476
rect 4712 14288 4764 14340
rect 4804 14220 4856 14272
rect 7564 14492 7616 14544
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 8944 14560 8996 14612
rect 9128 14492 9180 14544
rect 6644 14356 6696 14408
rect 6920 14356 6972 14408
rect 11428 14560 11480 14612
rect 13360 14560 13412 14612
rect 15016 14603 15068 14612
rect 15016 14569 15025 14603
rect 15025 14569 15059 14603
rect 15059 14569 15068 14603
rect 15016 14560 15068 14569
rect 16120 14560 16172 14612
rect 16212 14560 16264 14612
rect 17132 14560 17184 14612
rect 12808 14424 12860 14476
rect 14924 14424 14976 14476
rect 15108 14467 15160 14476
rect 15108 14433 15117 14467
rect 15117 14433 15151 14467
rect 15151 14433 15160 14467
rect 15108 14424 15160 14433
rect 15568 14492 15620 14544
rect 16764 14492 16816 14544
rect 11244 14356 11296 14408
rect 13268 14399 13320 14408
rect 7656 14220 7708 14272
rect 9772 14220 9824 14272
rect 9864 14220 9916 14272
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 16212 14424 16264 14476
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 15200 14288 15252 14340
rect 17224 14424 17276 14476
rect 17592 14492 17644 14544
rect 22652 14603 22704 14612
rect 22652 14569 22661 14603
rect 22661 14569 22695 14603
rect 22695 14569 22704 14603
rect 22652 14560 22704 14569
rect 18420 14492 18472 14544
rect 22468 14424 22520 14476
rect 23204 14424 23256 14476
rect 23296 14467 23348 14476
rect 23296 14433 23305 14467
rect 23305 14433 23339 14467
rect 23339 14433 23348 14467
rect 23296 14424 23348 14433
rect 23848 14492 23900 14544
rect 23940 14424 23992 14476
rect 14832 14220 14884 14272
rect 15108 14220 15160 14272
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 18696 14220 18748 14272
rect 23204 14220 23256 14272
rect 25504 14220 25556 14272
rect 26240 14263 26292 14272
rect 26240 14229 26249 14263
rect 26249 14229 26283 14263
rect 26283 14229 26292 14263
rect 26240 14220 26292 14229
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 2412 13948 2464 14000
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 3700 14016 3752 14068
rect 4344 14016 4396 14068
rect 7012 14016 7064 14068
rect 7564 14016 7616 14068
rect 13268 14016 13320 14068
rect 13912 14016 13964 14068
rect 4712 13991 4764 14000
rect 4712 13957 4721 13991
rect 4721 13957 4755 13991
rect 4755 13957 4764 13991
rect 4712 13948 4764 13957
rect 8024 13948 8076 14000
rect 4344 13787 4396 13796
rect 4344 13753 4353 13787
rect 4353 13753 4387 13787
rect 4387 13753 4396 13787
rect 4344 13744 4396 13753
rect 4804 13812 4856 13864
rect 4988 13855 5040 13864
rect 4988 13821 4997 13855
rect 4997 13821 5031 13855
rect 5031 13821 5040 13855
rect 4988 13812 5040 13821
rect 6460 13923 6512 13932
rect 6460 13889 6469 13923
rect 6469 13889 6503 13923
rect 6503 13889 6512 13923
rect 6460 13880 6512 13889
rect 7012 13812 7064 13864
rect 7104 13812 7156 13864
rect 7656 13812 7708 13864
rect 9036 13812 9088 13864
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 15384 14016 15436 14068
rect 18696 14016 18748 14068
rect 19064 14016 19116 14068
rect 16488 13948 16540 14000
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 18696 13855 18748 13864
rect 18696 13821 18705 13855
rect 18705 13821 18739 13855
rect 18739 13821 18748 13855
rect 18696 13812 18748 13821
rect 2780 13719 2832 13728
rect 2780 13685 2789 13719
rect 2789 13685 2823 13719
rect 2823 13685 2832 13719
rect 2780 13676 2832 13685
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 4068 13676 4120 13728
rect 4252 13676 4304 13728
rect 12900 13744 12952 13796
rect 15568 13744 15620 13796
rect 15752 13744 15804 13796
rect 18144 13787 18196 13796
rect 18144 13753 18162 13787
rect 18162 13753 18196 13787
rect 18144 13744 18196 13753
rect 18328 13744 18380 13796
rect 20260 13744 20312 13796
rect 24492 13812 24544 13864
rect 25044 13855 25096 13864
rect 25044 13821 25053 13855
rect 25053 13821 25087 13855
rect 25087 13821 25096 13855
rect 25044 13812 25096 13821
rect 25136 13855 25188 13864
rect 25136 13821 25150 13855
rect 25150 13821 25184 13855
rect 25184 13821 25188 13855
rect 25136 13812 25188 13821
rect 23296 13744 23348 13796
rect 24400 13744 24452 13796
rect 24952 13787 25004 13796
rect 24952 13753 24961 13787
rect 24961 13753 24995 13787
rect 24995 13753 25004 13787
rect 24952 13744 25004 13753
rect 4988 13676 5040 13728
rect 6368 13676 6420 13728
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 11520 13676 11572 13728
rect 14740 13676 14792 13728
rect 20076 13719 20128 13728
rect 20076 13685 20085 13719
rect 20085 13685 20119 13719
rect 20119 13685 20128 13719
rect 20076 13676 20128 13685
rect 20536 13676 20588 13728
rect 20628 13676 20680 13728
rect 24860 13676 24912 13728
rect 25596 13676 25648 13728
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 2780 13472 2832 13524
rect 2872 13472 2924 13524
rect 3056 13472 3108 13524
rect 7656 13404 7708 13456
rect 4160 13379 4212 13388
rect 4160 13345 4169 13379
rect 4169 13345 4203 13379
rect 4203 13345 4212 13379
rect 4160 13336 4212 13345
rect 4252 13336 4304 13388
rect 4712 13336 4764 13388
rect 8024 13336 8076 13388
rect 8760 13336 8812 13388
rect 9864 13336 9916 13388
rect 10600 13472 10652 13524
rect 10324 13447 10376 13456
rect 10324 13413 10333 13447
rect 10333 13413 10367 13447
rect 10367 13413 10376 13447
rect 10324 13404 10376 13413
rect 10784 13336 10836 13388
rect 11244 13379 11296 13388
rect 11244 13345 11278 13379
rect 11278 13345 11296 13379
rect 11244 13336 11296 13345
rect 11612 13336 11664 13388
rect 12716 13447 12768 13456
rect 12716 13413 12725 13447
rect 12725 13413 12759 13447
rect 12759 13413 12768 13447
rect 12716 13404 12768 13413
rect 15568 13472 15620 13524
rect 6920 13268 6972 13320
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 12716 13268 12768 13320
rect 13636 13336 13688 13388
rect 14096 13336 14148 13388
rect 24860 13472 24912 13524
rect 25136 13472 25188 13524
rect 12900 13200 12952 13252
rect 3516 13175 3568 13184
rect 3516 13141 3525 13175
rect 3525 13141 3559 13175
rect 3559 13141 3568 13175
rect 3516 13132 3568 13141
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 4804 13132 4856 13184
rect 5356 13132 5408 13184
rect 6644 13175 6696 13184
rect 6644 13141 6653 13175
rect 6653 13141 6687 13175
rect 6687 13141 6696 13175
rect 6644 13132 6696 13141
rect 10600 13132 10652 13184
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 12348 13175 12400 13184
rect 12348 13141 12357 13175
rect 12357 13141 12391 13175
rect 12391 13141 12400 13175
rect 12348 13132 12400 13141
rect 12992 13175 13044 13184
rect 12992 13141 13001 13175
rect 13001 13141 13035 13175
rect 13035 13141 13044 13175
rect 12992 13132 13044 13141
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 15384 13379 15436 13388
rect 15384 13345 15393 13379
rect 15393 13345 15427 13379
rect 15427 13345 15436 13379
rect 15384 13336 15436 13345
rect 15844 13336 15896 13388
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 16488 13336 16540 13388
rect 20352 13404 20404 13456
rect 20444 13447 20496 13456
rect 20444 13413 20453 13447
rect 20453 13413 20487 13447
rect 20487 13413 20496 13447
rect 20444 13404 20496 13413
rect 23204 13404 23256 13456
rect 18696 13336 18748 13388
rect 18788 13379 18840 13388
rect 18788 13345 18797 13379
rect 18797 13345 18831 13379
rect 18831 13345 18840 13379
rect 18788 13336 18840 13345
rect 18972 13379 19024 13388
rect 18972 13345 18981 13379
rect 18981 13345 19015 13379
rect 19015 13345 19024 13379
rect 18972 13336 19024 13345
rect 15568 13268 15620 13320
rect 19156 13379 19208 13388
rect 19156 13345 19165 13379
rect 19165 13345 19199 13379
rect 19199 13345 19208 13379
rect 19156 13336 19208 13345
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 20260 13379 20312 13388
rect 20260 13345 20270 13379
rect 20270 13345 20304 13379
rect 20304 13345 20312 13379
rect 20260 13336 20312 13345
rect 20536 13379 20588 13388
rect 20536 13345 20545 13379
rect 20545 13345 20579 13379
rect 20579 13345 20588 13379
rect 20536 13336 20588 13345
rect 20628 13379 20680 13388
rect 20628 13345 20642 13379
rect 20642 13345 20676 13379
rect 20676 13345 20680 13379
rect 20628 13336 20680 13345
rect 22008 13379 22060 13388
rect 22008 13345 22042 13379
rect 22042 13345 22060 13379
rect 22008 13336 22060 13345
rect 15660 13200 15712 13252
rect 14648 13132 14700 13184
rect 14924 13132 14976 13184
rect 20720 13268 20772 13320
rect 21272 13268 21324 13320
rect 23480 13379 23532 13388
rect 23480 13345 23514 13379
rect 23514 13345 23532 13379
rect 23480 13336 23532 13345
rect 26240 13404 26292 13456
rect 25136 13379 25188 13388
rect 25136 13345 25159 13379
rect 25159 13345 25188 13379
rect 25136 13336 25188 13345
rect 26148 13336 26200 13388
rect 17132 13132 17184 13184
rect 17316 13132 17368 13184
rect 21640 13200 21692 13252
rect 19340 13175 19392 13184
rect 19340 13141 19349 13175
rect 19349 13141 19383 13175
rect 19383 13141 19392 13175
rect 19340 13132 19392 13141
rect 19524 13132 19576 13184
rect 20628 13132 20680 13184
rect 20812 13175 20864 13184
rect 20812 13141 20821 13175
rect 20821 13141 20855 13175
rect 20855 13141 20864 13175
rect 20812 13132 20864 13141
rect 23112 13175 23164 13184
rect 23112 13141 23121 13175
rect 23121 13141 23155 13175
rect 23155 13141 23164 13175
rect 23112 13132 23164 13141
rect 23388 13132 23440 13184
rect 23940 13132 23992 13184
rect 24584 13175 24636 13184
rect 24584 13141 24593 13175
rect 24593 13141 24627 13175
rect 24627 13141 24636 13175
rect 24584 13132 24636 13141
rect 27804 13200 27856 13252
rect 26884 13132 26936 13184
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 11704 12928 11756 12980
rect 12716 12928 12768 12980
rect 13084 12928 13136 12980
rect 14004 12928 14056 12980
rect 11612 12860 11664 12912
rect 4160 12792 4212 12844
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 12808 12860 12860 12912
rect 6000 12724 6052 12776
rect 4160 12656 4212 12708
rect 5080 12656 5132 12708
rect 6828 12724 6880 12776
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 7748 12724 7800 12776
rect 6920 12656 6972 12708
rect 7472 12656 7524 12708
rect 10692 12724 10744 12776
rect 11520 12767 11572 12776
rect 11520 12733 11530 12767
rect 11530 12733 11564 12767
rect 11564 12733 11572 12767
rect 11520 12724 11572 12733
rect 11704 12767 11756 12776
rect 11704 12733 11713 12767
rect 11713 12733 11747 12767
rect 11747 12733 11756 12767
rect 11704 12724 11756 12733
rect 12348 12792 12400 12844
rect 16488 12928 16540 12980
rect 18788 12928 18840 12980
rect 19340 12928 19392 12980
rect 12072 12724 12124 12776
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 15844 12860 15896 12912
rect 17040 12860 17092 12912
rect 18144 12860 18196 12912
rect 19524 12860 19576 12912
rect 13084 12724 13136 12733
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 13728 12724 13780 12776
rect 16212 12835 16264 12844
rect 16212 12801 16221 12835
rect 16221 12801 16255 12835
rect 16255 12801 16264 12835
rect 16212 12792 16264 12801
rect 3608 12588 3660 12640
rect 5448 12631 5500 12640
rect 5448 12597 5457 12631
rect 5457 12597 5491 12631
rect 5491 12597 5500 12631
rect 5448 12588 5500 12597
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 5908 12588 5960 12640
rect 7104 12588 7156 12640
rect 7840 12588 7892 12640
rect 9680 12588 9732 12640
rect 12072 12631 12124 12640
rect 12072 12597 12081 12631
rect 12081 12597 12115 12631
rect 12115 12597 12124 12631
rect 12072 12588 12124 12597
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 13544 12588 13596 12640
rect 14096 12588 14148 12640
rect 14648 12631 14700 12640
rect 14648 12597 14657 12631
rect 14657 12597 14691 12631
rect 14691 12597 14700 12631
rect 14648 12588 14700 12597
rect 15844 12656 15896 12708
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 16580 12656 16632 12708
rect 16764 12699 16816 12708
rect 16764 12665 16773 12699
rect 16773 12665 16807 12699
rect 16807 12665 16816 12699
rect 16764 12656 16816 12665
rect 16304 12631 16356 12640
rect 16304 12597 16313 12631
rect 16313 12597 16347 12631
rect 16347 12597 16356 12631
rect 16304 12588 16356 12597
rect 17868 12656 17920 12708
rect 18420 12656 18472 12708
rect 19064 12656 19116 12708
rect 20812 12928 20864 12980
rect 22008 12928 22060 12980
rect 23112 12928 23164 12980
rect 23480 12971 23532 12980
rect 23480 12937 23489 12971
rect 23489 12937 23523 12971
rect 23523 12937 23532 12971
rect 23480 12928 23532 12937
rect 24492 12971 24544 12980
rect 24492 12937 24501 12971
rect 24501 12937 24535 12971
rect 24535 12937 24544 12971
rect 24492 12928 24544 12937
rect 25136 12928 25188 12980
rect 21640 12860 21692 12912
rect 22928 12860 22980 12912
rect 20996 12656 21048 12708
rect 21732 12767 21784 12776
rect 21732 12733 21741 12767
rect 21741 12733 21775 12767
rect 21775 12733 21784 12767
rect 21732 12724 21784 12733
rect 23020 12792 23072 12844
rect 23848 12860 23900 12912
rect 23296 12767 23348 12776
rect 23296 12733 23305 12767
rect 23305 12733 23339 12767
rect 23339 12733 23348 12767
rect 23296 12724 23348 12733
rect 24584 12792 24636 12844
rect 24308 12767 24360 12776
rect 24308 12733 24317 12767
rect 24317 12733 24351 12767
rect 24351 12733 24360 12767
rect 24308 12724 24360 12733
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 25964 12724 26016 12776
rect 26884 12767 26936 12776
rect 26884 12733 26893 12767
rect 26893 12733 26927 12767
rect 26927 12733 26936 12767
rect 26884 12724 26936 12733
rect 27068 12767 27120 12776
rect 27068 12733 27075 12767
rect 27075 12733 27120 12767
rect 27068 12724 27120 12733
rect 22376 12631 22428 12640
rect 22376 12597 22385 12631
rect 22385 12597 22419 12631
rect 22419 12597 22428 12631
rect 22376 12588 22428 12597
rect 24032 12656 24084 12708
rect 26424 12656 26476 12708
rect 27252 12699 27304 12708
rect 27252 12665 27261 12699
rect 27261 12665 27295 12699
rect 27295 12665 27304 12699
rect 27252 12656 27304 12665
rect 24860 12588 24912 12640
rect 26240 12588 26292 12640
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 4160 12384 4212 12436
rect 4620 12384 4672 12436
rect 5172 12384 5224 12436
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 5724 12384 5776 12436
rect 6828 12384 6880 12436
rect 6920 12384 6972 12436
rect 7472 12384 7524 12436
rect 3516 12316 3568 12368
rect 4620 12291 4672 12300
rect 4620 12257 4635 12291
rect 4635 12257 4669 12291
rect 4669 12257 4672 12291
rect 4620 12248 4672 12257
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 4896 12291 4948 12300
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 5540 12359 5592 12368
rect 5540 12325 5549 12359
rect 5549 12325 5583 12359
rect 5583 12325 5592 12359
rect 5540 12316 5592 12325
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 4068 12180 4120 12232
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 5356 12248 5408 12300
rect 5816 12281 5868 12300
rect 5816 12248 5825 12281
rect 5825 12248 5859 12281
rect 5859 12248 5868 12281
rect 6000 12248 6052 12300
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 6644 12291 6696 12300
rect 6644 12257 6653 12291
rect 6653 12257 6687 12291
rect 6687 12257 6696 12291
rect 6644 12248 6696 12257
rect 4804 12155 4856 12164
rect 4804 12121 4813 12155
rect 4813 12121 4847 12155
rect 4847 12121 4856 12155
rect 4804 12112 4856 12121
rect 5264 12112 5316 12164
rect 5816 12112 5868 12164
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 7012 12248 7064 12300
rect 7288 12291 7340 12300
rect 7288 12257 7297 12291
rect 7297 12257 7331 12291
rect 7331 12257 7340 12291
rect 7288 12248 7340 12257
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 11244 12384 11296 12436
rect 12532 12384 12584 12436
rect 13268 12427 13320 12436
rect 13268 12393 13277 12427
rect 13277 12393 13311 12427
rect 13311 12393 13320 12427
rect 13268 12384 13320 12393
rect 9680 12359 9732 12368
rect 9680 12325 9714 12359
rect 9714 12325 9732 12359
rect 9680 12316 9732 12325
rect 9864 12316 9916 12368
rect 11520 12316 11572 12368
rect 8024 12248 8076 12300
rect 8668 12248 8720 12300
rect 12072 12316 12124 12368
rect 12624 12359 12676 12368
rect 12624 12325 12633 12359
rect 12633 12325 12667 12359
rect 12667 12325 12676 12359
rect 12624 12316 12676 12325
rect 13176 12316 13228 12368
rect 6920 12112 6972 12164
rect 3608 12044 3660 12053
rect 6644 12044 6696 12096
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 11704 12180 11756 12232
rect 12808 12291 12860 12300
rect 12808 12257 12817 12291
rect 12817 12257 12851 12291
rect 12851 12257 12860 12291
rect 12808 12248 12860 12257
rect 13728 12384 13780 12436
rect 14004 12384 14056 12436
rect 16212 12427 16264 12436
rect 16212 12393 16221 12427
rect 16221 12393 16255 12427
rect 16255 12393 16264 12427
rect 16212 12384 16264 12393
rect 16304 12384 16356 12436
rect 14648 12316 14700 12368
rect 14832 12316 14884 12368
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 12440 12112 12492 12164
rect 12808 12112 12860 12164
rect 13084 12112 13136 12164
rect 13268 12112 13320 12164
rect 9588 12044 9640 12096
rect 9680 12044 9732 12096
rect 10692 12044 10744 12096
rect 10784 12087 10836 12096
rect 10784 12053 10793 12087
rect 10793 12053 10827 12087
rect 10827 12053 10836 12087
rect 10784 12044 10836 12053
rect 11520 12044 11572 12096
rect 15476 12087 15528 12096
rect 15476 12053 15485 12087
rect 15485 12053 15519 12087
rect 15519 12053 15528 12087
rect 15476 12044 15528 12053
rect 15844 12248 15896 12300
rect 16304 12291 16356 12300
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 16396 12248 16448 12300
rect 16580 12291 16632 12300
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 17868 12427 17920 12436
rect 17868 12393 17877 12427
rect 17877 12393 17911 12427
rect 17911 12393 17920 12427
rect 17868 12384 17920 12393
rect 17040 12291 17092 12300
rect 17040 12257 17049 12291
rect 17049 12257 17083 12291
rect 17083 12257 17092 12291
rect 17040 12248 17092 12257
rect 18696 12248 18748 12300
rect 17868 12180 17920 12232
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 17960 12112 18012 12164
rect 18880 12180 18932 12232
rect 19432 12248 19484 12300
rect 20076 12248 20128 12300
rect 20260 12248 20312 12300
rect 19892 12180 19944 12232
rect 19248 12044 19300 12096
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 21088 12291 21140 12300
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 21364 12248 21416 12300
rect 21640 12291 21692 12300
rect 21640 12257 21649 12291
rect 21649 12257 21683 12291
rect 21683 12257 21692 12291
rect 21640 12248 21692 12257
rect 21732 12248 21784 12300
rect 21456 12112 21508 12164
rect 22008 12291 22060 12300
rect 22008 12257 22017 12291
rect 22017 12257 22051 12291
rect 22051 12257 22060 12291
rect 22008 12248 22060 12257
rect 21824 12180 21876 12232
rect 22376 12316 22428 12368
rect 22560 12248 22612 12300
rect 22744 12291 22796 12300
rect 22744 12257 22753 12291
rect 22753 12257 22787 12291
rect 22787 12257 22796 12291
rect 22744 12248 22796 12257
rect 23020 12248 23072 12300
rect 23204 12291 23256 12300
rect 23204 12257 23213 12291
rect 23213 12257 23247 12291
rect 23247 12257 23256 12291
rect 23204 12248 23256 12257
rect 23848 12316 23900 12368
rect 23572 12248 23624 12300
rect 24124 12291 24176 12300
rect 24124 12257 24158 12291
rect 24158 12257 24176 12291
rect 24124 12248 24176 12257
rect 23848 12223 23900 12232
rect 23848 12189 23857 12223
rect 23857 12189 23891 12223
rect 23891 12189 23900 12223
rect 23848 12180 23900 12189
rect 25044 12316 25096 12368
rect 27252 12384 27304 12436
rect 25228 12248 25280 12300
rect 25504 12248 25556 12300
rect 25780 12291 25832 12300
rect 25780 12257 25794 12291
rect 25794 12257 25828 12291
rect 25828 12257 25832 12291
rect 25780 12248 25832 12257
rect 26148 12248 26200 12300
rect 27712 12248 27764 12300
rect 29276 12223 29328 12232
rect 29276 12189 29285 12223
rect 29285 12189 29319 12223
rect 29319 12189 29328 12223
rect 29276 12180 29328 12189
rect 19524 12044 19576 12096
rect 20260 12044 20312 12096
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 21272 12044 21324 12096
rect 22836 12044 22888 12096
rect 23204 12087 23256 12096
rect 23204 12053 23213 12087
rect 23213 12053 23247 12087
rect 23247 12053 23256 12087
rect 23204 12044 23256 12053
rect 23480 12087 23532 12096
rect 23480 12053 23489 12087
rect 23489 12053 23523 12087
rect 23523 12053 23532 12087
rect 23480 12044 23532 12053
rect 26332 12044 26384 12096
rect 27068 12044 27120 12096
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 5172 11840 5224 11892
rect 6092 11840 6144 11892
rect 7564 11840 7616 11892
rect 8668 11883 8720 11892
rect 8668 11849 8677 11883
rect 8677 11849 8711 11883
rect 8711 11849 8720 11883
rect 8668 11840 8720 11849
rect 11796 11840 11848 11892
rect 11888 11840 11940 11892
rect 12716 11840 12768 11892
rect 4712 11772 4764 11824
rect 6644 11772 6696 11824
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 4620 11704 4672 11756
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 7748 11772 7800 11824
rect 8576 11772 8628 11824
rect 9220 11772 9272 11824
rect 11060 11772 11112 11824
rect 11244 11772 11296 11824
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 10784 11704 10836 11756
rect 3516 11500 3568 11552
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 4988 11568 5040 11620
rect 5264 11568 5316 11620
rect 6736 11543 6788 11552
rect 6736 11509 6745 11543
rect 6745 11509 6779 11543
rect 6779 11509 6788 11543
rect 6736 11500 6788 11509
rect 7564 11568 7616 11620
rect 9588 11636 9640 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 11060 11679 11112 11688
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 9404 11568 9456 11620
rect 11888 11636 11940 11688
rect 12532 11704 12584 11756
rect 12992 11704 13044 11756
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 11336 11611 11388 11620
rect 11336 11577 11345 11611
rect 11345 11577 11379 11611
rect 11379 11577 11388 11611
rect 11336 11568 11388 11577
rect 11796 11611 11848 11620
rect 11796 11577 11805 11611
rect 11805 11577 11839 11611
rect 11839 11577 11848 11611
rect 11796 11568 11848 11577
rect 12440 11636 12492 11688
rect 12624 11679 12676 11688
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 13820 11636 13872 11688
rect 18236 11840 18288 11892
rect 18512 11840 18564 11892
rect 19156 11883 19208 11892
rect 19156 11849 19165 11883
rect 19165 11849 19199 11883
rect 19199 11849 19208 11883
rect 19156 11840 19208 11849
rect 15476 11636 15528 11688
rect 15844 11636 15896 11688
rect 7656 11500 7708 11552
rect 7932 11500 7984 11552
rect 9680 11500 9732 11552
rect 9864 11500 9916 11552
rect 10692 11500 10744 11552
rect 16396 11636 16448 11688
rect 17868 11679 17920 11688
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 18144 11772 18196 11824
rect 20076 11840 20128 11892
rect 20260 11840 20312 11892
rect 21088 11840 21140 11892
rect 21456 11840 21508 11892
rect 22008 11840 22060 11892
rect 23296 11883 23348 11892
rect 19524 11772 19576 11824
rect 22744 11772 22796 11824
rect 23296 11849 23305 11883
rect 23305 11849 23339 11883
rect 23339 11849 23348 11883
rect 23296 11840 23348 11849
rect 23480 11840 23532 11892
rect 24124 11840 24176 11892
rect 27712 11883 27764 11892
rect 27712 11849 27721 11883
rect 27721 11849 27755 11883
rect 27755 11849 27764 11883
rect 27712 11840 27764 11849
rect 23112 11772 23164 11824
rect 18144 11679 18196 11688
rect 18144 11645 18153 11679
rect 18153 11645 18187 11679
rect 18187 11645 18196 11679
rect 18144 11636 18196 11645
rect 18880 11636 18932 11688
rect 19248 11636 19300 11688
rect 19432 11636 19484 11688
rect 12072 11543 12124 11552
rect 12072 11509 12081 11543
rect 12081 11509 12115 11543
rect 12115 11509 12124 11543
rect 12072 11500 12124 11509
rect 12440 11500 12492 11552
rect 13820 11500 13872 11552
rect 14280 11500 14332 11552
rect 15384 11500 15436 11552
rect 15476 11500 15528 11552
rect 18052 11568 18104 11620
rect 19892 11679 19944 11688
rect 17684 11500 17736 11552
rect 19892 11645 19901 11679
rect 19901 11645 19935 11679
rect 19935 11645 19944 11679
rect 19892 11636 19944 11645
rect 22192 11636 22244 11688
rect 22928 11704 22980 11756
rect 22744 11679 22796 11688
rect 22744 11645 22753 11679
rect 22753 11645 22787 11679
rect 22787 11645 22796 11679
rect 22744 11636 22796 11645
rect 23664 11704 23716 11756
rect 23204 11636 23256 11688
rect 23572 11636 23624 11688
rect 20168 11611 20220 11620
rect 20168 11577 20202 11611
rect 20202 11577 20220 11611
rect 20168 11568 20220 11577
rect 20260 11500 20312 11552
rect 21824 11500 21876 11552
rect 22560 11543 22612 11552
rect 22560 11509 22569 11543
rect 22569 11509 22603 11543
rect 22603 11509 22612 11543
rect 22560 11500 22612 11509
rect 23020 11568 23072 11620
rect 22836 11500 22888 11552
rect 26240 11679 26292 11688
rect 26240 11645 26249 11679
rect 26249 11645 26283 11679
rect 26283 11645 26292 11679
rect 26240 11636 26292 11645
rect 26332 11636 26384 11688
rect 26700 11679 26752 11688
rect 26700 11645 26709 11679
rect 26709 11645 26743 11679
rect 26743 11645 26752 11679
rect 26700 11636 26752 11645
rect 27252 11679 27304 11688
rect 27252 11645 27261 11679
rect 27261 11645 27295 11679
rect 27295 11645 27304 11679
rect 27252 11636 27304 11645
rect 26148 11543 26200 11552
rect 26148 11509 26157 11543
rect 26157 11509 26191 11543
rect 26191 11509 26200 11543
rect 26148 11500 26200 11509
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 3424 11296 3476 11348
rect 3976 11296 4028 11348
rect 4620 11296 4672 11348
rect 4988 11339 5040 11348
rect 4988 11305 4997 11339
rect 4997 11305 5031 11339
rect 5031 11305 5040 11339
rect 4988 11296 5040 11305
rect 6000 11296 6052 11348
rect 7104 11296 7156 11348
rect 7288 11296 7340 11348
rect 7748 11296 7800 11348
rect 8300 11296 8352 11348
rect 3792 11228 3844 11280
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 3240 11092 3292 11144
rect 7840 11092 7892 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8208 11160 8260 11212
rect 8300 11203 8352 11212
rect 8300 11169 8309 11203
rect 8309 11169 8343 11203
rect 8343 11169 8352 11203
rect 8300 11160 8352 11169
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 8760 11203 8812 11212
rect 8760 11169 8769 11203
rect 8769 11169 8803 11203
rect 8803 11169 8812 11203
rect 8760 11160 8812 11169
rect 9036 11160 9088 11212
rect 9220 11228 9272 11280
rect 9404 11296 9456 11348
rect 10692 11296 10744 11348
rect 11796 11296 11848 11348
rect 12072 11296 12124 11348
rect 5172 10956 5224 11008
rect 5908 10956 5960 11008
rect 7932 10956 7984 11008
rect 8484 11024 8536 11076
rect 10600 11160 10652 11212
rect 11244 11203 11296 11212
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 8116 10956 8168 11008
rect 8300 10956 8352 11008
rect 8668 10956 8720 11008
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 11428 11160 11480 11212
rect 12440 11160 12492 11212
rect 13176 11296 13228 11348
rect 13820 11296 13872 11348
rect 16120 11296 16172 11348
rect 13360 11160 13412 11212
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 11428 10956 11480 11008
rect 11520 10956 11572 11008
rect 15108 11160 15160 11212
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 15292 11160 15344 11212
rect 16304 11228 16356 11280
rect 16396 11228 16448 11280
rect 16488 11271 16540 11280
rect 16488 11237 16497 11271
rect 16497 11237 16531 11271
rect 16531 11237 16540 11271
rect 16488 11228 16540 11237
rect 15476 11024 15528 11076
rect 18052 11296 18104 11348
rect 18144 11296 18196 11348
rect 19524 11296 19576 11348
rect 20168 11296 20220 11348
rect 20260 11296 20312 11348
rect 20628 11296 20680 11348
rect 21456 11296 21508 11348
rect 17224 11203 17276 11212
rect 17224 11169 17233 11203
rect 17233 11169 17267 11203
rect 17267 11169 17276 11203
rect 17224 11160 17276 11169
rect 17960 11160 18012 11212
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 21272 11160 21324 11212
rect 22836 11296 22888 11348
rect 22928 11296 22980 11348
rect 23020 11296 23072 11348
rect 22560 11228 22612 11280
rect 22192 11203 22244 11212
rect 22192 11169 22201 11203
rect 22201 11169 22235 11203
rect 22235 11169 22244 11203
rect 22192 11160 22244 11169
rect 20812 11092 20864 11144
rect 22836 11203 22888 11212
rect 22836 11169 22845 11203
rect 22845 11169 22879 11203
rect 22879 11169 22888 11203
rect 22836 11160 22888 11169
rect 20168 11024 20220 11076
rect 23020 11092 23072 11144
rect 25228 11160 25280 11212
rect 25780 11271 25832 11280
rect 25780 11237 25789 11271
rect 25789 11237 25823 11271
rect 25823 11237 25832 11271
rect 25780 11228 25832 11237
rect 26148 11228 26200 11280
rect 25964 11203 26016 11212
rect 25964 11169 25978 11203
rect 25978 11169 26012 11203
rect 26012 11169 26016 11203
rect 25964 11160 26016 11169
rect 28080 11160 28132 11212
rect 29276 11160 29328 11212
rect 23664 11092 23716 11144
rect 23848 11092 23900 11144
rect 27988 11092 28040 11144
rect 29000 11092 29052 11144
rect 15108 10999 15160 11008
rect 15108 10965 15117 10999
rect 15117 10965 15151 10999
rect 15151 10965 15160 10999
rect 15108 10956 15160 10965
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 16488 10956 16540 11008
rect 18788 10956 18840 11008
rect 21088 10956 21140 11008
rect 23020 10999 23072 11008
rect 23020 10965 23029 10999
rect 23029 10965 23063 10999
rect 23063 10965 23072 10999
rect 23020 10956 23072 10965
rect 23112 10999 23164 11008
rect 23112 10965 23121 10999
rect 23121 10965 23155 10999
rect 23155 10965 23164 10999
rect 23112 10956 23164 10965
rect 26148 10999 26200 11008
rect 26148 10965 26157 10999
rect 26157 10965 26191 10999
rect 26191 10965 26200 10999
rect 26148 10956 26200 10965
rect 27160 10956 27212 11008
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 848 10591 900 10600
rect 848 10557 857 10591
rect 857 10557 891 10591
rect 891 10557 900 10591
rect 848 10548 900 10557
rect 10140 10752 10192 10804
rect 10600 10752 10652 10804
rect 5264 10616 5316 10668
rect 7748 10616 7800 10668
rect 7932 10616 7984 10668
rect 8760 10616 8812 10668
rect 10692 10684 10744 10736
rect 15752 10752 15804 10804
rect 18236 10752 18288 10804
rect 22284 10752 22336 10804
rect 3516 10548 3568 10600
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 5908 10591 5960 10600
rect 5908 10557 5942 10591
rect 5942 10557 5960 10591
rect 5908 10548 5960 10557
rect 7840 10548 7892 10600
rect 4988 10455 5040 10464
rect 4988 10421 4997 10455
rect 4997 10421 5031 10455
rect 5031 10421 5040 10455
rect 4988 10412 5040 10421
rect 8484 10480 8536 10532
rect 10784 10548 10836 10600
rect 11152 10548 11204 10600
rect 11520 10616 11572 10668
rect 11428 10591 11480 10600
rect 11428 10557 11437 10591
rect 11437 10557 11471 10591
rect 11471 10557 11480 10591
rect 11428 10548 11480 10557
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 10600 10412 10652 10464
rect 11520 10480 11572 10532
rect 14004 10548 14056 10600
rect 20720 10684 20772 10736
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 15384 10616 15436 10668
rect 16120 10616 16172 10668
rect 14740 10548 14792 10600
rect 14924 10548 14976 10600
rect 15384 10480 15436 10532
rect 18420 10480 18472 10532
rect 18788 10548 18840 10600
rect 20812 10548 20864 10600
rect 25596 10659 25648 10668
rect 25596 10625 25605 10659
rect 25605 10625 25639 10659
rect 25639 10625 25648 10659
rect 25596 10616 25648 10625
rect 21732 10591 21784 10600
rect 21732 10557 21741 10591
rect 21741 10557 21775 10591
rect 21775 10557 21784 10591
rect 21732 10548 21784 10557
rect 21824 10548 21876 10600
rect 23020 10548 23072 10600
rect 23664 10591 23716 10600
rect 23664 10557 23673 10591
rect 23673 10557 23707 10591
rect 23707 10557 23716 10591
rect 23664 10548 23716 10557
rect 25136 10591 25188 10600
rect 25136 10557 25145 10591
rect 25145 10557 25179 10591
rect 25179 10557 25188 10591
rect 25136 10548 25188 10557
rect 25320 10591 25372 10600
rect 25320 10557 25329 10591
rect 25329 10557 25363 10591
rect 25363 10557 25372 10591
rect 25320 10548 25372 10557
rect 26148 10548 26200 10600
rect 14280 10412 14332 10464
rect 14648 10412 14700 10464
rect 15476 10412 15528 10464
rect 15568 10412 15620 10464
rect 16212 10412 16264 10464
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 20076 10412 20128 10421
rect 20904 10455 20956 10464
rect 20904 10421 20913 10455
rect 20913 10421 20947 10455
rect 20947 10421 20956 10455
rect 20904 10412 20956 10421
rect 21364 10455 21416 10464
rect 21364 10421 21373 10455
rect 21373 10421 21407 10455
rect 21407 10421 21416 10455
rect 21364 10412 21416 10421
rect 23112 10480 23164 10532
rect 31668 10480 31720 10532
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 4988 10208 5040 10260
rect 3148 10140 3200 10192
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 6736 10140 6788 10192
rect 5264 10072 5316 10124
rect 7196 10072 7248 10124
rect 8852 10140 8904 10192
rect 9680 10183 9732 10192
rect 9680 10149 9689 10183
rect 9689 10149 9723 10183
rect 9723 10149 9732 10183
rect 9680 10140 9732 10149
rect 9772 10183 9824 10192
rect 9772 10149 9781 10183
rect 9781 10149 9815 10183
rect 9815 10149 9824 10183
rect 9772 10140 9824 10149
rect 10692 10140 10744 10192
rect 7932 10115 7984 10124
rect 7932 10081 7966 10115
rect 7966 10081 7984 10115
rect 7932 10072 7984 10081
rect 8484 10072 8536 10124
rect 9220 10072 9272 10124
rect 9864 10115 9916 10124
rect 9864 10081 9878 10115
rect 9878 10081 9912 10115
rect 9912 10081 9916 10115
rect 9864 10072 9916 10081
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 10232 10072 10284 10124
rect 10600 10072 10652 10124
rect 12348 10140 12400 10192
rect 12992 10140 13044 10192
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 11520 10072 11572 10124
rect 14188 10208 14240 10260
rect 14556 10208 14608 10260
rect 15384 10208 15436 10260
rect 15568 10208 15620 10260
rect 16396 10208 16448 10260
rect 20076 10208 20128 10260
rect 20352 10251 20404 10260
rect 20352 10217 20361 10251
rect 20361 10217 20395 10251
rect 20395 10217 20404 10251
rect 20352 10208 20404 10217
rect 20904 10208 20956 10260
rect 21180 10208 21232 10260
rect 14004 10140 14056 10192
rect 14280 10072 14332 10124
rect 14740 10072 14792 10124
rect 16212 10115 16264 10124
rect 16212 10081 16221 10115
rect 16221 10081 16255 10115
rect 16255 10081 16264 10115
rect 16212 10072 16264 10081
rect 19432 10072 19484 10124
rect 10876 9936 10928 9988
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 18972 10004 19024 10056
rect 19156 10047 19208 10056
rect 19156 10013 19165 10047
rect 19165 10013 19199 10047
rect 19199 10013 19208 10047
rect 19156 10004 19208 10013
rect 16212 9936 16264 9988
rect 19984 9936 20036 9988
rect 16396 9868 16448 9920
rect 16580 9868 16632 9920
rect 20720 10115 20772 10124
rect 20720 10081 20729 10115
rect 20729 10081 20763 10115
rect 20763 10081 20772 10115
rect 20720 10072 20772 10081
rect 21364 10072 21416 10124
rect 22192 10208 22244 10260
rect 22284 10140 22336 10192
rect 22652 10072 22704 10124
rect 23112 10115 23164 10124
rect 23112 10081 23121 10115
rect 23121 10081 23155 10115
rect 23155 10081 23164 10115
rect 23112 10072 23164 10081
rect 23388 10115 23440 10124
rect 23388 10081 23422 10115
rect 23422 10081 23440 10115
rect 23388 10072 23440 10081
rect 25228 10140 25280 10192
rect 24860 10115 24912 10124
rect 24860 10081 24869 10115
rect 24869 10081 24903 10115
rect 24903 10081 24912 10115
rect 24860 10072 24912 10081
rect 25412 10115 25464 10124
rect 25412 10081 25421 10115
rect 25421 10081 25455 10115
rect 25455 10081 25464 10115
rect 25412 10072 25464 10081
rect 25596 10115 25648 10124
rect 25596 10081 25605 10115
rect 25605 10081 25639 10115
rect 25639 10081 25648 10115
rect 25596 10072 25648 10081
rect 26884 10115 26936 10124
rect 26884 10081 26918 10115
rect 26918 10081 26936 10115
rect 21180 10004 21232 10056
rect 24400 10004 24452 10056
rect 26884 10072 26936 10081
rect 27896 10072 27948 10124
rect 27988 10004 28040 10056
rect 22284 9868 22336 9920
rect 24676 9868 24728 9920
rect 25872 9911 25924 9920
rect 25872 9877 25881 9911
rect 25881 9877 25915 9911
rect 25915 9877 25924 9911
rect 25872 9868 25924 9877
rect 27988 9911 28040 9920
rect 27988 9877 27997 9911
rect 27997 9877 28031 9911
rect 28031 9877 28040 9911
rect 27988 9868 28040 9877
rect 29460 9911 29512 9920
rect 29460 9877 29469 9911
rect 29469 9877 29503 9911
rect 29503 9877 29512 9911
rect 29460 9868 29512 9877
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 3240 9596 3292 9648
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 9772 9664 9824 9716
rect 9864 9664 9916 9716
rect 14004 9664 14056 9716
rect 10600 9596 10652 9648
rect 11336 9596 11388 9648
rect 15660 9596 15712 9648
rect 5632 9460 5684 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 4804 9324 4856 9376
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 10876 9528 10928 9580
rect 12900 9528 12952 9580
rect 18144 9664 18196 9716
rect 20720 9664 20772 9716
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 11520 9460 11572 9512
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 15476 9503 15528 9512
rect 15476 9469 15485 9503
rect 15485 9469 15519 9503
rect 15519 9469 15528 9503
rect 15476 9460 15528 9469
rect 16580 9460 16632 9512
rect 17500 9460 17552 9512
rect 18604 9460 18656 9512
rect 18972 9460 19024 9512
rect 20168 9528 20220 9580
rect 20904 9596 20956 9648
rect 23388 9664 23440 9716
rect 25412 9664 25464 9716
rect 21732 9528 21784 9580
rect 21916 9528 21968 9580
rect 22192 9528 22244 9580
rect 24584 9596 24636 9648
rect 25780 9596 25832 9648
rect 26700 9664 26752 9716
rect 26884 9664 26936 9716
rect 27068 9664 27120 9716
rect 27896 9664 27948 9716
rect 27988 9664 28040 9716
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 9220 9324 9272 9376
rect 12256 9392 12308 9444
rect 17684 9392 17736 9444
rect 18420 9392 18472 9444
rect 19156 9392 19208 9444
rect 19984 9392 20036 9444
rect 9772 9324 9824 9376
rect 10968 9324 11020 9376
rect 11336 9324 11388 9376
rect 12900 9324 12952 9376
rect 13084 9324 13136 9376
rect 13636 9367 13688 9376
rect 13636 9333 13645 9367
rect 13645 9333 13679 9367
rect 13679 9333 13688 9367
rect 13636 9324 13688 9333
rect 14740 9324 14792 9376
rect 16764 9324 16816 9376
rect 19432 9324 19484 9376
rect 20628 9324 20680 9376
rect 21824 9435 21876 9444
rect 21824 9401 21833 9435
rect 21833 9401 21867 9435
rect 21867 9401 21876 9435
rect 21824 9392 21876 9401
rect 22192 9392 22244 9444
rect 24308 9528 24360 9580
rect 22376 9503 22428 9512
rect 22376 9469 22385 9503
rect 22385 9469 22419 9503
rect 22419 9469 22428 9503
rect 22376 9460 22428 9469
rect 22468 9503 22520 9512
rect 22468 9469 22477 9503
rect 22477 9469 22511 9503
rect 22511 9469 22520 9503
rect 22468 9460 22520 9469
rect 23020 9460 23072 9512
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 24492 9460 24544 9469
rect 24584 9503 24636 9512
rect 24584 9469 24593 9503
rect 24593 9469 24627 9503
rect 24627 9469 24636 9503
rect 24584 9460 24636 9469
rect 22468 9324 22520 9376
rect 24124 9324 24176 9376
rect 24676 9435 24728 9444
rect 24676 9401 24685 9435
rect 24685 9401 24719 9435
rect 24719 9401 24728 9435
rect 24676 9392 24728 9401
rect 25136 9460 25188 9512
rect 25964 9503 26016 9512
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 26056 9503 26108 9512
rect 26056 9469 26065 9503
rect 26065 9469 26099 9503
rect 26099 9469 26108 9503
rect 26056 9460 26108 9469
rect 26884 9460 26936 9512
rect 27344 9528 27396 9580
rect 26976 9324 27028 9376
rect 27436 9503 27488 9512
rect 27436 9469 27445 9503
rect 27445 9469 27479 9503
rect 27479 9469 27488 9503
rect 27436 9460 27488 9469
rect 27804 9460 27856 9512
rect 28080 9460 28132 9512
rect 29184 9503 29236 9512
rect 29184 9469 29193 9503
rect 29193 9469 29227 9503
rect 29227 9469 29236 9503
rect 29184 9460 29236 9469
rect 29460 9460 29512 9512
rect 29368 9435 29420 9444
rect 29368 9401 29377 9435
rect 29377 9401 29411 9435
rect 29411 9401 29420 9435
rect 29368 9392 29420 9401
rect 28080 9367 28132 9376
rect 28080 9333 28089 9367
rect 28089 9333 28123 9367
rect 28123 9333 28132 9367
rect 28080 9324 28132 9333
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 6000 9120 6052 9172
rect 7288 9120 7340 9172
rect 11336 9120 11388 9172
rect 3240 9027 3292 9036
rect 3240 8993 3249 9027
rect 3249 8993 3283 9027
rect 3283 8993 3292 9027
rect 3240 8984 3292 8993
rect 4988 8984 5040 9036
rect 7104 9052 7156 9104
rect 7196 9052 7248 9104
rect 10416 9095 10468 9104
rect 10416 9061 10425 9095
rect 10425 9061 10459 9095
rect 10459 9061 10468 9095
rect 10416 9052 10468 9061
rect 11152 9052 11204 9104
rect 11244 9052 11296 9104
rect 11612 9052 11664 9104
rect 9956 8984 10008 9036
rect 10140 8984 10192 9036
rect 13084 9095 13136 9104
rect 13084 9061 13093 9095
rect 13093 9061 13127 9095
rect 13127 9061 13136 9095
rect 13084 9052 13136 9061
rect 14556 9120 14608 9172
rect 15108 9120 15160 9172
rect 16488 9163 16540 9172
rect 16488 9129 16497 9163
rect 16497 9129 16531 9163
rect 16531 9129 16540 9163
rect 16488 9120 16540 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 12348 8984 12400 9036
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 12808 9027 12860 9036
rect 12808 8993 12817 9027
rect 12817 8993 12851 9027
rect 12851 8993 12860 9027
rect 12808 8984 12860 8993
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 13268 8984 13320 9036
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 13728 9027 13780 9036
rect 13728 8993 13737 9027
rect 13737 8993 13771 9027
rect 13771 8993 13780 9027
rect 13728 8984 13780 8993
rect 13820 8984 13872 9036
rect 14372 8984 14424 9036
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 15844 9052 15896 9104
rect 17132 9120 17184 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 17684 9163 17736 9172
rect 17684 9129 17693 9163
rect 17693 9129 17727 9163
rect 17727 9129 17736 9163
rect 17684 9120 17736 9129
rect 19340 9163 19392 9172
rect 19340 9129 19349 9163
rect 19349 9129 19383 9163
rect 19383 9129 19392 9163
rect 19340 9120 19392 9129
rect 19800 9120 19852 9172
rect 19984 9120 20036 9172
rect 20628 9120 20680 9172
rect 22376 9120 22428 9172
rect 15016 8984 15068 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 16212 8984 16264 9036
rect 17040 9052 17092 9104
rect 26332 9120 26384 9172
rect 4068 8916 4120 8968
rect 17592 8984 17644 9036
rect 17776 8984 17828 9036
rect 18328 8984 18380 9036
rect 18420 8959 18472 8968
rect 5724 8848 5776 8900
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 7288 8780 7340 8832
rect 7932 8780 7984 8832
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 11520 8780 11572 8832
rect 12256 8848 12308 8900
rect 13820 8848 13872 8900
rect 18420 8925 18429 8959
rect 18429 8925 18463 8959
rect 18463 8925 18472 8959
rect 18420 8916 18472 8925
rect 18604 8984 18656 9036
rect 18972 8916 19024 8968
rect 19432 9027 19484 9036
rect 19432 8993 19441 9027
rect 19441 8993 19475 9027
rect 19475 8993 19484 9027
rect 19432 8984 19484 8993
rect 20076 9027 20128 9036
rect 20076 8993 20085 9027
rect 20085 8993 20119 9027
rect 20119 8993 20128 9027
rect 20076 8984 20128 8993
rect 20904 8984 20956 9036
rect 21180 8984 21232 9036
rect 23020 9027 23072 9036
rect 23020 8993 23029 9027
rect 23029 8993 23063 9027
rect 23063 8993 23072 9027
rect 23020 8984 23072 8993
rect 23112 9027 23164 9036
rect 23112 8993 23121 9027
rect 23121 8993 23155 9027
rect 23155 8993 23164 9027
rect 23112 8984 23164 8993
rect 25596 9095 25648 9104
rect 25596 9061 25605 9095
rect 25605 9061 25639 9095
rect 25639 9061 25648 9095
rect 25596 9052 25648 9061
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 22836 8916 22888 8925
rect 15016 8780 15068 8832
rect 21088 8848 21140 8900
rect 23204 8848 23256 8900
rect 26424 8984 26476 9036
rect 26608 9052 26660 9104
rect 27068 9052 27120 9104
rect 26700 8984 26752 9036
rect 28080 9052 28132 9104
rect 29368 9052 29420 9104
rect 30012 9052 30064 9104
rect 24124 8959 24176 8968
rect 24124 8925 24133 8959
rect 24133 8925 24167 8959
rect 24167 8925 24176 8959
rect 24124 8916 24176 8925
rect 25228 8916 25280 8968
rect 26332 8916 26384 8968
rect 27988 8984 28040 9036
rect 29184 8984 29236 9036
rect 29736 8984 29788 9036
rect 30196 9027 30248 9036
rect 30196 8993 30205 9027
rect 30205 8993 30239 9027
rect 30239 8993 30248 9027
rect 30196 8984 30248 8993
rect 16856 8780 16908 8832
rect 19064 8780 19116 8832
rect 19616 8780 19668 8832
rect 22192 8780 22244 8832
rect 23664 8780 23716 8832
rect 26148 8848 26200 8900
rect 27804 8916 27856 8968
rect 28080 8916 28132 8968
rect 27068 8891 27120 8900
rect 24400 8780 24452 8832
rect 24492 8780 24544 8832
rect 26608 8780 26660 8832
rect 27068 8857 27077 8891
rect 27077 8857 27111 8891
rect 27111 8857 27120 8891
rect 27068 8848 27120 8857
rect 27344 8848 27396 8900
rect 27436 8891 27488 8900
rect 27436 8857 27445 8891
rect 27445 8857 27479 8891
rect 27479 8857 27488 8891
rect 27436 8848 27488 8857
rect 27528 8891 27580 8900
rect 27528 8857 27537 8891
rect 27537 8857 27571 8891
rect 27571 8857 27580 8891
rect 27528 8848 27580 8857
rect 27252 8780 27304 8832
rect 27896 8780 27948 8832
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 4804 8576 4856 8628
rect 4988 8619 5040 8628
rect 4988 8585 4997 8619
rect 4997 8585 5031 8619
rect 5031 8585 5040 8619
rect 4988 8576 5040 8585
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 7196 8576 7248 8628
rect 9036 8576 9088 8628
rect 11152 8576 11204 8628
rect 7012 8508 7064 8560
rect 4068 8372 4120 8424
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 6368 8440 6420 8492
rect 7104 8440 7156 8492
rect 13728 8576 13780 8628
rect 5908 8372 5960 8381
rect 6644 8372 6696 8424
rect 8484 8440 8536 8492
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 10232 8440 10284 8492
rect 10416 8440 10468 8492
rect 12072 8551 12124 8560
rect 12072 8517 12081 8551
rect 12081 8517 12115 8551
rect 12115 8517 12124 8551
rect 12072 8508 12124 8517
rect 12164 8551 12216 8560
rect 12164 8517 12173 8551
rect 12173 8517 12207 8551
rect 12207 8517 12216 8551
rect 19708 8576 19760 8628
rect 20076 8576 20128 8628
rect 21180 8619 21232 8628
rect 21180 8585 21189 8619
rect 21189 8585 21223 8619
rect 21223 8585 21232 8619
rect 21180 8576 21232 8585
rect 23020 8576 23072 8628
rect 12164 8508 12216 8517
rect 3240 8236 3292 8288
rect 6736 8304 6788 8356
rect 6920 8304 6972 8356
rect 9404 8372 9456 8424
rect 9956 8372 10008 8424
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 7380 8347 7432 8356
rect 7380 8313 7389 8347
rect 7389 8313 7423 8347
rect 7423 8313 7432 8347
rect 7380 8304 7432 8313
rect 11152 8415 11204 8424
rect 11152 8381 11161 8415
rect 11161 8381 11195 8415
rect 11195 8381 11204 8415
rect 11152 8372 11204 8381
rect 11336 8372 11388 8424
rect 12348 8440 12400 8492
rect 15476 8508 15528 8560
rect 10048 8236 10100 8288
rect 11152 8236 11204 8288
rect 12532 8372 12584 8424
rect 12072 8304 12124 8356
rect 13912 8372 13964 8424
rect 12808 8304 12860 8356
rect 14372 8372 14424 8424
rect 15844 8415 15896 8424
rect 15844 8381 15853 8415
rect 15853 8381 15887 8415
rect 15887 8381 15896 8415
rect 15844 8372 15896 8381
rect 17040 8508 17092 8560
rect 19340 8508 19392 8560
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 16488 8415 16540 8424
rect 16488 8381 16497 8415
rect 16497 8381 16531 8415
rect 16531 8381 16540 8415
rect 16488 8372 16540 8381
rect 16856 8372 16908 8424
rect 19524 8440 19576 8492
rect 19064 8415 19116 8424
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 19248 8415 19300 8424
rect 19248 8381 19257 8415
rect 19257 8381 19291 8415
rect 19291 8381 19300 8415
rect 19248 8372 19300 8381
rect 19340 8415 19392 8424
rect 19340 8381 19349 8415
rect 19349 8381 19383 8415
rect 19383 8381 19392 8415
rect 19340 8372 19392 8381
rect 17684 8304 17736 8356
rect 12164 8236 12216 8288
rect 12440 8236 12492 8288
rect 12532 8279 12584 8288
rect 12532 8245 12541 8279
rect 12541 8245 12575 8279
rect 12575 8245 12584 8279
rect 12532 8236 12584 8245
rect 16396 8236 16448 8288
rect 16580 8236 16632 8288
rect 18512 8279 18564 8288
rect 18512 8245 18521 8279
rect 18521 8245 18555 8279
rect 18555 8245 18564 8279
rect 18512 8236 18564 8245
rect 18696 8279 18748 8288
rect 18696 8245 18705 8279
rect 18705 8245 18739 8279
rect 18739 8245 18748 8279
rect 18696 8236 18748 8245
rect 18972 8347 19024 8356
rect 18972 8313 18981 8347
rect 18981 8313 19015 8347
rect 19015 8313 19024 8347
rect 18972 8304 19024 8313
rect 19156 8304 19208 8356
rect 19984 8440 20036 8492
rect 19708 8372 19760 8424
rect 22468 8508 22520 8560
rect 24492 8576 24544 8628
rect 25320 8576 25372 8628
rect 25780 8576 25832 8628
rect 23664 8508 23716 8560
rect 23848 8508 23900 8560
rect 21088 8372 21140 8424
rect 22744 8415 22796 8424
rect 22744 8381 22753 8415
rect 22753 8381 22787 8415
rect 22787 8381 22796 8415
rect 22744 8372 22796 8381
rect 22468 8304 22520 8356
rect 23204 8440 23256 8492
rect 23112 8415 23164 8424
rect 23112 8381 23121 8415
rect 23121 8381 23155 8415
rect 23155 8381 23164 8415
rect 23112 8372 23164 8381
rect 21732 8236 21784 8288
rect 23204 8347 23256 8356
rect 23204 8313 23213 8347
rect 23213 8313 23247 8347
rect 23247 8313 23256 8347
rect 23204 8304 23256 8313
rect 23756 8236 23808 8288
rect 23940 8236 23992 8288
rect 24400 8415 24452 8424
rect 24400 8381 24409 8415
rect 24409 8381 24443 8415
rect 24443 8381 24452 8415
rect 24400 8372 24452 8381
rect 25688 8415 25740 8424
rect 25688 8381 25697 8415
rect 25697 8381 25731 8415
rect 25731 8381 25740 8415
rect 25688 8372 25740 8381
rect 25872 8415 25924 8424
rect 25872 8381 25881 8415
rect 25881 8381 25915 8415
rect 25915 8381 25924 8415
rect 25872 8372 25924 8381
rect 25964 8415 26016 8424
rect 25964 8381 25973 8415
rect 25973 8381 26007 8415
rect 26007 8381 26016 8415
rect 25964 8372 26016 8381
rect 27252 8576 27304 8628
rect 27804 8576 27856 8628
rect 30196 8576 30248 8628
rect 27620 8508 27672 8560
rect 26884 8415 26936 8424
rect 26884 8381 26893 8415
rect 26893 8381 26927 8415
rect 26927 8381 26936 8415
rect 26884 8372 26936 8381
rect 26148 8236 26200 8288
rect 26792 8279 26844 8288
rect 26792 8245 26801 8279
rect 26801 8245 26835 8279
rect 26835 8245 26844 8279
rect 26792 8236 26844 8245
rect 26884 8236 26936 8288
rect 27068 8372 27120 8424
rect 27160 8372 27212 8424
rect 27896 8415 27948 8424
rect 27896 8381 27905 8415
rect 27905 8381 27939 8415
rect 27939 8381 27948 8415
rect 27896 8372 27948 8381
rect 29000 8415 29052 8424
rect 29000 8381 29009 8415
rect 29009 8381 29043 8415
rect 29043 8381 29052 8415
rect 29000 8372 29052 8381
rect 27068 8236 27120 8288
rect 27160 8279 27212 8288
rect 27160 8245 27169 8279
rect 27169 8245 27203 8279
rect 27203 8245 27212 8279
rect 27160 8236 27212 8245
rect 27252 8236 27304 8288
rect 27620 8236 27672 8288
rect 27804 8236 27856 8288
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 5908 8032 5960 8084
rect 7012 8032 7064 8084
rect 7932 8032 7984 8084
rect 6644 7896 6696 7948
rect 6736 7939 6788 7948
rect 6736 7905 6745 7939
rect 6745 7905 6779 7939
rect 6779 7905 6788 7939
rect 6736 7896 6788 7905
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 7748 7896 7800 7948
rect 7012 7828 7064 7880
rect 9680 8032 9732 8084
rect 10048 7964 10100 8016
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 11060 8032 11112 8084
rect 10692 7964 10744 8016
rect 11520 8032 11572 8084
rect 6552 7760 6604 7812
rect 9680 7828 9732 7880
rect 10508 7828 10560 7880
rect 11336 7896 11388 7948
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 12532 7964 12584 8016
rect 13544 8032 13596 8084
rect 13636 8032 13688 8084
rect 14280 8032 14332 8084
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 16488 8032 16540 8084
rect 16764 8032 16816 8084
rect 13820 8007 13872 8016
rect 13820 7973 13829 8007
rect 13829 7973 13863 8007
rect 13863 7973 13872 8007
rect 13820 7964 13872 7973
rect 15108 7964 15160 8016
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 13636 7939 13688 7948
rect 13636 7905 13640 7939
rect 13640 7905 13674 7939
rect 13674 7905 13688 7939
rect 13636 7896 13688 7905
rect 13176 7828 13228 7880
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 16580 7896 16632 7948
rect 11152 7760 11204 7812
rect 5448 7692 5500 7744
rect 6184 7692 6236 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 13544 7692 13596 7744
rect 15292 7828 15344 7880
rect 16120 7828 16172 7880
rect 17684 8075 17736 8084
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 18420 8032 18472 8084
rect 19248 8032 19300 8084
rect 17040 7964 17092 8016
rect 19432 8032 19484 8084
rect 22744 8032 22796 8084
rect 23204 8032 23256 8084
rect 25688 8075 25740 8084
rect 25688 8041 25697 8075
rect 25697 8041 25731 8075
rect 25731 8041 25740 8075
rect 25688 8032 25740 8041
rect 25964 8032 26016 8084
rect 17132 7896 17184 7948
rect 17684 7896 17736 7948
rect 17868 7939 17920 7948
rect 17868 7905 17877 7939
rect 17877 7905 17911 7939
rect 17911 7905 17920 7939
rect 17868 7896 17920 7905
rect 18236 7896 18288 7948
rect 19524 7896 19576 7948
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 18420 7828 18472 7880
rect 20076 7896 20128 7948
rect 16212 7692 16264 7744
rect 22652 7871 22704 7880
rect 22652 7837 22661 7871
rect 22661 7837 22695 7871
rect 22695 7837 22704 7871
rect 22652 7828 22704 7837
rect 23020 7896 23072 7948
rect 23296 7828 23348 7880
rect 23848 7896 23900 7948
rect 24032 7939 24084 7948
rect 24032 7905 24041 7939
rect 24041 7905 24075 7939
rect 24075 7905 24084 7939
rect 24032 7896 24084 7905
rect 24124 7896 24176 7948
rect 26792 7964 26844 8016
rect 24400 7896 24452 7948
rect 26884 7896 26936 7948
rect 27160 7896 27212 7948
rect 27252 7939 27304 7948
rect 27252 7905 27261 7939
rect 27261 7905 27295 7939
rect 27295 7905 27304 7939
rect 27252 7896 27304 7905
rect 27804 7964 27856 8016
rect 30380 7964 30432 8016
rect 26148 7828 26200 7880
rect 27988 7939 28040 7948
rect 27988 7905 27997 7939
rect 27997 7905 28031 7939
rect 28031 7905 28040 7939
rect 27988 7896 28040 7905
rect 28080 7939 28132 7948
rect 28080 7905 28089 7939
rect 28089 7905 28123 7939
rect 28123 7905 28132 7939
rect 28080 7896 28132 7905
rect 28172 7896 28224 7948
rect 29736 7939 29788 7948
rect 29736 7905 29745 7939
rect 29745 7905 29779 7939
rect 29779 7905 29788 7939
rect 29736 7896 29788 7905
rect 30012 7896 30064 7948
rect 18880 7692 18932 7744
rect 20628 7735 20680 7744
rect 20628 7701 20637 7735
rect 20637 7701 20671 7735
rect 20671 7701 20680 7735
rect 20628 7692 20680 7701
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 23756 7735 23808 7744
rect 23756 7701 23765 7735
rect 23765 7701 23799 7735
rect 23799 7701 23808 7735
rect 23756 7692 23808 7701
rect 24032 7692 24084 7744
rect 24952 7692 25004 7744
rect 26240 7760 26292 7812
rect 27528 7803 27580 7812
rect 27528 7769 27537 7803
rect 27537 7769 27571 7803
rect 27571 7769 27580 7803
rect 27528 7760 27580 7769
rect 27160 7692 27212 7744
rect 27988 7803 28040 7812
rect 27988 7769 27997 7803
rect 27997 7769 28031 7803
rect 28031 7769 28040 7803
rect 27988 7760 28040 7769
rect 30748 7939 30800 7948
rect 30748 7905 30757 7939
rect 30757 7905 30791 7939
rect 30791 7905 30800 7939
rect 30748 7896 30800 7905
rect 31024 7871 31076 7880
rect 31024 7837 31033 7871
rect 31033 7837 31067 7871
rect 31067 7837 31076 7871
rect 31024 7828 31076 7837
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 6184 7488 6236 7540
rect 6736 7488 6788 7540
rect 6828 7488 6880 7540
rect 7656 7488 7708 7540
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 10416 7531 10468 7540
rect 10416 7497 10425 7531
rect 10425 7497 10459 7531
rect 10459 7497 10468 7531
rect 10416 7488 10468 7497
rect 10508 7531 10560 7540
rect 10508 7497 10517 7531
rect 10517 7497 10551 7531
rect 10551 7497 10560 7531
rect 10508 7488 10560 7497
rect 11428 7488 11480 7540
rect 15016 7488 15068 7540
rect 16120 7488 16172 7540
rect 16580 7488 16632 7540
rect 17316 7488 17368 7540
rect 17868 7488 17920 7540
rect 20628 7488 20680 7540
rect 21272 7488 21324 7540
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 4068 7352 4120 7404
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 7012 7420 7064 7472
rect 4252 7216 4304 7268
rect 6552 7216 6604 7268
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 9864 7420 9916 7472
rect 7656 7284 7708 7336
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 8208 7284 8260 7336
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9956 7284 10008 7336
rect 11612 7352 11664 7404
rect 10600 7284 10652 7336
rect 7380 7216 7432 7268
rect 10048 7259 10100 7268
rect 10048 7225 10057 7259
rect 10057 7225 10091 7259
rect 10091 7225 10100 7259
rect 10048 7216 10100 7225
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 11244 7284 11296 7336
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 13636 7327 13688 7336
rect 13636 7293 13646 7327
rect 13646 7293 13680 7327
rect 13680 7293 13688 7327
rect 13636 7284 13688 7293
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 14004 7327 14056 7336
rect 14004 7293 14018 7327
rect 14018 7293 14052 7327
rect 14052 7293 14056 7327
rect 14004 7284 14056 7293
rect 14464 7284 14516 7336
rect 14832 7327 14884 7336
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 17684 7420 17736 7472
rect 20536 7420 20588 7472
rect 16764 7327 16816 7336
rect 16764 7293 16773 7327
rect 16773 7293 16807 7327
rect 16807 7293 16816 7327
rect 16764 7284 16816 7293
rect 17316 7327 17368 7336
rect 8484 7148 8536 7200
rect 9036 7148 9088 7200
rect 13728 7148 13780 7200
rect 14004 7148 14056 7200
rect 14372 7148 14424 7200
rect 16212 7148 16264 7200
rect 16580 7148 16632 7200
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 17132 7259 17184 7268
rect 17132 7225 17141 7259
rect 17141 7225 17175 7259
rect 17175 7225 17184 7259
rect 17132 7216 17184 7225
rect 17684 7327 17736 7336
rect 17684 7293 17693 7327
rect 17693 7293 17727 7327
rect 17727 7293 17736 7327
rect 17684 7284 17736 7293
rect 17776 7327 17828 7336
rect 17776 7293 17785 7327
rect 17785 7293 17819 7327
rect 17819 7293 17828 7327
rect 17776 7284 17828 7293
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 18788 7352 18840 7404
rect 19984 7284 20036 7336
rect 23848 7463 23900 7472
rect 23848 7429 23857 7463
rect 23857 7429 23891 7463
rect 23891 7429 23900 7463
rect 23848 7420 23900 7429
rect 24400 7531 24452 7540
rect 24400 7497 24409 7531
rect 24409 7497 24443 7531
rect 24443 7497 24452 7531
rect 24400 7488 24452 7497
rect 25872 7488 25924 7540
rect 28172 7488 28224 7540
rect 30380 7531 30432 7540
rect 30380 7497 30389 7531
rect 30389 7497 30423 7531
rect 30423 7497 30432 7531
rect 30380 7488 30432 7497
rect 21456 7327 21508 7336
rect 21456 7293 21463 7327
rect 21463 7293 21508 7327
rect 21456 7284 21508 7293
rect 21732 7327 21784 7336
rect 21732 7293 21746 7327
rect 21746 7293 21780 7327
rect 21780 7293 21784 7327
rect 21732 7284 21784 7293
rect 20720 7216 20772 7268
rect 23756 7352 23808 7404
rect 23112 7284 23164 7336
rect 26056 7420 26108 7472
rect 24032 7352 24084 7404
rect 17592 7148 17644 7200
rect 18788 7191 18840 7200
rect 18788 7157 18797 7191
rect 18797 7157 18831 7191
rect 18831 7157 18840 7191
rect 18788 7148 18840 7157
rect 23940 7216 23992 7268
rect 24952 7327 25004 7336
rect 24952 7293 24961 7327
rect 24961 7293 24995 7327
rect 24995 7293 25004 7327
rect 24952 7284 25004 7293
rect 25044 7327 25096 7336
rect 25044 7293 25054 7327
rect 25054 7293 25088 7327
rect 25088 7293 25096 7327
rect 25044 7284 25096 7293
rect 29000 7395 29052 7404
rect 29000 7361 29009 7395
rect 29009 7361 29043 7395
rect 29043 7361 29052 7395
rect 29000 7352 29052 7361
rect 24860 7148 24912 7200
rect 25320 7259 25372 7268
rect 25320 7225 25329 7259
rect 25329 7225 25363 7259
rect 25363 7225 25372 7259
rect 25320 7216 25372 7225
rect 26240 7327 26292 7336
rect 26240 7293 26249 7327
rect 26249 7293 26283 7327
rect 26283 7293 26292 7327
rect 26240 7284 26292 7293
rect 26424 7284 26476 7336
rect 26976 7284 27028 7336
rect 27160 7284 27212 7336
rect 27988 7284 28040 7336
rect 26608 7216 26660 7268
rect 27252 7216 27304 7268
rect 27712 7259 27764 7268
rect 27712 7225 27721 7259
rect 27721 7225 27755 7259
rect 27755 7225 27764 7259
rect 27712 7216 27764 7225
rect 26148 7191 26200 7200
rect 26148 7157 26157 7191
rect 26157 7157 26191 7191
rect 26191 7157 26200 7191
rect 26148 7148 26200 7157
rect 26792 7191 26844 7200
rect 26792 7157 26801 7191
rect 26801 7157 26835 7191
rect 26835 7157 26844 7191
rect 26792 7148 26844 7157
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 4252 6987 4304 6996
rect 4252 6953 4261 6987
rect 4261 6953 4295 6987
rect 4295 6953 4304 6987
rect 4252 6944 4304 6953
rect 6828 6944 6880 6996
rect 7380 6944 7432 6996
rect 5448 6876 5500 6928
rect 5908 6808 5960 6860
rect 6920 6808 6972 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 11336 6944 11388 6996
rect 8024 6808 8076 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 11612 6808 11664 6860
rect 11704 6851 11756 6860
rect 11704 6817 11713 6851
rect 11713 6817 11747 6851
rect 11747 6817 11756 6851
rect 11704 6808 11756 6817
rect 7380 6672 7432 6724
rect 9864 6740 9916 6792
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 8668 6672 8720 6724
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 6552 6604 6604 6656
rect 6828 6604 6880 6656
rect 10324 6604 10376 6656
rect 11060 6604 11112 6656
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 11888 6604 11940 6656
rect 12900 6604 12952 6656
rect 13544 6851 13596 6860
rect 13544 6817 13578 6851
rect 13578 6817 13596 6851
rect 13544 6808 13596 6817
rect 14464 6944 14516 6996
rect 16580 6944 16632 6996
rect 17132 6944 17184 6996
rect 17684 6944 17736 6996
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 19340 6944 19392 6996
rect 19524 6944 19576 6996
rect 14648 6808 14700 6860
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 13268 6672 13320 6724
rect 15292 6740 15344 6792
rect 17592 6808 17644 6860
rect 18788 6876 18840 6928
rect 23296 6944 23348 6996
rect 25320 6944 25372 6996
rect 26884 6944 26936 6996
rect 18144 6851 18196 6860
rect 18144 6817 18153 6851
rect 18153 6817 18187 6851
rect 18187 6817 18196 6851
rect 18144 6808 18196 6817
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 18052 6740 18104 6792
rect 19984 6808 20036 6860
rect 20628 6851 20680 6860
rect 20628 6817 20635 6851
rect 20635 6817 20680 6851
rect 20628 6808 20680 6817
rect 20720 6851 20772 6860
rect 20720 6817 20729 6851
rect 20729 6817 20763 6851
rect 20763 6817 20772 6851
rect 20720 6808 20772 6817
rect 20812 6851 20864 6860
rect 20812 6817 20821 6851
rect 20821 6817 20855 6851
rect 20855 6817 20864 6851
rect 20812 6808 20864 6817
rect 20904 6851 20956 6860
rect 20904 6817 20918 6851
rect 20918 6817 20952 6851
rect 20952 6817 20956 6851
rect 20904 6808 20956 6817
rect 23204 6851 23256 6860
rect 14740 6604 14792 6656
rect 15108 6647 15160 6656
rect 15108 6613 15117 6647
rect 15117 6613 15151 6647
rect 15151 6613 15160 6647
rect 15108 6604 15160 6613
rect 17776 6604 17828 6656
rect 21732 6783 21784 6792
rect 21732 6749 21741 6783
rect 21741 6749 21775 6783
rect 21775 6749 21784 6783
rect 21732 6740 21784 6749
rect 18604 6604 18656 6656
rect 19064 6604 19116 6656
rect 20352 6604 20404 6656
rect 23204 6817 23213 6851
rect 23213 6817 23247 6851
rect 23247 6817 23256 6851
rect 23204 6808 23256 6817
rect 23940 6808 23992 6860
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 24124 6808 24176 6860
rect 26148 6876 26200 6928
rect 22284 6740 22336 6792
rect 22744 6783 22796 6792
rect 22744 6749 22753 6783
rect 22753 6749 22787 6783
rect 22787 6749 22796 6783
rect 22744 6740 22796 6749
rect 22928 6715 22980 6724
rect 22928 6681 22937 6715
rect 22937 6681 22971 6715
rect 22971 6681 22980 6715
rect 22928 6672 22980 6681
rect 23480 6783 23532 6792
rect 23480 6749 23489 6783
rect 23489 6749 23523 6783
rect 23523 6749 23532 6783
rect 23480 6740 23532 6749
rect 26792 6808 26844 6860
rect 27252 6876 27304 6928
rect 27160 6851 27212 6860
rect 27160 6817 27169 6851
rect 27169 6817 27203 6851
rect 27203 6817 27212 6851
rect 27160 6808 27212 6817
rect 26424 6740 26476 6792
rect 28080 6808 28132 6860
rect 28724 6851 28776 6860
rect 28724 6817 28733 6851
rect 28733 6817 28767 6851
rect 28767 6817 28776 6851
rect 28724 6808 28776 6817
rect 30012 6876 30064 6928
rect 29092 6851 29144 6860
rect 29092 6817 29101 6851
rect 29101 6817 29135 6851
rect 29135 6817 29144 6851
rect 29092 6808 29144 6817
rect 29736 6808 29788 6860
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 29368 6715 29420 6724
rect 29368 6681 29377 6715
rect 29377 6681 29411 6715
rect 29411 6681 29420 6715
rect 29368 6672 29420 6681
rect 27160 6604 27212 6656
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 5448 6196 5500 6248
rect 5816 6196 5868 6248
rect 3608 6171 3660 6180
rect 3608 6137 3617 6171
rect 3617 6137 3651 6171
rect 3651 6137 3660 6171
rect 3608 6128 3660 6137
rect 5908 6128 5960 6180
rect 6000 6171 6052 6180
rect 6000 6137 6009 6171
rect 6009 6137 6043 6171
rect 6043 6137 6052 6171
rect 6000 6128 6052 6137
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 9864 6400 9916 6452
rect 11796 6400 11848 6452
rect 13084 6400 13136 6452
rect 13544 6443 13596 6452
rect 13544 6409 13553 6443
rect 13553 6409 13587 6443
rect 13587 6409 13596 6443
rect 13544 6400 13596 6409
rect 12900 6332 12952 6384
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 11060 6239 11112 6248
rect 11060 6205 11094 6239
rect 11094 6205 11112 6239
rect 3516 6060 3568 6112
rect 5724 6060 5776 6112
rect 8576 6060 8628 6112
rect 11060 6196 11112 6205
rect 11520 6196 11572 6248
rect 12992 6264 13044 6316
rect 12716 6196 12768 6248
rect 14004 6264 14056 6316
rect 15200 6375 15252 6384
rect 15200 6341 15209 6375
rect 15209 6341 15243 6375
rect 15243 6341 15252 6375
rect 15200 6332 15252 6341
rect 16396 6400 16448 6452
rect 16764 6400 16816 6452
rect 17592 6400 17644 6452
rect 18604 6400 18656 6452
rect 20812 6400 20864 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 24124 6400 24176 6452
rect 25228 6400 25280 6452
rect 25964 6400 26016 6452
rect 27252 6400 27304 6452
rect 28724 6400 28776 6452
rect 15108 6264 15160 6316
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 14096 6128 14148 6180
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 14740 6239 14792 6248
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 15292 6239 15344 6248
rect 15292 6205 15301 6239
rect 15301 6205 15335 6239
rect 15335 6205 15344 6239
rect 15292 6196 15344 6205
rect 17684 6264 17736 6316
rect 15200 6128 15252 6180
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 14648 6060 14700 6112
rect 18144 6060 18196 6112
rect 19156 6060 19208 6112
rect 20352 6239 20404 6248
rect 20352 6205 20386 6239
rect 20386 6205 20404 6239
rect 20352 6196 20404 6205
rect 20720 6196 20772 6248
rect 22928 6239 22980 6248
rect 22928 6205 22937 6239
rect 22937 6205 22971 6239
rect 22971 6205 22980 6239
rect 22928 6196 22980 6205
rect 23848 6239 23900 6248
rect 23848 6205 23857 6239
rect 23857 6205 23891 6239
rect 23891 6205 23900 6239
rect 23848 6196 23900 6205
rect 24124 6239 24176 6248
rect 24124 6205 24133 6239
rect 24133 6205 24167 6239
rect 24167 6205 24176 6239
rect 24124 6196 24176 6205
rect 24860 6264 24912 6316
rect 25964 6239 26016 6248
rect 25964 6205 25973 6239
rect 25973 6205 26007 6239
rect 26007 6205 26016 6239
rect 25964 6196 26016 6205
rect 23112 6103 23164 6112
rect 23112 6069 23121 6103
rect 23121 6069 23155 6103
rect 23155 6069 23164 6103
rect 23112 6060 23164 6069
rect 24400 6171 24452 6180
rect 24400 6137 24409 6171
rect 24409 6137 24443 6171
rect 24443 6137 24452 6171
rect 24400 6128 24452 6137
rect 26240 6239 26292 6248
rect 26240 6205 26249 6239
rect 26249 6205 26283 6239
rect 26283 6205 26292 6239
rect 26240 6196 26292 6205
rect 26976 6196 27028 6248
rect 27160 6239 27212 6248
rect 27160 6205 27169 6239
rect 27169 6205 27203 6239
rect 27203 6205 27212 6239
rect 27160 6196 27212 6205
rect 26516 6171 26568 6180
rect 26516 6137 26525 6171
rect 26525 6137 26559 6171
rect 26559 6137 26568 6171
rect 26516 6128 26568 6137
rect 26700 6060 26752 6112
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 5816 5856 5868 5908
rect 5908 5856 5960 5908
rect 8576 5856 8628 5908
rect 10140 5856 10192 5908
rect 2780 5720 2832 5772
rect 3516 5763 3568 5772
rect 3516 5729 3525 5763
rect 3525 5729 3559 5763
rect 3559 5729 3568 5763
rect 3516 5720 3568 5729
rect 10324 5856 10376 5908
rect 11704 5856 11756 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 5724 5516 5776 5568
rect 10968 5720 11020 5772
rect 13636 5720 13688 5772
rect 14096 5720 14148 5772
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 6644 5652 6696 5704
rect 10232 5652 10284 5704
rect 14280 5652 14332 5704
rect 17592 5856 17644 5908
rect 17868 5856 17920 5908
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 20628 5856 20680 5908
rect 23112 5856 23164 5908
rect 24124 5856 24176 5908
rect 24400 5856 24452 5908
rect 26516 5856 26568 5908
rect 16764 5720 16816 5772
rect 16948 5720 17000 5772
rect 18696 5788 18748 5840
rect 19156 5788 19208 5840
rect 18604 5720 18656 5772
rect 19340 5720 19392 5772
rect 22100 5763 22152 5772
rect 22100 5729 22123 5763
rect 22123 5729 22152 5763
rect 22100 5720 22152 5729
rect 11520 5516 11572 5568
rect 13268 5516 13320 5568
rect 14832 5584 14884 5636
rect 15292 5584 15344 5636
rect 16488 5652 16540 5704
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 15016 5516 15068 5568
rect 15660 5516 15712 5568
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 29092 5856 29144 5908
rect 23388 5720 23440 5772
rect 23940 5720 23992 5772
rect 24032 5720 24084 5772
rect 26424 5720 26476 5772
rect 26700 5720 26752 5772
rect 27344 5763 27396 5772
rect 27344 5729 27353 5763
rect 27353 5729 27387 5763
rect 27387 5729 27396 5763
rect 27344 5720 27396 5729
rect 29000 5720 29052 5772
rect 26608 5516 26660 5568
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 5908 5312 5960 5364
rect 6828 5312 6880 5364
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 4068 5176 4120 5228
rect 6092 5244 6144 5296
rect 6644 5244 6696 5296
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 7288 5176 7340 5228
rect 5724 5108 5776 5160
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 3608 5083 3660 5092
rect 3608 5049 3617 5083
rect 3617 5049 3651 5083
rect 3651 5049 3660 5083
rect 3608 5040 3660 5049
rect 4344 5040 4396 5092
rect 6092 5151 6144 5160
rect 6092 5117 6101 5151
rect 6101 5117 6135 5151
rect 6135 5117 6144 5151
rect 6092 5108 6144 5117
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 7840 5312 7892 5364
rect 8944 5312 8996 5364
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 12716 5312 12768 5364
rect 13176 5355 13228 5364
rect 13176 5321 13185 5355
rect 13185 5321 13219 5355
rect 13219 5321 13228 5355
rect 13176 5312 13228 5321
rect 11520 5176 11572 5228
rect 16212 5244 16264 5296
rect 16488 5355 16540 5364
rect 16488 5321 16497 5355
rect 16497 5321 16531 5355
rect 16531 5321 16540 5355
rect 16488 5312 16540 5321
rect 16948 5312 17000 5364
rect 19340 5312 19392 5364
rect 20076 5355 20128 5364
rect 20076 5321 20085 5355
rect 20085 5321 20119 5355
rect 20119 5321 20128 5355
rect 20076 5312 20128 5321
rect 21456 5312 21508 5364
rect 9864 5040 9916 5092
rect 10692 5040 10744 5092
rect 13912 5040 13964 5092
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 17960 5151 18012 5160
rect 17960 5117 17969 5151
rect 17969 5117 18003 5151
rect 18003 5117 18012 5151
rect 17960 5108 18012 5117
rect 18696 5151 18748 5160
rect 18696 5117 18705 5151
rect 18705 5117 18739 5151
rect 18739 5117 18748 5151
rect 27252 5312 27304 5364
rect 27712 5355 27764 5364
rect 27712 5321 27721 5355
rect 27721 5321 27755 5355
rect 27755 5321 27764 5355
rect 27712 5312 27764 5321
rect 18696 5108 18748 5117
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 5816 4972 5868 5024
rect 5908 5015 5960 5024
rect 5908 4981 5917 5015
rect 5917 4981 5951 5015
rect 5951 4981 5960 5015
rect 5908 4972 5960 4981
rect 7104 4972 7156 5024
rect 7932 4972 7984 5024
rect 8760 4972 8812 5024
rect 9404 4972 9456 5024
rect 9680 4972 9732 5024
rect 13268 4972 13320 5024
rect 14280 5015 14332 5024
rect 14280 4981 14289 5015
rect 14289 4981 14323 5015
rect 14323 4981 14332 5015
rect 14280 4972 14332 4981
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 14740 4972 14792 5024
rect 18420 5040 18472 5092
rect 15660 4972 15712 5024
rect 16580 4972 16632 5024
rect 17960 4972 18012 5024
rect 20536 4972 20588 5024
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 3608 4768 3660 4820
rect 4344 4768 4396 4820
rect 5356 4768 5408 4820
rect 5908 4768 5960 4820
rect 6828 4768 6880 4820
rect 7104 4700 7156 4752
rect 7288 4768 7340 4820
rect 12716 4768 12768 4820
rect 13268 4768 13320 4820
rect 13728 4768 13780 4820
rect 7932 4700 7984 4752
rect 5448 4564 5500 4616
rect 6460 4564 6512 4616
rect 10692 4700 10744 4752
rect 12348 4700 12400 4752
rect 14556 4768 14608 4820
rect 14740 4768 14792 4820
rect 18420 4811 18472 4820
rect 9036 4675 9088 4684
rect 9036 4641 9045 4675
rect 9045 4641 9079 4675
rect 9079 4641 9088 4675
rect 9036 4632 9088 4641
rect 9404 4675 9456 4684
rect 9404 4641 9413 4675
rect 9413 4641 9447 4675
rect 9447 4641 9456 4675
rect 9404 4632 9456 4641
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 11060 4632 11112 4684
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 11520 4632 11572 4684
rect 12440 4675 12492 4684
rect 12440 4641 12474 4675
rect 12474 4641 12492 4675
rect 13912 4743 13964 4752
rect 13912 4709 13921 4743
rect 13921 4709 13955 4743
rect 13955 4709 13964 4743
rect 13912 4700 13964 4709
rect 14556 4675 14608 4684
rect 12440 4632 12492 4641
rect 14556 4641 14565 4675
rect 14565 4641 14599 4675
rect 14599 4641 14608 4675
rect 14556 4632 14608 4641
rect 15108 4632 15160 4684
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 20536 4768 20588 4820
rect 9864 4564 9916 4616
rect 10784 4539 10836 4548
rect 10784 4505 10793 4539
rect 10793 4505 10827 4539
rect 10827 4505 10836 4539
rect 10784 4496 10836 4505
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 14464 4496 14516 4548
rect 15108 4496 15160 4548
rect 17960 4700 18012 4752
rect 19524 4700 19576 4752
rect 20444 4700 20496 4752
rect 25044 4768 25096 4820
rect 18604 4675 18656 4684
rect 18604 4641 18613 4675
rect 18613 4641 18647 4675
rect 18647 4641 18656 4675
rect 18604 4632 18656 4641
rect 21456 4675 21508 4684
rect 21456 4641 21465 4675
rect 21465 4641 21499 4675
rect 21499 4641 21508 4675
rect 21456 4632 21508 4641
rect 23388 4700 23440 4752
rect 16580 4564 16632 4616
rect 20812 4564 20864 4616
rect 20996 4539 21048 4548
rect 20996 4505 21005 4539
rect 21005 4505 21039 4539
rect 21039 4505 21048 4539
rect 22652 4632 22704 4684
rect 20996 4496 21048 4505
rect 22192 4496 22244 4548
rect 23572 4632 23624 4684
rect 12532 4428 12584 4480
rect 20628 4428 20680 4480
rect 21456 4428 21508 4480
rect 21916 4428 21968 4480
rect 22468 4428 22520 4480
rect 22560 4471 22612 4480
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 22560 4428 22612 4437
rect 22928 4471 22980 4480
rect 22928 4437 22937 4471
rect 22937 4437 22971 4471
rect 22971 4437 22980 4471
rect 22928 4428 22980 4437
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 8760 4224 8812 4276
rect 4068 4156 4120 4208
rect 11152 4224 11204 4276
rect 7104 4088 7156 4140
rect 7748 4020 7800 4072
rect 11060 4156 11112 4208
rect 8944 4020 8996 4072
rect 9036 3952 9088 4004
rect 9680 4020 9732 4072
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 10784 4088 10836 4140
rect 11336 4224 11388 4276
rect 12532 4224 12584 4276
rect 14096 4224 14148 4276
rect 14556 4224 14608 4276
rect 10508 4020 10560 4072
rect 11244 4020 11296 4072
rect 11612 4088 11664 4140
rect 11336 3952 11388 4004
rect 12348 4020 12400 4072
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 19524 4224 19576 4276
rect 15108 4156 15160 4208
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 15844 4088 15896 4140
rect 18236 4156 18288 4208
rect 18604 4156 18656 4208
rect 20812 4224 20864 4276
rect 23388 4224 23440 4276
rect 16212 4020 16264 4072
rect 16488 4063 16540 4072
rect 16488 4029 16497 4063
rect 16497 4029 16531 4063
rect 16531 4029 16540 4063
rect 16488 4020 16540 4029
rect 19340 4020 19392 4072
rect 20536 4020 20588 4072
rect 20628 4063 20680 4072
rect 20628 4029 20637 4063
rect 20637 4029 20671 4063
rect 20671 4029 20680 4063
rect 20628 4020 20680 4029
rect 22560 4088 22612 4140
rect 23572 4088 23624 4140
rect 20996 4020 21048 4072
rect 11060 3927 11112 3936
rect 11060 3893 11069 3927
rect 11069 3893 11103 3927
rect 11103 3893 11112 3927
rect 11244 3927 11296 3936
rect 11060 3884 11112 3893
rect 11244 3893 11271 3927
rect 11271 3893 11296 3927
rect 11244 3884 11296 3893
rect 12532 3884 12584 3936
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 22100 3952 22152 4004
rect 22928 3952 22980 4004
rect 23848 3952 23900 4004
rect 18236 3884 18288 3893
rect 18972 3884 19024 3936
rect 20444 3884 20496 3936
rect 21088 3884 21140 3936
rect 26240 3927 26292 3936
rect 26240 3893 26249 3927
rect 26249 3893 26283 3927
rect 26283 3893 26292 3927
rect 26240 3884 26292 3893
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 9680 3680 9732 3732
rect 11612 3680 11664 3732
rect 12440 3680 12492 3732
rect 13728 3680 13780 3732
rect 15568 3680 15620 3732
rect 21456 3680 21508 3732
rect 23940 3680 23992 3732
rect 9128 3612 9180 3664
rect 7748 3544 7800 3596
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 11060 3544 11112 3596
rect 11244 3544 11296 3596
rect 11520 3612 11572 3664
rect 12256 3612 12308 3664
rect 12532 3544 12584 3596
rect 12716 3544 12768 3596
rect 13912 3612 13964 3664
rect 16764 3612 16816 3664
rect 14924 3544 14976 3596
rect 15660 3544 15712 3596
rect 12348 3476 12400 3528
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 10140 3340 10192 3392
rect 11336 3340 11388 3392
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 13728 3476 13780 3528
rect 18420 3544 18472 3596
rect 20076 3612 20128 3664
rect 21088 3655 21140 3664
rect 21088 3621 21097 3655
rect 21097 3621 21131 3655
rect 21131 3621 21140 3655
rect 21088 3612 21140 3621
rect 18972 3544 19024 3596
rect 14648 3408 14700 3460
rect 16488 3476 16540 3528
rect 21824 3519 21876 3528
rect 21824 3485 21833 3519
rect 21833 3485 21867 3519
rect 21867 3485 21876 3519
rect 21824 3476 21876 3485
rect 22192 3476 22244 3528
rect 16212 3340 16264 3392
rect 16948 3340 17000 3392
rect 21916 3340 21968 3392
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 8116 3068 8168 3120
rect 12716 3179 12768 3188
rect 12716 3145 12725 3179
rect 12725 3145 12759 3179
rect 12759 3145 12768 3179
rect 12716 3136 12768 3145
rect 16488 3136 16540 3188
rect 20076 3136 20128 3188
rect 21824 3136 21876 3188
rect 23848 3136 23900 3188
rect 18420 3111 18472 3120
rect 18420 3077 18429 3111
rect 18429 3077 18463 3111
rect 18463 3077 18472 3111
rect 18420 3068 18472 3077
rect 11612 3000 11664 3052
rect 16212 3000 16264 3052
rect 21456 3000 21508 3052
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 14924 2932 14976 2984
rect 19340 2932 19392 2984
rect 16948 2907 17000 2916
rect 16948 2873 16957 2907
rect 16957 2873 16991 2907
rect 16991 2873 17000 2907
rect 16948 2864 17000 2873
rect 21088 2932 21140 2984
rect 22192 2864 22244 2916
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 16304 960 16356 1012
rect 16396 1003 16448 1012
rect 16396 969 16405 1003
rect 16405 969 16439 1003
rect 16439 969 16448 1003
rect 16396 960 16448 969
rect 16856 1003 16908 1012
rect 16856 969 16865 1003
rect 16865 969 16899 1003
rect 16899 969 16908 1003
rect 16856 960 16908 969
rect 6552 799 6604 808
rect 6552 765 6561 799
rect 6561 765 6595 799
rect 6595 765 6604 799
rect 6552 756 6604 765
rect 14280 799 14332 808
rect 14280 765 14289 799
rect 14289 765 14323 799
rect 14323 765 14332 799
rect 14280 756 14332 765
rect 15568 799 15620 808
rect 15568 765 15577 799
rect 15577 765 15611 799
rect 15611 765 15620 799
rect 15568 756 15620 765
rect 16212 799 16264 808
rect 16212 765 16221 799
rect 16221 765 16255 799
rect 16255 765 16264 799
rect 16212 756 16264 765
rect 16764 756 16816 808
rect 18788 799 18840 808
rect 18788 765 18797 799
rect 18797 765 18831 799
rect 18831 765 18840 799
rect 18788 756 18840 765
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
<< metal2 >>
rect 10322 19600 10378 20000
rect 10966 19600 11022 20000
rect 11610 19600 11666 20000
rect 12254 19600 12310 20000
rect 12898 19600 12954 20000
rect 15474 19600 15530 20000
rect 16118 19600 16174 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 19338 19600 19394 20000
rect 19982 19600 20038 20000
rect 20626 19600 20682 20000
rect 21270 19600 21326 20000
rect 21914 19600 21970 20000
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 10336 18834 10364 19600
rect 10980 18834 11008 19600
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 4250 18459 4558 18468
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 11520 16720 11572 16726
rect 11624 16708 11652 19600
rect 12268 18834 12296 19600
rect 12912 18834 12940 19600
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 12624 16720 12676 16726
rect 11624 16680 11744 16708
rect 11520 16662 11572 16668
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6656 15502 6684 16186
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 4250 15260 4558 15269
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 6104 15026 6132 15438
rect 7944 15162 7972 15574
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 848 14476 900 14482
rect 848 14418 900 14424
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 860 14385 888 14418
rect 846 14376 902 14385
rect 846 14311 902 14320
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2424 14006 2452 14282
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2792 13530 2820 13670
rect 2884 13530 2912 13806
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13530 3096 13670
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 848 10600 900 10606
rect 848 10542 900 10548
rect 860 10305 888 10542
rect 846 10296 902 10305
rect 846 10231 902 10240
rect 3160 10198 3188 14418
rect 3252 12782 3280 14894
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 3424 14544 3476 14550
rect 3424 14486 3476 14492
rect 3436 14074 3464 14486
rect 4080 14482 4108 14826
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3712 14074 3740 14350
rect 4724 14346 4752 14758
rect 4816 14618 4844 14826
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4896 14476 4948 14482
rect 6104 14464 6132 14962
rect 8956 14958 8984 16594
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 15978 9168 16390
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9048 15706 9076 15846
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9048 15026 9076 15642
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9140 15094 9168 15506
rect 9600 15502 9628 16594
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9784 16114 9812 16390
rect 10336 16250 10364 16594
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10428 15706 10456 15982
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10888 15570 10916 16050
rect 11440 16046 11468 16390
rect 11532 16182 11560 16662
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11624 16250 11652 16526
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11520 16176 11572 16182
rect 11520 16118 11572 16124
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 9600 15366 9628 15438
rect 10336 15366 10364 15438
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 9128 15088 9180 15094
rect 10140 15088 10192 15094
rect 9128 15030 9180 15036
rect 9968 15048 10140 15076
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 6288 14618 6316 14894
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14618 6408 14758
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6276 14476 6328 14482
rect 6104 14436 6276 14464
rect 4896 14418 4948 14424
rect 6276 14418 6328 14424
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4356 13802 4384 14010
rect 4724 14006 4752 14282
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 4816 13870 4844 14214
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4068 13728 4120 13734
rect 4252 13728 4304 13734
rect 4120 13676 4200 13682
rect 4068 13670 4200 13676
rect 4252 13670 4304 13676
rect 4080 13654 4200 13670
rect 4172 13394 4200 13654
rect 4264 13394 4292 13670
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4066 13288 4122 13297
rect 4066 13223 4068 13232
rect 4120 13223 4122 13232
rect 4068 13194 4120 13200
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3252 11150 3280 12718
rect 3528 12481 3556 13126
rect 4172 12850 4200 13126
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3514 12472 3570 12481
rect 3514 12407 3570 12416
rect 3528 12374 3556 12407
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3620 12102 3648 12582
rect 4172 12442 4200 12650
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4632 12306 4660 12378
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11370 3556 11494
rect 3436 11354 3556 11370
rect 3424 11348 3556 11354
rect 3476 11342 3556 11348
rect 3424 11290 3476 11296
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9466 3188 9862
rect 3252 9654 3280 11086
rect 3528 10606 3556 11342
rect 3804 11286 3832 11698
rect 4080 11694 4108 12174
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 4632 11762 4660 12242
rect 4724 11830 4752 13330
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4816 12306 4844 13126
rect 4908 12306 4936 14418
rect 4988 13864 5040 13870
rect 5040 13812 5120 13818
rect 4988 13806 5120 13812
rect 5000 13790 5120 13806
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5000 12986 5028 13670
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5092 12714 5120 13790
rect 6380 13734 6408 14554
rect 6472 13938 6500 14894
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6656 14618 6684 14758
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6748 14498 6776 14554
rect 6656 14470 6776 14498
rect 6656 14414 6684 14470
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4802 12200 4858 12209
rect 4802 12135 4804 12144
rect 4856 12135 4858 12144
rect 4804 12106 4856 12112
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11354 4016 11494
rect 4632 11354 4660 11698
rect 5092 11642 5120 12650
rect 5276 12442 5304 12718
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5184 12322 5212 12378
rect 5184 12294 5304 12322
rect 5368 12306 5396 13126
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5460 12345 5488 12582
rect 5540 12368 5592 12374
rect 5446 12336 5502 12345
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5184 11898 5212 12174
rect 5276 12170 5304 12294
rect 5356 12300 5408 12306
rect 5644 12356 5672 12582
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5592 12328 5672 12356
rect 5540 12310 5592 12316
rect 5446 12271 5502 12280
rect 5356 12242 5408 12248
rect 5264 12164 5316 12170
rect 5736 12152 5764 12378
rect 5816 12300 5868 12306
rect 5920 12288 5948 12582
rect 6012 12306 6040 12718
rect 6656 12434 6684 13126
rect 6840 12782 6868 13670
rect 6932 13326 6960 14350
rect 7024 14074 7052 14758
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 8956 14618 8984 14894
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7576 14074 7604 14486
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7024 13870 7052 14010
rect 7668 13870 7696 14214
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6932 12714 6960 13262
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 7116 12646 7144 13806
rect 7668 13462 7696 13806
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 8036 13394 8064 13942
rect 9048 13870 9076 14962
rect 9140 14550 9168 15030
rect 9968 14822 9996 15048
rect 10140 15030 10192 15036
rect 10336 14890 10364 15302
rect 10520 15162 10548 15506
rect 11072 15502 11100 15914
rect 11440 15706 11468 15982
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10520 14958 10548 15098
rect 11072 14958 11100 15438
rect 11440 14958 11468 15642
rect 11532 14958 11560 16118
rect 11716 15706 11744 16680
rect 12624 16662 12676 16668
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 12636 16250 12664 16662
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12728 15706 12756 16050
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 11440 14618 11468 14894
rect 11624 14822 11652 15506
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11808 14890 11836 15302
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 6564 12406 6684 12434
rect 6826 12472 6882 12481
rect 6826 12407 6828 12416
rect 6564 12306 6592 12406
rect 6880 12407 6882 12416
rect 6920 12436 6972 12442
rect 6828 12378 6880 12384
rect 6920 12378 6972 12384
rect 5868 12260 5948 12288
rect 6000 12300 6052 12306
rect 5816 12242 5868 12248
rect 6000 12242 6052 12248
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 5816 12164 5868 12170
rect 5736 12124 5816 12152
rect 5264 12106 5316 12112
rect 5816 12106 5868 12112
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5092 11626 5304 11642
rect 4988 11620 5040 11626
rect 5092 11620 5316 11626
rect 5092 11614 5264 11620
rect 4988 11562 5040 11568
rect 5264 11562 5316 11568
rect 5000 11354 5028 11562
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 5184 10606 5212 10950
rect 5276 10674 5304 11562
rect 6012 11354 6040 12242
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6104 11898 6132 12174
rect 6656 12102 6684 12242
rect 6932 12170 6960 12378
rect 7012 12300 7064 12306
rect 7116 12288 7144 12582
rect 7484 12442 7512 12650
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7064 12260 7144 12288
rect 7012 12242 7064 12248
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6656 11830 6684 12038
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5000 10266 5028 10406
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5276 10130 5304 10610
rect 5920 10606 5948 10950
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6748 10198 6776 11494
rect 7116 11354 7144 12260
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7300 11665 7328 12242
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7576 11898 7604 12174
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7668 11694 7696 12718
rect 7760 11830 7788 12718
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12306 7880 12582
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 8680 12434 8708 13262
rect 8772 12986 8800 13330
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 8680 12406 8892 12434
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 8036 11694 8064 12242
rect 8680 11898 8708 12242
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 7656 11688 7708 11694
rect 7286 11656 7342 11665
rect 7656 11630 7708 11636
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7286 11591 7342 11600
rect 7564 11620 7616 11626
rect 7300 11354 7328 11591
rect 7564 11562 7616 11568
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7576 11218 7604 11562
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7668 10554 7696 11494
rect 7760 11354 7788 11630
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7760 11234 7788 11290
rect 7760 11206 7880 11234
rect 7760 10674 7788 11206
rect 7852 11150 7880 11206
rect 7944 11150 7972 11494
rect 8036 11257 8064 11630
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8022 11248 8078 11257
rect 8312 11218 8340 11290
rect 8208 11212 8260 11218
rect 8022 11183 8078 11192
rect 8128 11172 8208 11200
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7932 11144 7984 11150
rect 8128 11121 8156 11172
rect 8208 11154 8260 11160
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 7932 11086 7984 11092
rect 8114 11112 8170 11121
rect 8114 11047 8170 11056
rect 8484 11076 8536 11082
rect 8588 11064 8616 11766
rect 8666 11656 8722 11665
rect 8666 11591 8722 11600
rect 8680 11218 8708 11591
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8536 11036 8616 11064
rect 8484 11018 8536 11024
rect 8680 11014 8708 11154
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 8116 11008 8168 11014
rect 8300 11008 8352 11014
rect 8168 10968 8300 10996
rect 8116 10950 8168 10956
rect 8300 10950 8352 10956
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 7944 10674 7972 10950
rect 8772 10674 8800 11154
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 7840 10600 7892 10606
rect 7668 10548 7840 10554
rect 7668 10542 7892 10548
rect 7668 10526 7880 10542
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 7944 10130 7972 10406
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 8102 10299 8410 10308
rect 8496 10130 8524 10474
rect 8864 10198 8892 12406
rect 9692 12374 9720 12582
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9232 11286 9260 11766
rect 9600 11694 9628 12038
rect 9692 11694 9720 12038
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 11354 9444 11562
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9220 11280 9272 11286
rect 9126 11248 9182 11257
rect 9048 11218 9126 11234
rect 9036 11212 9126 11218
rect 9088 11206 9126 11212
rect 9220 11222 9272 11228
rect 9126 11183 9182 11192
rect 9036 11154 9088 11160
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 5644 9518 5672 9862
rect 3240 9512 3292 9518
rect 3160 9460 3240 9466
rect 3160 9454 3292 9460
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 3160 9438 3280 9454
rect 3252 9042 3280 9438
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8430 4108 8910
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 4816 8634 4844 9318
rect 6012 9178 6040 9318
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 7116 9110 7144 9454
rect 7208 9110 7236 10066
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9178 7328 9318
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8634 5028 8978
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5736 8634 5764 8842
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 7012 8560 7064 8566
rect 6380 8498 6960 8514
rect 7012 8502 7064 8508
rect 6368 8492 6960 8498
rect 6420 8486 6960 8492
rect 6368 8434 6420 8440
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 5778 2820 7346
rect 3252 7342 3280 8230
rect 4080 7410 4108 8366
rect 5920 8090 5948 8366
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 6656 7954 6684 8366
rect 6932 8362 6960 8486
rect 6736 8356 6788 8362
rect 6920 8356 6972 8362
rect 6788 8316 6868 8344
rect 6736 8298 6788 8304
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3252 6236 3280 7278
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4264 7002 4292 7210
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 5460 6934 5488 7686
rect 6196 7546 6224 7686
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6458 7304 6514 7313
rect 6564 7274 6592 7754
rect 6748 7546 6776 7890
rect 6840 7546 6868 8316
rect 6920 8298 6972 8304
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6458 7239 6514 7248
rect 6552 7268 6604 7274
rect 6472 7206 6500 7239
rect 6552 7210 6604 7216
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 5460 6254 5488 6870
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 3332 6248 3384 6254
rect 3252 6208 3332 6236
rect 3332 6190 3384 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 3344 5234 3372 6190
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5778 3556 6054
rect 3620 5914 3648 6122
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3620 4826 3648 5034
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 4080 4214 4108 5170
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4356 4826 4384 5034
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4826 5396 4966
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5460 4622 5488 6190
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5574 5764 6054
rect 5828 5914 5856 6190
rect 5920 6186 5948 6802
rect 6564 6662 6592 7210
rect 6840 7002 6868 7278
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6932 6866 6960 8298
rect 7024 8090 7052 8502
rect 7116 8498 7144 9046
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7208 8634 7236 8774
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7300 8514 7328 8774
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7208 8486 7328 8514
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7116 7954 7144 8434
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7478 7052 7822
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6254 6868 6598
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5920 5914 5948 6122
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 5166 5764 5510
rect 5920 5370 5948 5850
rect 6012 5710 6040 6122
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5724 5160 5776 5166
rect 5908 5160 5960 5166
rect 5724 5102 5776 5108
rect 5828 5108 5908 5114
rect 6012 5148 6040 5646
rect 6656 5302 6684 5646
rect 6840 5370 6868 6190
rect 7208 5681 7236 8486
rect 7378 8392 7434 8401
rect 7378 8327 7380 8336
rect 7432 8327 7434 8336
rect 7380 8298 7432 8304
rect 7944 8090 7972 8774
rect 8864 8498 8892 10134
rect 9036 8628 9088 8634
rect 9140 8616 9168 11183
rect 9232 11121 9260 11222
rect 9404 11144 9456 11150
rect 9218 11112 9274 11121
rect 9692 11098 9720 11494
rect 9456 11092 9720 11098
rect 9404 11086 9720 11092
rect 9416 11070 9720 11086
rect 9218 11047 9274 11056
rect 9784 10198 9812 14214
rect 9876 13870 9904 14214
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9876 13394 9904 13806
rect 10782 13560 10838 13569
rect 10600 13524 10652 13530
rect 11256 13546 11284 14350
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11256 13518 11468 13546
rect 10782 13495 10838 13504
rect 10600 13466 10652 13472
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 12374 9904 13330
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9876 11558 9904 12310
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9232 9518 9260 10066
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9382 9260 9454
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9088 8588 9168 8616
rect 9036 8570 9088 8576
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 8496 8004 8524 8434
rect 8404 7976 8524 8004
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7546 7788 7890
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7668 7342 7696 7482
rect 8404 7342 8432 7976
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 8024 7336 8076 7342
rect 8208 7336 8260 7342
rect 8024 7278 8076 7284
rect 8206 7304 8208 7313
rect 8392 7336 8444 7342
rect 8260 7304 8262 7313
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7392 7002 7420 7210
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7392 6730 7420 6938
rect 8036 6866 8064 7278
rect 8444 7284 8800 7290
rect 8392 7278 8800 7284
rect 8404 7262 8800 7278
rect 8206 7239 8262 7248
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 8496 6866 8524 7142
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7194 5672 7250 5681
rect 7194 5607 7250 5616
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6104 5166 6132 5238
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 5960 5120 6040 5148
rect 6092 5160 6144 5166
rect 5828 5102 5960 5108
rect 6092 5102 6144 5108
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 5828 5086 5948 5102
rect 5828 5030 5856 5086
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4826 5948 4966
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6472 4622 6500 5102
rect 6840 4826 6868 5170
rect 7208 5166 7236 5607
rect 7852 5370 7880 6802
rect 8680 6730 8708 6802
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8772 6322 8800 7262
rect 9048 7206 9076 8570
rect 9416 8430 9444 8774
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9692 8090 9720 10134
rect 10152 10130 10180 10746
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 9876 9722 9904 10066
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9784 9382 9812 9658
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 8588 5914 8616 6054
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 7116 4758 7144 4966
rect 7300 4826 7328 5170
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7944 4758 7972 4966
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 7116 4146 7144 4694
rect 8772 4282 8800 4966
rect 8956 4672 8984 5306
rect 9692 5030 9720 7822
rect 9876 7478 9904 9658
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 10060 9518 10088 9551
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 10140 9036 10192 9042
rect 10244 9024 10272 10066
rect 10336 9674 10364 13398
rect 10612 13190 10640 13466
rect 10796 13394 10824 13495
rect 11440 13433 11468 13518
rect 11426 13424 11482 13433
rect 10784 13388 10836 13394
rect 11244 13388 11296 13394
rect 10836 13348 11192 13376
rect 10784 13330 10836 13336
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12782 10732 13126
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10704 11558 10732 12038
rect 10796 11762 10824 12038
rect 11060 11824 11112 11830
rect 11058 11792 11060 11801
rect 11112 11792 11114 11801
rect 10784 11756 10836 11762
rect 11058 11727 11114 11736
rect 10784 11698 10836 11704
rect 11060 11688 11112 11694
rect 11058 11656 11060 11665
rect 11112 11656 11114 11665
rect 11058 11591 11114 11600
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 11354 10732 11494
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10612 10810 10640 11154
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10130 10640 10406
rect 10704 10198 10732 10678
rect 10796 10606 10824 10950
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10600 10124 10652 10130
rect 10520 10084 10600 10112
rect 10336 9646 10456 9674
rect 10428 9110 10456 9646
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10192 8996 10272 9024
rect 10140 8978 10192 8984
rect 9968 8430 9996 8978
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 10048 8288 10100 8294
rect 9954 8256 10010 8265
rect 10048 8230 10100 8236
rect 9954 8191 10010 8200
rect 9968 7954 9996 8191
rect 10060 8022 10088 8230
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10152 7834 10180 8978
rect 10428 8498 10456 9046
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10060 7806 10180 7834
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 6458 9904 6734
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9968 5370 9996 7278
rect 10060 7274 10088 7806
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5914 10180 6054
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10244 5817 10272 8434
rect 10520 8265 10548 10084
rect 10600 10066 10652 10072
rect 10876 9988 10928 9994
rect 10876 9930 10928 9936
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10506 8256 10562 8265
rect 10506 8191 10562 8200
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7546 10456 7686
rect 10520 7546 10548 7822
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10612 7342 10640 9590
rect 10888 9586 10916 9930
rect 11072 9602 11100 11591
rect 11164 11098 11192 13348
rect 11426 13359 11482 13368
rect 11244 13330 11296 13336
rect 11256 12442 11284 13330
rect 11440 12594 11468 13359
rect 11532 12782 11560 13670
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11624 12918 11652 13330
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11716 12782 11744 12922
rect 12360 12850 12388 13126
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11704 12776 11756 12782
rect 12072 12776 12124 12782
rect 11704 12718 11756 12724
rect 12070 12744 12072 12753
rect 12440 12776 12492 12782
rect 12124 12744 12126 12753
rect 12126 12702 12388 12730
rect 12440 12718 12492 12724
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12070 12679 12126 12688
rect 12072 12640 12124 12646
rect 11440 12566 11652 12594
rect 12072 12582 12124 12588
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11532 12102 11560 12310
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11256 11218 11284 11766
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11164 11070 11284 11098
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10980 9574 11100 9602
rect 10980 9382 11008 9574
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10704 8022 10732 8366
rect 11072 8090 11100 9454
rect 11164 9110 11192 10542
rect 11256 9110 11284 11070
rect 11348 9654 11376 11562
rect 11426 11248 11482 11257
rect 11426 11183 11428 11192
rect 11480 11183 11482 11192
rect 11428 11154 11480 11160
rect 11532 11014 11560 12038
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11440 10606 11468 10950
rect 11532 10674 11560 10950
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11532 10130 11560 10474
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11348 9382 11376 9590
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11244 9104 11296 9110
rect 11348 9081 11376 9114
rect 11244 9046 11296 9052
rect 11334 9072 11390 9081
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 8430 11192 8570
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 11164 7818 11192 8230
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11256 7342 11284 9046
rect 11334 9007 11390 9016
rect 11532 8838 11560 9454
rect 11624 9110 11652 12566
rect 12084 12374 12112 12582
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11348 7954 11376 8366
rect 11532 8090 11560 8774
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 5914 10364 6598
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10230 5808 10286 5817
rect 10980 5778 11008 7278
rect 11348 7002 11376 7890
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11440 7546 11468 7822
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6254 11100 6598
rect 11532 6254 11560 8026
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 6866 11652 7346
rect 11716 7018 11744 12174
rect 11808 11898 11836 12242
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11900 11694 11928 11834
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11808 11354 11836 11562
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 11354 12112 11494
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11955 10843 12263 10852
rect 12360 10198 12388 12702
rect 12452 12170 12480 12718
rect 12544 12442 12572 12718
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12636 12374 12664 15642
rect 12820 15434 12848 15982
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12820 14482 12848 15370
rect 13556 14822 13584 15914
rect 14660 15706 14688 15914
rect 14924 15904 14976 15910
rect 15028 15892 15056 16118
rect 14976 15864 15056 15892
rect 14924 15846 14976 15852
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13740 14958 13768 15370
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13372 14618 13400 14758
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 14936 14482 14964 14962
rect 15028 14618 15056 15864
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12728 13462 12756 14214
rect 13280 14074 13308 14350
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12728 12986 12756 13262
rect 12912 13258 12940 13738
rect 13726 13424 13782 13433
rect 13648 13394 13726 13410
rect 13636 13388 13726 13394
rect 13688 13382 13726 13388
rect 13726 13359 13782 13368
rect 13636 13330 13688 13336
rect 13542 13288 13598 13297
rect 12900 13252 12952 13258
rect 13542 13223 13598 13232
rect 12900 13194 12952 13200
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12624 12368 12676 12374
rect 12624 12310 12676 12316
rect 12820 12306 12848 12854
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12452 11694 12480 12106
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12622 11792 12678 11801
rect 12532 11756 12584 11762
rect 12622 11727 12678 11736
rect 12532 11698 12584 11704
rect 12440 11688 12492 11694
rect 12544 11665 12572 11698
rect 12636 11694 12664 11727
rect 12624 11688 12676 11694
rect 12440 11630 12492 11636
rect 12530 11656 12586 11665
rect 12728 11665 12756 11834
rect 12624 11630 12676 11636
rect 12714 11656 12770 11665
rect 12530 11591 12586 11600
rect 12714 11591 12770 11600
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12452 11218 12480 11494
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12728 9926 12756 11591
rect 12820 11257 12848 12106
rect 12912 11744 12940 13194
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13004 11914 13032 13126
rect 13096 12986 13124 13126
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13096 12170 13124 12718
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12374 13216 12582
rect 13280 12442 13308 12718
rect 13556 12646 13584 13223
rect 13728 12776 13780 12782
rect 13924 12730 13952 14010
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13728 12718 13780 12724
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13740 12442 13768 12718
rect 13832 12702 13952 12730
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13280 12170 13308 12378
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13556 11937 13584 12174
rect 13542 11928 13598 11937
rect 13004 11886 13124 11914
rect 12992 11756 13044 11762
rect 12912 11716 12992 11744
rect 12992 11698 13044 11704
rect 12806 11248 12862 11257
rect 12806 11183 12862 11192
rect 13096 10713 13124 11886
rect 13542 11863 13598 11872
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13188 11354 13216 11698
rect 13832 11694 13860 12702
rect 14016 12442 14044 12922
rect 14108 12646 14136 13330
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 13025 14688 13126
rect 14646 13016 14702 13025
rect 14646 12951 14702 12960
rect 14660 12730 14688 12951
rect 14568 12702 14688 12730
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 13832 11354 13860 11494
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13372 11121 13400 11154
rect 13358 11112 13414 11121
rect 13358 11047 13414 11056
rect 13818 11112 13874 11121
rect 13818 11047 13874 11056
rect 13082 10704 13138 10713
rect 13082 10639 13138 10648
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12268 8906 12296 9386
rect 12912 9382 12940 9522
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12806 9072 12862 9081
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12532 9036 12584 9042
rect 13004 9042 13032 10134
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13096 9110 13124 9318
rect 13648 9160 13676 9318
rect 13464 9132 13676 9160
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13266 9072 13322 9081
rect 12806 9007 12808 9016
rect 12532 8978 12584 8984
rect 12860 9007 12862 9016
rect 12992 9036 13044 9042
rect 12808 8978 12860 8984
rect 13266 9007 13268 9016
rect 12992 8978 13044 8984
rect 13320 9007 13322 9016
rect 13268 8978 13320 8984
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12084 8362 12112 8502
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12176 8294 12204 8502
rect 12360 8498 12388 8978
rect 12438 8664 12494 8673
rect 12438 8599 12494 8608
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12452 8294 12480 8599
rect 12544 8430 12572 8978
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12544 8022 12572 8230
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11808 7857 11836 7890
rect 11794 7848 11850 7857
rect 11794 7783 11850 7792
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 11716 6990 11836 7018
rect 11808 6882 11836 6990
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11704 6860 11756 6866
rect 11808 6854 11928 6882
rect 11704 6802 11756 6808
rect 11716 6769 11744 6802
rect 11796 6792 11848 6798
rect 11702 6760 11758 6769
rect 11796 6734 11848 6740
rect 11702 6695 11758 6704
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 10230 5743 10286 5752
rect 10968 5772 11020 5778
rect 10244 5710 10272 5743
rect 10968 5714 11020 5720
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 11532 5574 11560 6190
rect 11716 5914 11744 6598
rect 11808 6458 11836 6734
rect 11900 6662 11928 6854
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11955 6491 12263 6500
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 11532 5234 11560 5510
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 12728 5370 12756 6190
rect 12820 5914 12848 8298
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 6390 12940 6598
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 13004 6322 13032 8978
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6458 13124 6734
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13188 5370 13216 7822
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13280 5574 13308 6666
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9416 4690 9444 4966
rect 9036 4684 9088 4690
rect 8956 4644 9036 4672
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 8956 4078 8984 4644
rect 9036 4626 9088 4632
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9876 4622 9904 5034
rect 10704 4758 10732 5034
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 11532 4690 11560 5170
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4826 13308 4966
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 7760 3602 7788 4014
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 8128 3126 8156 3538
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 9048 2990 9076 3946
rect 9692 3738 9720 4014
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9140 3194 9168 3606
rect 9876 3398 9904 4558
rect 9968 4078 9996 4626
rect 10520 4078 10548 4626
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4146 10824 4490
rect 11072 4214 11100 4626
rect 11164 4282 11192 4626
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11060 4208 11112 4214
rect 11060 4154 11112 4156
rect 11060 4150 11192 4154
rect 10784 4140 10836 4146
rect 11072 4126 11192 4150
rect 10784 4082 10836 4088
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 11060 3936 11112 3942
rect 11164 3924 11192 4126
rect 11256 4078 11284 4422
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11348 4154 11376 4218
rect 11348 4126 11560 4154
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11244 3936 11296 3942
rect 11164 3896 11244 3924
rect 11060 3878 11112 3884
rect 11244 3878 11296 3884
rect 11072 3602 11100 3878
rect 11256 3602 11284 3878
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10152 3398 10180 3538
rect 11348 3398 11376 3946
rect 11532 3670 11560 4126
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11624 3738 11652 4082
rect 12360 4078 12388 4694
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12452 4162 12480 4626
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4282 12572 4422
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12452 4134 12572 4162
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12268 3505 12296 3606
rect 12360 3534 12388 4014
rect 12452 3738 12480 4014
rect 12544 3942 12572 4134
rect 12728 4078 12756 4762
rect 13464 4154 13492 9132
rect 13832 9042 13860 11047
rect 14292 10674 14320 11494
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 10198 14044 10542
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 14016 9722 14044 10134
rect 14004 9716 14056 9722
rect 14200 9674 14228 10202
rect 14292 10130 14320 10406
rect 14568 10266 14596 12702
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14660 12374 14688 12582
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14752 10606 14780 13670
rect 14844 12374 14872 14214
rect 15028 13870 15056 14554
rect 15120 14482 15148 16594
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15396 15638 15424 16186
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15396 15094 15424 15574
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15396 14906 15424 15030
rect 15212 14890 15424 14906
rect 15200 14884 15424 14890
rect 15252 14878 15424 14884
rect 15200 14826 15252 14832
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15120 14278 15148 14418
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14936 10606 14964 13126
rect 15212 11218 15240 14282
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 13938 15332 14214
rect 15396 14074 15424 14878
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15382 13560 15438 13569
rect 15382 13495 15438 13504
rect 15396 13394 15424 13495
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15396 11914 15424 13330
rect 15488 12288 15516 19600
rect 16132 19258 16160 19600
rect 16132 19230 16252 19258
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 16224 18834 16252 19230
rect 18064 18834 18092 19600
rect 18708 18834 18736 19600
rect 19352 18834 19380 19600
rect 19996 18834 20024 19600
rect 20640 18834 20668 19600
rect 21284 18834 21312 19600
rect 21928 18834 21956 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 31217 19068 31525 19077
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 31036 18465 31064 18566
rect 31022 18456 31078 18465
rect 31022 18391 31078 18400
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18248 16114 18276 16730
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 15672 15706 15700 16050
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15672 14890 15700 15506
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15948 14822 15976 15098
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15580 14550 15608 14758
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 16224 14618 16252 14894
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 15568 14544 15620 14550
rect 16132 14521 16160 14554
rect 15568 14486 15620 14492
rect 16118 14512 16174 14521
rect 16316 14498 16344 14962
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14521 16620 14758
rect 16776 14550 16804 14894
rect 17144 14618 17172 14962
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16764 14544 16816 14550
rect 16224 14482 16344 14498
rect 16578 14512 16634 14521
rect 16118 14447 16174 14456
rect 16212 14476 16344 14482
rect 16264 14470 16344 14476
rect 16488 14476 16540 14482
rect 16212 14418 16264 14424
rect 16764 14486 16816 14492
rect 17236 14482 17264 16050
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17972 15434 18000 15982
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17498 15056 17554 15065
rect 17498 14991 17554 15000
rect 17512 14958 17540 14991
rect 18156 14958 18184 15302
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 16578 14447 16634 14456
rect 17224 14476 17276 14482
rect 16488 14418 16540 14424
rect 17224 14418 17276 14424
rect 16500 14006 16528 14418
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 15672 13802 15792 13818
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15672 13796 15804 13802
rect 15672 13790 15752 13796
rect 15580 13530 15608 13738
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15580 13326 15608 13466
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15672 13258 15700 13790
rect 15752 13738 15804 13744
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 17512 13433 17540 14894
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17604 14550 17632 14758
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17498 13424 17554 13433
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16488 13388 16540 13394
rect 17498 13359 17554 13368
rect 16488 13330 16540 13336
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15856 12918 15884 13330
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 15672 12714 15884 12730
rect 15672 12708 15896 12714
rect 15672 12702 15844 12708
rect 15672 12434 15700 12702
rect 15844 12650 15896 12656
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 16224 12442 16252 12786
rect 16316 12782 16344 13330
rect 16500 12986 16528 13330
rect 17314 13288 17370 13297
rect 17314 13223 17370 13232
rect 17328 13190 17356 13223
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16304 12776 16356 12782
rect 16356 12736 16436 12764
rect 16304 12718 16356 12724
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12442 16344 12582
rect 16212 12436 16264 12442
rect 15672 12406 15792 12434
rect 15488 12260 15700 12288
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15304 11886 15424 11914
rect 15304 11393 15332 11886
rect 15488 11694 15516 12038
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15290 11384 15346 11393
rect 15290 11319 15346 11328
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15120 11014 15148 11154
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15304 10554 15332 11154
rect 15396 10674 15424 11494
rect 15488 11082 15516 11494
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15304 10538 15424 10554
rect 15304 10532 15436 10538
rect 15304 10526 15384 10532
rect 15384 10474 15436 10480
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14004 9658 14056 9664
rect 14016 9194 14044 9658
rect 13924 9166 14044 9194
rect 14108 9646 14228 9674
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13556 8090 13584 8978
rect 13740 8634 13768 8978
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13648 7954 13676 8026
rect 13832 8022 13860 8842
rect 13924 8430 13952 9166
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13924 7970 13952 8366
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7342 13584 7686
rect 13832 7342 13860 7958
rect 13924 7942 14044 7970
rect 14016 7342 14044 7942
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14004 7336 14056 7342
rect 14108 7313 14136 9646
rect 14292 8090 14320 10066
rect 14660 9518 14688 10406
rect 15396 10266 15424 10474
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14568 9178 14596 9454
rect 14752 9382 14780 10066
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14752 9042 14780 9318
rect 15028 9042 15056 9998
rect 15488 9518 15516 10406
rect 15580 10266 15608 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15672 9654 15700 12260
rect 15764 12209 15792 12406
rect 16212 12378 16264 12384
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 15842 12336 15898 12345
rect 16316 12306 16344 12378
rect 16408 12306 16436 12736
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16592 12306 16620 12650
rect 16776 12594 16804 12650
rect 16776 12566 16988 12594
rect 15842 12271 15844 12280
rect 15896 12271 15898 12280
rect 16304 12300 16356 12306
rect 15844 12242 15896 12248
rect 16304 12242 16356 12248
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 15750 12200 15806 12209
rect 15750 12135 15806 12144
rect 16408 11694 16436 12242
rect 15844 11688 15896 11694
rect 15750 11656 15806 11665
rect 15806 11636 15844 11642
rect 15806 11630 15896 11636
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 15806 11614 15884 11630
rect 15750 11591 15806 11600
rect 15807 11452 16115 11461
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15807 11387 16115 11396
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 10810 15792 10950
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16132 10674 16160 11290
rect 16408 11286 16436 11630
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 15807 10364 16115 10373
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 16224 10130 16252 10406
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14384 8430 14412 8978
rect 15028 8838 15056 8978
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14004 7278 14056 7284
rect 14094 7304 14150 7313
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13556 6458 13584 6802
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13648 5778 13676 7278
rect 14094 7239 14150 7248
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13740 4826 13768 7142
rect 14016 6322 14044 7142
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14108 6186 14136 7239
rect 14384 7206 14412 8366
rect 15120 8022 15148 9114
rect 15396 8090 15424 9454
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15488 8566 15516 8978
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15856 8430 15884 9046
rect 16224 9042 16252 9930
rect 16316 9674 16344 11222
rect 16500 11014 16528 11222
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10266 16436 10406
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16408 9674 16436 9862
rect 16316 9646 16436 9674
rect 16302 9072 16358 9081
rect 16212 9036 16264 9042
rect 16302 9007 16358 9016
rect 16212 8978 16264 8984
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15807 8123 16115 8132
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15028 7546 15056 7890
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16224 7834 16252 8978
rect 16316 7954 16344 9007
rect 16408 8294 16436 9646
rect 16592 9518 16620 9862
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16500 8430 16528 9114
rect 16684 9081 16712 9114
rect 16670 9072 16726 9081
rect 16670 9007 16726 9016
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16500 8090 16528 8366
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14476 7002 14504 7278
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14660 6254 14688 6802
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6254 14780 6598
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14660 6118 14688 6190
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13924 4758 13952 5034
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 13464 4126 13584 4154
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 3602 12572 3878
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12348 3528 12400 3534
rect 12254 3496 12310 3505
rect 12348 3470 12400 3476
rect 12254 3431 12310 3440
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 11624 3058 11652 3334
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 12728 3194 12756 3538
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 6552 808 6604 814
rect 6552 750 6604 756
rect 6564 490 6592 750
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 6472 462 6592 490
rect 6472 400 6500 462
rect 13556 400 13584 4126
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13740 3534 13768 3674
rect 13924 3670 13952 4694
rect 14108 4282 14136 5714
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14292 5030 14320 5646
rect 14844 5642 14872 7278
rect 15014 6896 15070 6905
rect 15014 6831 15016 6840
rect 15068 6831 15070 6840
rect 15016 6802 15068 6808
rect 15304 6798 15332 7822
rect 16132 7546 16160 7822
rect 16224 7806 16344 7834
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16224 7206 16252 7686
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15120 6322 15148 6598
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15212 6186 15240 6326
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 5681 15148 5714
rect 15106 5672 15162 5681
rect 14832 5636 14884 5642
rect 15304 5642 15332 6190
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 15106 5607 15162 5616
rect 15292 5636 15344 5642
rect 14832 5578 14884 5584
rect 15292 5578 15344 5584
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4554 14504 4966
rect 14568 4826 14596 5510
rect 15028 5234 15056 5510
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 15672 5030 15700 5510
rect 16224 5302 16252 5510
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 14752 4826 14780 4966
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14568 4282 14596 4626
rect 15120 4554 15148 4626
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 15120 4214 15148 4490
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15844 4140 15896 4146
rect 15672 4100 15844 4128
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15580 3738 15608 4014
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 15672 3602 15700 4100
rect 15844 4082 15896 4088
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 14646 3496 14702 3505
rect 14646 3431 14648 3440
rect 14700 3431 14702 3440
rect 14648 3402 14700 3408
rect 14936 2990 14964 3538
rect 16224 3398 16252 4014
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16224 3058 16252 3334
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 16316 1018 16344 7806
rect 16408 6458 16436 7890
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16500 6338 16528 8026
rect 16592 7954 16620 8230
rect 16776 8090 16804 9318
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 8430 16896 8774
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16578 7848 16634 7857
rect 16578 7783 16634 7792
rect 16592 7546 16620 7783
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16592 7002 16620 7142
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16776 6458 16804 7278
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16408 6310 16528 6338
rect 16408 1018 16436 6310
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16500 5370 16528 5646
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4622 16620 4966
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16592 4196 16620 4558
rect 16500 4168 16620 4196
rect 16500 4078 16528 4168
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16776 3670 16804 5714
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16500 3194 16528 3470
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16868 1018 16896 8366
rect 16960 7834 16988 12566
rect 17052 12306 17080 12854
rect 17144 12782 17172 13126
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17604 11540 17632 14486
rect 18156 13802 18184 14894
rect 18340 14521 18368 15846
rect 18984 15706 19012 15914
rect 19168 15910 19196 16526
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 19168 15570 19196 15846
rect 19444 15706 19472 15914
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 20272 15570 20300 15846
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18432 14550 18460 14758
rect 18420 14544 18472 14550
rect 18326 14512 18382 14521
rect 18420 14486 18472 14492
rect 18326 14447 18382 14456
rect 18340 13802 18368 14447
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 14074 18736 14214
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18708 13870 18736 14010
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18800 13512 18828 14894
rect 19168 14890 19196 15506
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 20088 15094 20116 15506
rect 20548 15502 20576 15846
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 19892 14952 19944 14958
rect 20272 14906 20300 15030
rect 19944 14900 20300 14906
rect 19892 14894 20300 14900
rect 19156 14884 19208 14890
rect 19904 14878 20300 14894
rect 19156 14826 19208 14832
rect 20272 14822 20300 14878
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 20260 14816 20312 14822
rect 20364 14804 20392 15302
rect 20548 15162 20576 15438
rect 20640 15162 20668 15506
rect 20824 15366 20852 15506
rect 20916 15502 20944 15914
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 21008 15162 21036 15506
rect 21468 15434 21496 16050
rect 21560 15978 21588 16390
rect 22480 16114 22508 16526
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 21548 15972 21600 15978
rect 21548 15914 21600 15920
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20456 15042 20484 15098
rect 20456 15014 20760 15042
rect 21468 15026 21496 15370
rect 20732 14890 20760 15014
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20444 14816 20496 14822
rect 20364 14776 20444 14804
rect 20260 14758 20312 14764
rect 20444 14758 20496 14764
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18708 13484 18828 13512
rect 18708 13394 18736 13484
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18142 13016 18198 13025
rect 18800 12986 18828 13330
rect 18142 12951 18198 12960
rect 18788 12980 18840 12986
rect 18156 12918 18184 12951
rect 18788 12922 18840 12928
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 17868 12708 17920 12714
rect 17868 12650 17920 12656
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 17880 12442 17908 12650
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11694 17908 12174
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17972 11812 18000 12106
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18144 11824 18196 11830
rect 17972 11784 18144 11812
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17684 11552 17736 11558
rect 17604 11512 17684 11540
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17236 11121 17264 11154
rect 17222 11112 17278 11121
rect 17222 11047 17278 11056
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17512 9178 17540 9454
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17052 8673 17080 9046
rect 17038 8664 17094 8673
rect 17038 8599 17094 8608
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17052 8022 17080 8502
rect 17144 8498 17172 9114
rect 17604 9042 17632 11512
rect 17684 11494 17736 11500
rect 17972 11218 18000 11784
rect 18144 11766 18196 11772
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 18064 11354 18092 11562
rect 18156 11354 18184 11630
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 18248 10810 18276 11834
rect 18432 11150 18460 12650
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18524 11898 18552 12174
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18708 11676 18736 12242
rect 18880 12232 18932 12238
rect 18878 12200 18880 12209
rect 18932 12200 18934 12209
rect 18878 12135 18934 12144
rect 18880 11688 18932 11694
rect 18708 11648 18880 11676
rect 18984 11665 19012 13330
rect 19076 12714 19104 14010
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19168 12753 19196 13330
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12986 19380 13126
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19154 12744 19210 12753
rect 19064 12708 19116 12714
rect 19154 12679 19210 12688
rect 19064 12650 19116 12656
rect 19444 12306 19472 14758
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 20272 13802 20300 14758
rect 22480 14482 22508 16050
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22848 15638 22876 15846
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 22652 14884 22704 14890
rect 22652 14826 22704 14832
rect 22664 14618 22692 14826
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 23308 14482 23336 15370
rect 23676 15065 23704 15506
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 23662 15056 23718 15065
rect 23662 14991 23718 15000
rect 24136 14958 24164 15302
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 23860 14550 23888 14758
rect 23848 14544 23900 14550
rect 23848 14486 23900 14492
rect 23952 14482 23980 14894
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23216 14278 23244 14418
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20088 13546 20116 13670
rect 20088 13518 20300 13546
rect 20272 13394 20300 13518
rect 20352 13456 20404 13462
rect 20444 13456 20496 13462
rect 20404 13424 20444 13444
rect 20496 13424 20498 13433
rect 20404 13416 20442 13424
rect 20352 13398 20404 13404
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20260 13388 20312 13394
rect 20548 13394 20576 13670
rect 20640 13394 20668 13670
rect 23216 13462 23244 14214
rect 23308 13802 23336 14418
rect 25056 13870 25084 14758
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 26240 14272 26292 14278
rect 26240 14214 26292 14220
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 24400 13796 24452 13802
rect 24400 13738 24452 13744
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 20442 13359 20498 13368
rect 20536 13388 20588 13394
rect 20260 13330 20312 13336
rect 20536 13330 20588 13336
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19536 12918 19564 13126
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 20180 12434 20208 13330
rect 20640 13190 20668 13330
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20732 12753 20760 13262
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20824 12986 20852 13126
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20718 12744 20774 12753
rect 20718 12679 20774 12688
rect 20996 12708 21048 12714
rect 19996 12406 20208 12434
rect 19890 12336 19946 12345
rect 19432 12300 19484 12306
rect 19890 12271 19946 12280
rect 19432 12242 19484 12248
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19154 11928 19210 11937
rect 19154 11863 19156 11872
rect 19208 11863 19210 11872
rect 19156 11834 19208 11840
rect 19260 11694 19288 12038
rect 19444 11694 19472 12242
rect 19904 12238 19932 12271
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11830 19564 12038
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19248 11688 19300 11694
rect 18880 11630 18932 11636
rect 18970 11656 19026 11665
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18248 10062 18276 10746
rect 18432 10538 18460 11086
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10606 18828 10950
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18892 10418 18920 11630
rect 19248 11630 19300 11636
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 18970 11591 19026 11600
rect 19536 11354 19564 11766
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19904 11121 19932 11630
rect 19890 11112 19946 11121
rect 19890 11047 19946 11056
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 18800 10390 18920 10418
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18156 9722 18184 9998
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 17696 9178 17724 9386
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17696 8090 17724 8298
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17144 7834 17172 7890
rect 16960 7806 17172 7834
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17328 7342 17356 7482
rect 17696 7478 17724 7890
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17788 7342 17816 8978
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 17880 7546 17908 7890
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17684 7336 17736 7342
rect 17684 7278 17736 7284
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 17144 7002 17172 7210
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17604 6866 17632 7142
rect 17696 7002 17724 7278
rect 17788 7002 17816 7278
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 6458 17632 6802
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17604 5914 17632 6394
rect 17696 6322 17724 6734
rect 17788 6662 17816 6938
rect 18064 6798 18092 7278
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 18156 6118 18184 6802
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18248 5914 18276 7890
rect 18340 7886 18368 8978
rect 18432 8974 18460 9386
rect 18616 9042 18644 9454
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18432 8090 18460 8910
rect 18512 8288 18564 8294
rect 18510 8256 18512 8265
rect 18564 8256 18566 8265
rect 18510 8191 18566 8200
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18432 7886 18460 8026
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18616 6662 18644 8978
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 6769 18736 8230
rect 18800 7410 18828 10390
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18984 9518 19012 9998
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 8974 19012 9454
rect 19168 9450 19196 9998
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 19444 9382 19472 10066
rect 19996 9994 20024 12406
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20088 11898 20116 12242
rect 20272 12102 20300 12242
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20272 11898 20300 12038
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20180 11354 20208 11562
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 11354 20300 11494
rect 20640 11354 20668 12038
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20088 10266 20116 10406
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 20180 9586 20208 11018
rect 20732 10742 20760 12679
rect 20996 12650 21048 12656
rect 20902 12336 20958 12345
rect 20902 12271 20904 12280
rect 20956 12271 20958 12280
rect 20904 12242 20956 12248
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20720 10736 20772 10742
rect 20350 10704 20406 10713
rect 20720 10678 20772 10684
rect 20350 10639 20406 10648
rect 20364 10266 20392 10639
rect 20824 10606 20852 11086
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20916 10266 20944 10406
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20732 9722 20760 10066
rect 20720 9716 20772 9722
rect 21008 9674 21036 12650
rect 21284 12434 21312 13262
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21652 12918 21680 13194
rect 22020 12986 22048 13330
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23124 12986 23152 13126
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 21192 12406 21312 12434
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21100 11898 21128 12242
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21100 11014 21128 11834
rect 21192 11121 21220 12406
rect 21652 12306 21680 12854
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21744 12306 21772 12718
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22940 12594 22968 12854
rect 23020 12844 23072 12850
rect 23072 12804 23152 12832
rect 23020 12786 23072 12792
rect 22388 12374 22416 12582
rect 22940 12566 23060 12594
rect 22376 12368 22428 12374
rect 22376 12310 22428 12316
rect 23032 12306 23060 12566
rect 21364 12300 21416 12306
rect 21284 12260 21364 12288
rect 21284 12102 21312 12260
rect 21364 12242 21416 12248
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22744 12300 22796 12306
rect 23020 12300 23072 12306
rect 22744 12242 22796 12248
rect 22940 12260 23020 12288
rect 21824 12232 21876 12238
rect 21638 12200 21694 12209
rect 21456 12164 21508 12170
rect 21694 12180 21824 12186
rect 21694 12174 21876 12180
rect 21694 12158 21864 12174
rect 21638 12135 21694 12144
rect 21456 12106 21508 12112
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21284 11218 21312 12038
rect 21468 11898 21496 12106
rect 22020 11898 22048 12242
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 21468 11354 21496 11834
rect 22572 11801 22600 12242
rect 22650 11928 22706 11937
rect 22650 11863 22706 11872
rect 22558 11792 22614 11801
rect 22558 11727 22614 11736
rect 22192 11688 22244 11694
rect 21730 11656 21786 11665
rect 22192 11630 22244 11636
rect 21730 11591 21786 11600
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21178 11112 21234 11121
rect 21178 11047 21234 11056
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21192 10266 21220 11047
rect 21744 10606 21772 11591
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21836 10606 21864 11494
rect 22204 11218 22232 11630
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22572 11286 22600 11494
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22664 10996 22692 11863
rect 22756 11830 22784 12242
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 22756 11694 22784 11766
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22848 11558 22876 12038
rect 22940 11762 22968 12260
rect 23020 12242 23072 12248
rect 23124 12288 23152 12804
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23204 12300 23256 12306
rect 23124 12260 23204 12288
rect 23018 11928 23074 11937
rect 23124 11914 23152 12260
rect 23204 12242 23256 12248
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23074 11886 23152 11914
rect 23018 11863 23074 11872
rect 23112 11824 23164 11830
rect 23032 11784 23112 11812
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22940 11354 22968 11698
rect 23032 11626 23060 11784
rect 23112 11766 23164 11772
rect 23216 11694 23244 12038
rect 23308 11898 23336 12718
rect 23400 12434 23428 13126
rect 23492 12986 23520 13330
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 23400 12406 23704 12434
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23492 11898 23520 12038
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23584 11694 23612 12242
rect 23676 12220 23704 12406
rect 23860 12374 23888 12854
rect 23952 12696 23980 13126
rect 24308 12776 24360 12782
rect 24306 12744 24308 12753
rect 24360 12744 24362 12753
rect 24032 12708 24084 12714
rect 23952 12668 24032 12696
rect 23848 12368 23900 12374
rect 23848 12310 23900 12316
rect 23848 12232 23900 12238
rect 23676 12192 23848 12220
rect 23848 12174 23900 12180
rect 23662 11792 23718 11801
rect 23662 11727 23664 11736
rect 23716 11727 23718 11736
rect 23664 11698 23716 11704
rect 23204 11688 23256 11694
rect 23204 11630 23256 11636
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23020 11620 23072 11626
rect 23020 11562 23072 11568
rect 23032 11354 23060 11562
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 22848 11218 22876 11290
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 23860 11150 23888 12174
rect 23952 11665 23980 12668
rect 24306 12679 24362 12688
rect 24032 12650 24084 12656
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24136 11898 24164 12242
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 23938 11656 23994 11665
rect 23938 11591 23994 11600
rect 23020 11144 23072 11150
rect 23664 11144 23716 11150
rect 23072 11092 23152 11098
rect 23020 11086 23152 11092
rect 23664 11086 23716 11092
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23032 11070 23152 11086
rect 23124 11014 23152 11070
rect 23020 11008 23072 11014
rect 22664 10968 22784 10996
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 21732 10600 21784 10606
rect 21732 10542 21784 10548
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 21192 10062 21220 10202
rect 21376 10130 21404 10406
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22204 10146 22232 10202
rect 22296 10198 22324 10746
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 22112 10118 22232 10146
rect 22284 10192 22336 10198
rect 22284 10134 22336 10140
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 20720 9658 20772 9664
rect 20916 9654 21036 9674
rect 20904 9648 21036 9654
rect 20956 9646 21036 9648
rect 20904 9590 20956 9596
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 19984 9444 20036 9450
rect 19812 9404 19984 9432
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18984 8820 19012 8910
rect 19064 8832 19116 8838
rect 18984 8792 19064 8820
rect 19064 8774 19116 8780
rect 19352 8566 19380 9114
rect 19444 9042 19472 9318
rect 19812 9178 19840 9404
rect 19984 9386 20036 9392
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 9178 20668 9318
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19340 8560 19392 8566
rect 18984 8486 19196 8514
rect 19340 8502 19392 8508
rect 18984 8362 19012 8486
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 19076 8265 19104 8366
rect 19168 8362 19196 8486
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19062 8256 19118 8265
rect 19062 8191 19118 8200
rect 19260 8090 19288 8366
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 18880 7744 18932 7750
rect 19352 7698 19380 8366
rect 19444 8090 19472 8978
rect 19616 8832 19668 8838
rect 19536 8792 19616 8820
rect 19536 8498 19564 8792
rect 19616 8774 19668 8780
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19720 8430 19748 8570
rect 19996 8498 20024 9114
rect 20916 9042 20944 9590
rect 21732 9580 21784 9586
rect 21916 9580 21968 9586
rect 21784 9540 21916 9568
rect 21732 9522 21784 9528
rect 21916 9522 21968 9528
rect 22112 9466 22140 10118
rect 22296 10010 22324 10134
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22204 9982 22324 10010
rect 22204 9586 22232 9982
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 21836 9450 22140 9466
rect 21824 9444 22140 9450
rect 21876 9438 22140 9444
rect 22192 9444 22244 9450
rect 21824 9386 21876 9392
rect 22192 9386 22244 9392
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 21180 9036 21232 9042
rect 21180 8978 21232 8984
rect 20088 8634 20116 8978
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 18932 7692 19380 7698
rect 18880 7686 19380 7692
rect 18892 7670 19380 7686
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18800 6934 18828 7142
rect 19352 7002 19380 7670
rect 19536 7002 19564 7890
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 19996 6866 20024 7278
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 18694 6760 18750 6769
rect 18694 6695 18750 6704
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18616 6458 18644 6598
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16960 5370 16988 5714
rect 17880 5534 17908 5850
rect 18616 5778 18644 6394
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18972 6248 19024 6254
rect 19076 6236 19104 6598
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 19024 6208 19104 6236
rect 18972 6190 19024 6196
rect 18708 5846 18736 6190
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19168 5846 19196 6054
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 18616 5534 18644 5714
rect 17880 5506 18000 5534
rect 18616 5506 18736 5534
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 17972 5166 18000 5506
rect 18708 5166 18736 5506
rect 19352 5370 19380 5714
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 20088 5370 20116 7890
rect 20534 7848 20590 7857
rect 20534 7783 20590 7792
rect 20548 7478 20576 7783
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20640 7546 20668 7686
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20718 7304 20774 7313
rect 20718 7239 20720 7248
rect 20772 7239 20774 7248
rect 20720 7210 20772 7216
rect 20916 6866 20944 8978
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 21100 8430 21128 8842
rect 21192 8634 21220 8978
rect 22204 8838 22232 9386
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21284 7546 21312 7686
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21744 7342 21772 8230
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20364 6254 20392 6598
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20640 5914 20668 6802
rect 20732 6254 20760 6802
rect 20824 6458 20852 6802
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20732 5817 20760 6190
rect 20718 5808 20774 5817
rect 20718 5743 20774 5752
rect 21468 5370 21496 7278
rect 22296 6798 22324 9862
rect 22376 9512 22428 9518
rect 22376 9454 22428 9460
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22388 9178 22416 9454
rect 22480 9382 22508 9454
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 22480 8362 22508 8502
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22664 7886 22692 10066
rect 22756 8430 22784 10968
rect 23020 10950 23072 10956
rect 23112 11008 23164 11014
rect 23112 10950 23164 10956
rect 23032 10606 23060 10950
rect 23676 10606 23704 11086
rect 23020 10600 23072 10606
rect 23020 10542 23072 10548
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23112 10532 23164 10538
rect 23112 10474 23164 10480
rect 23124 10130 23152 10474
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23400 9722 23428 10066
rect 24412 10062 24440 13738
rect 24504 12986 24532 13806
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 24872 13530 24900 13670
rect 24964 13546 24992 13738
rect 24860 13524 24912 13530
rect 24964 13518 25084 13546
rect 25148 13530 25176 13806
rect 24860 13466 24912 13472
rect 25056 13433 25084 13518
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25042 13424 25098 13433
rect 25042 13359 25098 13368
rect 25136 13388 25188 13394
rect 24584 13184 24636 13190
rect 24584 13126 24636 13132
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24596 12850 24624 13126
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24780 12345 24808 12718
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24766 12336 24822 12345
rect 24766 12271 24822 12280
rect 24872 10130 24900 12582
rect 25056 12374 25084 13359
rect 25136 13330 25188 13336
rect 25148 12986 25176 13330
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 25516 12306 25544 14214
rect 25596 13728 25648 13734
rect 25596 13670 25648 13676
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25240 11218 25268 12242
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 24412 9674 24440 9998
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24412 9646 24532 9674
rect 24308 9580 24360 9586
rect 24308 9522 24360 9528
rect 23020 9512 23072 9518
rect 24320 9489 24348 9522
rect 24504 9518 24532 9646
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24596 9518 24624 9590
rect 24492 9512 24544 9518
rect 23020 9454 23072 9460
rect 24306 9480 24362 9489
rect 23032 9042 23060 9454
rect 24492 9454 24544 9460
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24688 9450 24716 9862
rect 25148 9518 25176 10542
rect 25240 10198 25268 11154
rect 25608 10674 25636 13670
rect 26252 13462 26280 14214
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 31217 13628 31525 13637
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 25780 12300 25832 12306
rect 25780 12242 25832 12248
rect 25792 11286 25820 12242
rect 25780 11280 25832 11286
rect 25976 11257 26004 12718
rect 26160 12306 26188 13330
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 26884 13184 26936 13190
rect 26884 13126 26936 13132
rect 26896 12782 26924 13126
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 26884 12776 26936 12782
rect 26884 12718 26936 12724
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 26424 12708 26476 12714
rect 26424 12650 26476 12656
rect 26240 12640 26292 12646
rect 26240 12582 26292 12588
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 26252 11694 26280 12582
rect 26332 12096 26384 12102
rect 26332 12038 26384 12044
rect 26344 11694 26372 12038
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26160 11286 26188 11494
rect 26148 11280 26200 11286
rect 25780 11222 25832 11228
rect 25962 11248 26018 11257
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25228 10192 25280 10198
rect 25228 10134 25280 10140
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 24306 9415 24362 9424
rect 24676 9444 24728 9450
rect 24676 9386 24728 9392
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22744 8424 22796 8430
rect 22848 8401 22876 8910
rect 23032 8634 23060 8978
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 22744 8366 22796 8372
rect 22834 8392 22890 8401
rect 22756 8090 22784 8366
rect 22834 8327 22890 8336
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 23032 7954 23060 8570
rect 23124 8430 23152 8978
rect 24136 8974 24164 9318
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 23204 8900 23256 8906
rect 23204 8842 23256 8848
rect 23216 8498 23244 8842
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23676 8566 23704 8774
rect 23664 8560 23716 8566
rect 23848 8560 23900 8566
rect 23664 8502 23716 8508
rect 23768 8508 23848 8514
rect 23768 8502 23900 8508
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23768 8486 23888 8502
rect 23112 8424 23164 8430
rect 23112 8366 23164 8372
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 23124 7342 23152 8366
rect 23204 8356 23256 8362
rect 23204 8298 23256 8304
rect 23216 8090 23244 8298
rect 23768 8294 23796 8486
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23860 7954 23888 8486
rect 23940 8288 23992 8294
rect 23992 8248 24072 8276
rect 23940 8230 23992 8236
rect 24044 7954 24072 8248
rect 24136 7954 24164 8910
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24412 8430 24440 8774
rect 24504 8634 24532 8774
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24400 7948 24452 7954
rect 24400 7890 24452 7896
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23112 7336 23164 7342
rect 22742 7304 22798 7313
rect 23164 7296 23244 7324
rect 23112 7278 23164 7284
rect 22742 7239 22798 7248
rect 22756 6798 22784 7239
rect 23216 6866 23244 7296
rect 23308 7002 23336 7822
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 23768 7410 23796 7686
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 21732 6792 21784 6798
rect 21730 6760 21732 6769
rect 22284 6792 22336 6798
rect 21784 6760 21786 6769
rect 22284 6734 22336 6740
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 21730 6695 21786 6704
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 22940 6254 22968 6666
rect 23492 6458 23520 6734
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23860 6254 23888 7414
rect 24044 7410 24072 7686
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 23952 6866 23980 7210
rect 24136 7018 24164 7890
rect 24412 7546 24440 7890
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24964 7342 24992 7686
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 24044 6990 24164 7018
rect 24044 6866 24072 6990
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23124 5914 23152 6054
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 24044 5930 24072 6802
rect 24136 6458 24164 6802
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24872 6322 24900 7142
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24124 6248 24176 6254
rect 24124 6190 24176 6196
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23860 5902 24072 5930
rect 24136 5914 24164 6190
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 24412 5914 24440 6122
rect 23860 5794 23888 5902
rect 23400 5778 23888 5794
rect 24044 5778 24072 5902
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 23388 5772 23888 5778
rect 23440 5766 23888 5772
rect 23388 5714 23440 5720
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18420 5092 18472 5098
rect 18420 5034 18472 5040
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17972 4758 18000 4966
rect 18432 4826 18460 5034
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4826 20576 4966
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18616 4214 18644 4626
rect 19536 4282 19564 4694
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18248 3942 18276 4150
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18984 3602 19012 3878
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 2922 16988 3334
rect 18432 3126 18460 3538
rect 18420 3120 18472 3126
rect 18420 3062 18472 3068
rect 19352 2990 19380 4014
rect 20456 3942 20484 4694
rect 20548 4078 20576 4762
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4078 20668 4422
rect 20824 4282 20852 4558
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 21008 4078 21036 4490
rect 21468 4486 21496 4626
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 3670 21128 3878
rect 21468 3738 21496 4422
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 21088 3664 21140 3670
rect 21088 3606 21140 3612
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 20088 3194 20116 3606
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 21100 2990 21128 3606
rect 21468 3058 21496 3674
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21836 3194 21864 3470
rect 21928 3398 21956 4422
rect 22112 4010 22140 5714
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 23388 4752 23440 4758
rect 23388 4694 23440 4700
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22664 4570 22692 4626
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 22480 4542 22692 4570
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 22204 3534 22232 4490
rect 22480 4486 22508 4542
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22572 4146 22600 4422
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22940 4010 22968 4422
rect 23400 4282 23428 4694
rect 23572 4684 23624 4690
rect 23860 4672 23888 5766
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 23624 4644 23888 4672
rect 23572 4626 23624 4632
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23584 4146 23612 4626
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 22204 2922 22232 3470
rect 23860 3194 23888 3946
rect 23952 3738 23980 5714
rect 25056 4826 25084 7278
rect 25240 6458 25268 8910
rect 25332 8634 25360 10542
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25424 9722 25452 10066
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25608 9110 25636 10066
rect 25792 9654 25820 11222
rect 26148 11222 26200 11228
rect 25962 11183 25964 11192
rect 26016 11183 26018 11192
rect 25964 11154 26016 11160
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 26160 10606 26188 10950
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 25872 9920 25924 9926
rect 25872 9862 25924 9868
rect 25780 9648 25832 9654
rect 25884 9625 25912 9862
rect 25780 9590 25832 9596
rect 25870 9616 25926 9625
rect 25596 9104 25648 9110
rect 25596 9046 25648 9052
rect 25792 8634 25820 9590
rect 25870 9551 25926 9560
rect 25964 9512 26016 9518
rect 25962 9480 25964 9489
rect 26056 9512 26108 9518
rect 26016 9480 26018 9489
rect 26056 9454 26108 9460
rect 25962 9415 26018 9424
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25688 8424 25740 8430
rect 25688 8366 25740 8372
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 25700 8090 25728 8366
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25884 7546 25912 8366
rect 25976 8090 26004 8366
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 26068 7478 26096 9454
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26344 8974 26372 9114
rect 26436 9042 26464 12650
rect 27080 12102 27108 12718
rect 27252 12708 27304 12714
rect 27252 12650 27304 12656
rect 27264 12442 27292 12650
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 27250 12336 27306 12345
rect 27250 12271 27306 12280
rect 27712 12300 27764 12306
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 27264 11694 27292 12271
rect 27712 12242 27764 12248
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 27724 11898 27752 12242
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 26712 9722 26740 11630
rect 27160 11008 27212 11014
rect 27160 10950 27212 10956
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26896 9722 26924 10066
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 27068 9716 27120 9722
rect 27068 9658 27120 9664
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26608 9104 26660 9110
rect 26608 9046 26660 9052
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 26148 8900 26200 8906
rect 26148 8842 26200 8848
rect 26160 8294 26188 8842
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26160 7886 26188 8230
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 26056 7472 26108 7478
rect 26056 7414 26108 7420
rect 26252 7342 26280 7754
rect 26436 7342 26464 8978
rect 26620 8838 26648 9046
rect 26700 9036 26752 9042
rect 26700 8978 26752 8984
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26712 7834 26740 8978
rect 26896 8945 26924 9454
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 26882 8936 26938 8945
rect 26882 8871 26938 8880
rect 26896 8430 26924 8871
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26884 8288 26936 8294
rect 26988 8242 27016 9318
rect 27080 9110 27108 9658
rect 27172 9466 27200 10950
rect 27365 10908 27673 10917
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27172 9438 27292 9466
rect 27068 9104 27120 9110
rect 27264 9058 27292 9438
rect 27068 9046 27120 9052
rect 27172 9030 27292 9058
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 27080 8430 27108 8842
rect 27172 8430 27200 9030
rect 27356 8906 27384 9522
rect 27816 9518 27844 13194
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 29276 12232 29328 12238
rect 29276 12174 29328 12180
rect 29288 11218 29316 12174
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 28080 11212 28132 11218
rect 28080 11154 28132 11160
rect 29276 11212 29328 11218
rect 29276 11154 29328 11160
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27896 10124 27948 10130
rect 27896 10066 27948 10072
rect 27908 9722 27936 10066
rect 28000 10062 28028 11086
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 28000 9722 28028 9862
rect 27896 9716 27948 9722
rect 27896 9658 27948 9664
rect 27988 9716 28040 9722
rect 27988 9658 28040 9664
rect 28092 9518 28120 11154
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 27448 8906 27476 9454
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 28092 9110 28120 9318
rect 28080 9104 28132 9110
rect 28080 9046 28132 9052
rect 27988 9036 28040 9042
rect 27988 8978 28040 8984
rect 27804 8968 27856 8974
rect 27526 8936 27582 8945
rect 27344 8900 27396 8906
rect 27344 8842 27396 8848
rect 27436 8900 27488 8906
rect 27804 8910 27856 8916
rect 27526 8871 27528 8880
rect 27436 8842 27488 8848
rect 27580 8871 27582 8880
rect 27528 8842 27580 8848
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27264 8634 27292 8774
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 27816 8634 27844 8910
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27252 8628 27304 8634
rect 27252 8570 27304 8576
rect 27804 8628 27856 8634
rect 27804 8570 27856 8576
rect 27620 8560 27672 8566
rect 27620 8502 27672 8508
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 27172 8294 27200 8366
rect 27632 8294 27660 8502
rect 27908 8430 27936 8774
rect 27896 8424 27948 8430
rect 27896 8366 27948 8372
rect 26936 8236 27016 8242
rect 26884 8230 27016 8236
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 27160 8288 27212 8294
rect 27160 8230 27212 8236
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 26804 8022 26832 8230
rect 26896 8214 27016 8230
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 26896 7954 26924 8214
rect 27080 8129 27108 8230
rect 27066 8120 27122 8129
rect 27264 8106 27292 8230
rect 27066 8055 27122 8064
rect 27172 8078 27292 8106
rect 27172 7954 27200 8078
rect 27816 8022 27844 8230
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 28000 7954 28028 8978
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28092 7954 28120 8910
rect 29012 8430 29040 11086
rect 31668 10532 31720 10538
rect 31668 10474 31720 10480
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31680 10305 31708 10474
rect 31666 10296 31722 10305
rect 31666 10231 31722 10240
rect 29460 9920 29512 9926
rect 29460 9862 29512 9868
rect 29472 9518 29500 9862
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 29460 9512 29512 9518
rect 29460 9454 29512 9460
rect 29196 9042 29224 9454
rect 29368 9444 29420 9450
rect 29368 9386 29420 9392
rect 29380 9110 29408 9386
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 31217 9211 31525 9220
rect 29368 9104 29420 9110
rect 29368 9046 29420 9052
rect 30012 9104 30064 9110
rect 30012 9046 30064 9052
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29736 9036 29788 9042
rect 29736 8978 29788 8984
rect 29000 8424 29052 8430
rect 29000 8366 29052 8372
rect 26884 7948 26936 7954
rect 26884 7890 26936 7896
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 27252 7948 27304 7954
rect 27252 7890 27304 7896
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 28080 7948 28132 7954
rect 28080 7890 28132 7896
rect 28172 7948 28224 7954
rect 28172 7890 28224 7896
rect 26712 7806 26832 7834
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 25320 7268 25372 7274
rect 25320 7210 25372 7216
rect 26608 7268 26660 7274
rect 26608 7210 26660 7216
rect 25332 7002 25360 7210
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 26160 6934 26188 7142
rect 26148 6928 26200 6934
rect 26148 6870 26200 6876
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 25976 6254 26004 6394
rect 25964 6248 26016 6254
rect 25964 6190 26016 6196
rect 26240 6248 26292 6254
rect 26240 6190 26292 6196
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 26252 3942 26280 6190
rect 26436 5778 26464 6734
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 26528 5914 26556 6122
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26620 5574 26648 7210
rect 26804 7206 26832 7806
rect 26792 7200 26844 7206
rect 26792 7142 26844 7148
rect 26804 6866 26832 7142
rect 26896 7002 26924 7890
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 27172 7342 27200 7686
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 26884 6996 26936 7002
rect 26884 6938 26936 6944
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26712 6118 26740 6666
rect 26988 6254 27016 7278
rect 27172 6866 27200 7278
rect 27264 7274 27292 7890
rect 27526 7848 27582 7857
rect 27526 7783 27528 7792
rect 27580 7783 27582 7792
rect 27986 7848 28042 7857
rect 27986 7783 27988 7792
rect 27528 7754 27580 7760
rect 28040 7783 28042 7792
rect 27988 7754 28040 7760
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 27365 7579 27673 7588
rect 28000 7342 28028 7754
rect 27988 7336 28040 7342
rect 27988 7278 28040 7284
rect 27252 7268 27304 7274
rect 27252 7210 27304 7216
rect 27712 7268 27764 7274
rect 27712 7210 27764 7216
rect 27252 6928 27304 6934
rect 27724 6905 27752 7210
rect 27252 6870 27304 6876
rect 27710 6896 27766 6905
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 27160 6656 27212 6662
rect 27160 6598 27212 6604
rect 27172 6254 27200 6598
rect 27264 6458 27292 6870
rect 28092 6866 28120 7890
rect 28184 7546 28212 7890
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 29012 7410 29040 8366
rect 29748 7954 29776 8978
rect 30024 7954 30052 9046
rect 30196 9036 30248 9042
rect 30196 8978 30248 8984
rect 30208 8634 30236 8978
rect 30196 8628 30248 8634
rect 30196 8570 30248 8576
rect 31217 8188 31525 8197
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 30746 8120 30802 8129
rect 31217 8123 31525 8132
rect 30746 8055 30802 8064
rect 30380 8016 30432 8022
rect 30380 7958 30432 7964
rect 29736 7948 29788 7954
rect 29736 7890 29788 7896
rect 30012 7948 30064 7954
rect 30012 7890 30064 7896
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 27710 6831 27766 6840
rect 28080 6860 28132 6866
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 27160 6248 27212 6254
rect 27160 6190 27212 6196
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 26712 5778 26740 6054
rect 26700 5772 26752 5778
rect 26700 5714 26752 5720
rect 27344 5772 27396 5778
rect 27344 5714 27396 5720
rect 26608 5568 26660 5574
rect 27356 5534 27384 5714
rect 26608 5510 26660 5516
rect 27264 5506 27384 5534
rect 27264 5370 27292 5506
rect 27365 5468 27673 5477
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 27724 5370 27752 6831
rect 28080 6802 28132 6808
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28736 6458 28764 6802
rect 28724 6452 28776 6458
rect 28724 6394 28776 6400
rect 29012 5778 29040 7346
rect 29748 6866 29776 7890
rect 30024 6934 30052 7890
rect 30392 7546 30420 7958
rect 30760 7954 30788 8055
rect 30748 7948 30800 7954
rect 30748 7890 30800 7896
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31036 7585 31064 7822
rect 31022 7576 31078 7585
rect 30380 7540 30432 7546
rect 31022 7511 31078 7520
rect 30380 7482 30432 7488
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 30012 6928 30064 6934
rect 30012 6870 30064 6876
rect 29092 6860 29144 6866
rect 29092 6802 29144 6808
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 29104 5914 29132 6802
rect 29366 6760 29422 6769
rect 29366 6695 29368 6704
rect 29420 6695 29422 6704
rect 29368 6666 29420 6672
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 29092 5908 29144 5914
rect 29092 5850 29144 5856
rect 29000 5772 29052 5778
rect 29000 5714 29052 5720
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27712 5364 27764 5370
rect 27712 5306 27764 5312
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 31217 2748 31525 2757
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 16304 1012 16356 1018
rect 16304 954 16356 960
rect 16396 1012 16448 1018
rect 16396 954 16448 960
rect 16856 1012 16908 1018
rect 16856 954 16908 960
rect 14280 808 14332 814
rect 14280 750 14332 756
rect 15568 808 15620 814
rect 15568 750 15620 756
rect 16212 808 16264 814
rect 16764 808 16816 814
rect 16264 768 16344 796
rect 16212 750 16264 756
rect 14292 490 14320 750
rect 15580 490 15608 750
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 14200 462 14320 490
rect 15488 462 15608 490
rect 14200 400 14228 462
rect 15488 400 15516 462
rect 18 0 74 400
rect 662 0 718 400
rect 1306 0 1362 400
rect 1950 0 2006 400
rect 2594 0 2650 400
rect 3238 0 3294 400
rect 3882 0 3938 400
rect 4526 0 4582 400
rect 5170 0 5226 400
rect 5814 0 5870 400
rect 6458 0 6514 400
rect 7102 0 7158 400
rect 7746 0 7802 400
rect 8390 0 8446 400
rect 13542 0 13598 400
rect 14186 0 14242 400
rect 15474 0 15530 400
rect 16118 354 16174 400
rect 16316 354 16344 768
rect 16764 750 16816 756
rect 18788 808 18840 814
rect 18788 750 18840 756
rect 16776 400 16804 750
rect 18800 490 18828 750
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 18708 462 18828 490
rect 18708 400 18736 462
rect 16118 326 16344 354
rect 16118 0 16174 326
rect 16762 0 16818 400
rect 18694 0 18750 400
<< via2 >>
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 846 14320 902 14376
rect 846 10240 902 10296
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 4066 13252 4122 13288
rect 4066 13232 4068 13252
rect 4068 13232 4120 13252
rect 4120 13232 4122 13252
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 3514 12416 3570 12472
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 4802 12164 4858 12200
rect 4802 12144 4804 12164
rect 4804 12144 4856 12164
rect 4856 12144 4858 12164
rect 5446 12280 5502 12336
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 6826 12436 6882 12472
rect 6826 12416 6828 12436
rect 6828 12416 6880 12436
rect 6880 12416 6882 12436
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 7286 11600 7342 11656
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 8022 11192 8078 11248
rect 8114 11056 8170 11112
rect 8666 11600 8722 11656
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 9126 11192 9182 11248
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 6458 7248 6514 7304
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 7378 8356 7434 8392
rect 7378 8336 7380 8356
rect 7380 8336 7432 8356
rect 7432 8336 7434 8356
rect 9218 11056 9274 11112
rect 10782 13504 10838 13560
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 8206 7284 8208 7304
rect 8208 7284 8260 7304
rect 8260 7284 8262 7304
rect 8206 7248 8262 7284
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 7194 5616 7250 5672
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 10046 9560 10102 9616
rect 11058 11772 11060 11792
rect 11060 11772 11112 11792
rect 11112 11772 11114 11792
rect 11058 11736 11114 11772
rect 11058 11636 11060 11656
rect 11060 11636 11112 11656
rect 11112 11636 11114 11656
rect 11058 11600 11114 11636
rect 9954 8200 10010 8256
rect 10506 8200 10562 8256
rect 11426 13368 11482 13424
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 12070 12724 12072 12744
rect 12072 12724 12124 12744
rect 12124 12724 12126 12744
rect 12070 12688 12126 12724
rect 11426 11212 11482 11248
rect 11426 11192 11428 11212
rect 11428 11192 11480 11212
rect 11480 11192 11482 11212
rect 11334 9016 11390 9072
rect 10230 5752 10286 5808
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 13726 13368 13782 13424
rect 13542 13232 13598 13288
rect 12622 11736 12678 11792
rect 12530 11600 12586 11656
rect 12714 11600 12770 11656
rect 12806 11192 12862 11248
rect 13542 11872 13598 11928
rect 14646 12960 14702 13016
rect 13358 11056 13414 11112
rect 13818 11056 13874 11112
rect 13082 10648 13138 10704
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 12806 9036 12862 9072
rect 12806 9016 12808 9036
rect 12808 9016 12860 9036
rect 12860 9016 12862 9036
rect 13266 9036 13322 9072
rect 13266 9016 13268 9036
rect 13268 9016 13320 9036
rect 13320 9016 13322 9036
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 12438 8608 12494 8664
rect 11794 7792 11850 7848
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 11702 6704 11758 6760
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 15382 13504 15438 13560
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 31022 18400 31078 18456
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 16118 14456 16174 14512
rect 16578 14456 16634 14512
rect 17498 15000 17554 15056
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 17498 13368 17554 13424
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 17314 13232 17370 13288
rect 15290 11328 15346 11384
rect 15842 12300 15898 12336
rect 15842 12280 15844 12300
rect 15844 12280 15896 12300
rect 15896 12280 15898 12300
rect 15750 12144 15806 12200
rect 15750 11600 15806 11656
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 14094 7248 14150 7304
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 16302 9016 16358 9072
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 16670 9016 16726 9072
rect 12254 3440 12310 3496
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 15014 6860 15070 6896
rect 15014 6840 15016 6860
rect 15016 6840 15068 6860
rect 15068 6840 15070 6860
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15106 5616 15162 5672
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 14646 3460 14702 3496
rect 14646 3440 14648 3460
rect 14648 3440 14700 3460
rect 14700 3440 14702 3460
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 16578 7792 16634 7848
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 18326 14456 18382 14512
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 18142 12960 18198 13016
rect 17222 11056 17278 11112
rect 17038 8608 17094 8664
rect 18878 12180 18880 12200
rect 18880 12180 18932 12200
rect 18932 12180 18934 12200
rect 18878 12144 18934 12180
rect 19154 12688 19210 12744
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 23662 15000 23718 15056
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 20442 13404 20444 13424
rect 20444 13404 20496 13424
rect 20496 13404 20498 13424
rect 20442 13368 20498 13404
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 20718 12688 20774 12744
rect 19890 12280 19946 12336
rect 19154 11892 19210 11928
rect 19154 11872 19156 11892
rect 19156 11872 19208 11892
rect 19208 11872 19210 11892
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 18970 11600 19026 11656
rect 19890 11056 19946 11112
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 18510 8236 18512 8256
rect 18512 8236 18564 8256
rect 18564 8236 18566 8256
rect 18510 8200 18566 8236
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 20902 12300 20958 12336
rect 20902 12280 20904 12300
rect 20904 12280 20956 12300
rect 20956 12280 20958 12300
rect 20350 10648 20406 10704
rect 21638 12144 21694 12200
rect 22650 11872 22706 11928
rect 22558 11736 22614 11792
rect 21730 11600 21786 11656
rect 21178 11056 21234 11112
rect 23018 11872 23074 11928
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 24306 12724 24308 12744
rect 24308 12724 24360 12744
rect 24360 12724 24362 12744
rect 23662 11756 23718 11792
rect 23662 11736 23664 11756
rect 23664 11736 23716 11756
rect 23716 11736 23718 11756
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 24306 12688 24362 12724
rect 23938 11600 23994 11656
rect 19062 8200 19118 8256
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 18694 6704 18750 6760
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 20534 7792 20590 7848
rect 20718 7268 20774 7304
rect 20718 7248 20720 7268
rect 20720 7248 20772 7268
rect 20772 7248 20774 7268
rect 20718 5752 20774 5808
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 25042 13368 25098 13424
rect 24766 12280 24822 12336
rect 24306 9424 24362 9480
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 22834 8336 22890 8392
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 22742 7248 22798 7304
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 21730 6740 21732 6760
rect 21732 6740 21784 6760
rect 21784 6740 21786 6760
rect 21730 6704 21786 6740
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 25962 11212 26018 11248
rect 25962 11192 25964 11212
rect 25964 11192 26016 11212
rect 26016 11192 26018 11212
rect 25870 9560 25926 9616
rect 25962 9460 25964 9480
rect 25964 9460 26016 9480
rect 26016 9460 26018 9480
rect 25962 9424 26018 9460
rect 27250 12280 27306 12336
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 26882 8880 26938 8936
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 27526 8900 27582 8936
rect 27526 8880 27528 8900
rect 27528 8880 27580 8900
rect 27580 8880 27582 8900
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 27066 8064 27122 8120
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10240 31722 10296
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 27526 7812 27582 7848
rect 27526 7792 27528 7812
rect 27528 7792 27580 7812
rect 27580 7792 27582 7812
rect 27986 7812 28042 7848
rect 27986 7792 27988 7812
rect 27988 7792 28040 7812
rect 28040 7792 28042 7812
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 27710 6840 27766 6896
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 30746 8064 30802 8120
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 31022 7520 31078 7576
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 29366 6724 29422 6760
rect 29366 6704 29368 6724
rect 29368 6704 29420 6724
rect 29420 6704 29422 6724
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
<< metal3 >>
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31213 19007 31529 19008
rect 4246 18528 4562 18529
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 31017 18458 31083 18461
rect 31600 18458 32000 18488
rect 31017 18456 32000 18458
rect 31017 18400 31022 18456
rect 31078 18400 32000 18456
rect 31017 18398 32000 18400
rect 31017 18395 31083 18398
rect 31600 18368 32000 18398
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 17493 15058 17559 15061
rect 23657 15058 23723 15061
rect 17493 15056 23723 15058
rect 17493 15000 17498 15056
rect 17554 15000 23662 15056
rect 23718 15000 23723 15056
rect 17493 14998 23723 15000
rect 17493 14995 17559 14998
rect 23657 14995 23723 14998
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 16113 14514 16179 14517
rect 16573 14514 16639 14517
rect 18321 14514 18387 14517
rect 16113 14512 18387 14514
rect 16113 14456 16118 14512
rect 16174 14456 16578 14512
rect 16634 14456 18326 14512
rect 18382 14456 18387 14512
rect 16113 14454 18387 14456
rect 16113 14451 16179 14454
rect 16573 14451 16639 14454
rect 18321 14451 18387 14454
rect 0 14378 400 14408
rect 841 14378 907 14381
rect 0 14376 907 14378
rect 0 14320 846 14376
rect 902 14320 907 14376
rect 0 14318 907 14320
rect 0 14288 400 14318
rect 841 14315 907 14318
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31213 13567 31529 13568
rect 10777 13562 10843 13565
rect 15377 13562 15443 13565
rect 10777 13560 15443 13562
rect 10777 13504 10782 13560
rect 10838 13504 15382 13560
rect 15438 13504 15443 13560
rect 10777 13502 15443 13504
rect 10777 13499 10843 13502
rect 15377 13499 15443 13502
rect 11421 13426 11487 13429
rect 13721 13426 13787 13429
rect 17493 13426 17559 13429
rect 11421 13424 17559 13426
rect 11421 13368 11426 13424
rect 11482 13368 13726 13424
rect 13782 13368 17498 13424
rect 17554 13368 17559 13424
rect 11421 13366 17559 13368
rect 11421 13363 11487 13366
rect 13721 13363 13787 13366
rect 17493 13363 17559 13366
rect 20437 13426 20503 13429
rect 25037 13426 25103 13429
rect 20437 13424 25103 13426
rect 20437 13368 20442 13424
rect 20498 13368 25042 13424
rect 25098 13368 25103 13424
rect 20437 13366 25103 13368
rect 20437 13363 20503 13366
rect 25037 13363 25103 13366
rect 4061 13290 4127 13293
rect 13537 13290 13603 13293
rect 17309 13290 17375 13293
rect 4061 13288 17375 13290
rect 4061 13232 4066 13288
rect 4122 13232 13542 13288
rect 13598 13232 17314 13288
rect 17370 13232 17375 13288
rect 4061 13230 17375 13232
rect 4061 13227 4127 13230
rect 13537 13227 13603 13230
rect 17309 13227 17375 13230
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 14641 13018 14707 13021
rect 18137 13018 18203 13021
rect 14641 13016 18203 13018
rect 14641 12960 14646 13016
rect 14702 12960 18142 13016
rect 18198 12960 18203 13016
rect 14641 12958 18203 12960
rect 14641 12955 14707 12958
rect 18137 12955 18203 12958
rect 12065 12746 12131 12749
rect 19149 12746 19215 12749
rect 12065 12744 19215 12746
rect 12065 12688 12070 12744
rect 12126 12688 19154 12744
rect 19210 12688 19215 12744
rect 12065 12686 19215 12688
rect 12065 12683 12131 12686
rect 19149 12683 19215 12686
rect 20713 12746 20779 12749
rect 24301 12746 24367 12749
rect 20713 12744 24367 12746
rect 20713 12688 20718 12744
rect 20774 12688 24306 12744
rect 24362 12688 24367 12744
rect 20713 12686 24367 12688
rect 20713 12683 20779 12686
rect 24301 12683 24367 12686
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 3509 12474 3575 12477
rect 6821 12474 6887 12477
rect 3509 12472 6887 12474
rect 3509 12416 3514 12472
rect 3570 12416 6826 12472
rect 6882 12416 6887 12472
rect 3509 12414 6887 12416
rect 3509 12411 3575 12414
rect 6821 12411 6887 12414
rect 5441 12338 5507 12341
rect 15837 12338 15903 12341
rect 5441 12336 15903 12338
rect 5441 12280 5446 12336
rect 5502 12280 15842 12336
rect 15898 12280 15903 12336
rect 5441 12278 15903 12280
rect 5441 12275 5507 12278
rect 15837 12275 15903 12278
rect 19885 12338 19951 12341
rect 20897 12338 20963 12341
rect 24761 12338 24827 12341
rect 19885 12336 24827 12338
rect 19885 12280 19890 12336
rect 19946 12280 20902 12336
rect 20958 12280 24766 12336
rect 24822 12280 24827 12336
rect 19885 12278 24827 12280
rect 19885 12275 19951 12278
rect 20897 12275 20963 12278
rect 24761 12275 24827 12278
rect 27245 12338 27311 12341
rect 31600 12338 32000 12368
rect 27245 12336 32000 12338
rect 27245 12280 27250 12336
rect 27306 12280 32000 12336
rect 27245 12278 32000 12280
rect 27245 12275 27311 12278
rect 31600 12248 32000 12278
rect 4797 12202 4863 12205
rect 15745 12202 15811 12205
rect 4797 12200 15811 12202
rect 4797 12144 4802 12200
rect 4858 12144 15750 12200
rect 15806 12144 15811 12200
rect 4797 12142 15811 12144
rect 4797 12139 4863 12142
rect 15745 12139 15811 12142
rect 18873 12202 18939 12205
rect 21633 12202 21699 12205
rect 18873 12200 21699 12202
rect 18873 12144 18878 12200
rect 18934 12144 21638 12200
rect 21694 12144 21699 12200
rect 18873 12142 21699 12144
rect 18873 12139 18939 12142
rect 21633 12139 21699 12142
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 13537 11930 13603 11933
rect 19149 11930 19215 11933
rect 13537 11928 19215 11930
rect 13537 11872 13542 11928
rect 13598 11872 19154 11928
rect 19210 11872 19215 11928
rect 13537 11870 19215 11872
rect 13537 11867 13603 11870
rect 19149 11867 19215 11870
rect 22645 11930 22711 11933
rect 23013 11930 23079 11933
rect 22645 11928 23079 11930
rect 22645 11872 22650 11928
rect 22706 11872 23018 11928
rect 23074 11872 23079 11928
rect 22645 11870 23079 11872
rect 22645 11867 22711 11870
rect 23013 11867 23079 11870
rect 11053 11794 11119 11797
rect 12617 11794 12683 11797
rect 11053 11792 12683 11794
rect 11053 11736 11058 11792
rect 11114 11736 12622 11792
rect 12678 11736 12683 11792
rect 11053 11734 12683 11736
rect 11053 11731 11119 11734
rect 12617 11731 12683 11734
rect 22553 11794 22619 11797
rect 23657 11794 23723 11797
rect 22553 11792 23723 11794
rect 22553 11736 22558 11792
rect 22614 11736 23662 11792
rect 23718 11736 23723 11792
rect 22553 11734 23723 11736
rect 22553 11731 22619 11734
rect 23657 11731 23723 11734
rect 7281 11658 7347 11661
rect 8661 11658 8727 11661
rect 7281 11656 8727 11658
rect 7281 11600 7286 11656
rect 7342 11600 8666 11656
rect 8722 11600 8727 11656
rect 7281 11598 8727 11600
rect 7281 11595 7347 11598
rect 8661 11595 8727 11598
rect 11053 11658 11119 11661
rect 12525 11658 12591 11661
rect 11053 11656 12591 11658
rect 11053 11600 11058 11656
rect 11114 11600 12530 11656
rect 12586 11600 12591 11656
rect 11053 11598 12591 11600
rect 11053 11595 11119 11598
rect 12525 11595 12591 11598
rect 12709 11658 12775 11661
rect 15745 11658 15811 11661
rect 18965 11658 19031 11661
rect 21725 11658 21791 11661
rect 23933 11658 23999 11661
rect 12709 11656 23999 11658
rect 12709 11600 12714 11656
rect 12770 11600 15750 11656
rect 15806 11600 18970 11656
rect 19026 11600 21730 11656
rect 21786 11600 23938 11656
rect 23994 11600 23999 11656
rect 12709 11598 23999 11600
rect 12709 11595 12775 11598
rect 15745 11595 15811 11598
rect 18965 11595 19031 11598
rect 21725 11595 21791 11598
rect 23933 11595 23999 11598
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 15285 11384 15351 11389
rect 15285 11328 15290 11384
rect 15346 11328 15351 11384
rect 15285 11323 15351 11328
rect 8017 11250 8083 11253
rect 9121 11250 9187 11253
rect 11421 11250 11487 11253
rect 12801 11250 12867 11253
rect 8017 11248 12867 11250
rect 8017 11192 8022 11248
rect 8078 11192 9126 11248
rect 9182 11192 11426 11248
rect 11482 11192 12806 11248
rect 12862 11192 12867 11248
rect 8017 11190 12867 11192
rect 15288 11250 15348 11323
rect 25957 11250 26023 11253
rect 15288 11248 26023 11250
rect 15288 11192 25962 11248
rect 26018 11192 26023 11248
rect 15288 11190 26023 11192
rect 8017 11187 8083 11190
rect 9121 11187 9187 11190
rect 11421 11187 11487 11190
rect 12801 11187 12867 11190
rect 25957 11187 26023 11190
rect 8109 11114 8175 11117
rect 9213 11114 9279 11117
rect 8109 11112 9279 11114
rect 8109 11056 8114 11112
rect 8170 11056 9218 11112
rect 9274 11056 9279 11112
rect 8109 11054 9279 11056
rect 8109 11051 8175 11054
rect 9213 11051 9279 11054
rect 13353 11114 13419 11117
rect 13813 11114 13879 11117
rect 17217 11114 17283 11117
rect 13353 11112 17283 11114
rect 13353 11056 13358 11112
rect 13414 11056 13818 11112
rect 13874 11056 17222 11112
rect 17278 11056 17283 11112
rect 13353 11054 17283 11056
rect 13353 11051 13419 11054
rect 13813 11051 13879 11054
rect 17217 11051 17283 11054
rect 19885 11114 19951 11117
rect 21173 11114 21239 11117
rect 19885 11112 21239 11114
rect 19885 11056 19890 11112
rect 19946 11056 21178 11112
rect 21234 11056 21239 11112
rect 19885 11054 21239 11056
rect 19885 11051 19951 11054
rect 21173 11051 21239 11054
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 27361 10847 27677 10848
rect 13077 10706 13143 10709
rect 20345 10706 20411 10709
rect 13077 10704 20411 10706
rect 13077 10648 13082 10704
rect 13138 10648 20350 10704
rect 20406 10648 20411 10704
rect 13077 10646 20411 10648
rect 13077 10643 13143 10646
rect 20345 10643 20411 10646
rect 8098 10368 8414 10369
rect 0 10298 400 10328
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 841 10298 907 10301
rect 0 10296 907 10298
rect 0 10240 846 10296
rect 902 10240 907 10296
rect 0 10238 907 10240
rect 0 10208 400 10238
rect 841 10235 907 10238
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 0 9618 400 9648
rect 10041 9618 10107 9621
rect 0 9616 10107 9618
rect 0 9560 10046 9616
rect 10102 9560 10107 9616
rect 0 9558 10107 9560
rect 0 9528 400 9558
rect 10041 9555 10107 9558
rect 25865 9618 25931 9621
rect 31600 9618 32000 9648
rect 25865 9616 32000 9618
rect 25865 9560 25870 9616
rect 25926 9560 32000 9616
rect 25865 9558 32000 9560
rect 25865 9555 25931 9558
rect 31600 9528 32000 9558
rect 24301 9482 24367 9485
rect 25957 9482 26023 9485
rect 24301 9480 26023 9482
rect 24301 9424 24306 9480
rect 24362 9424 25962 9480
rect 26018 9424 26023 9480
rect 24301 9422 26023 9424
rect 24301 9419 24367 9422
rect 25957 9419 26023 9422
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 11329 9074 11395 9077
rect 12801 9074 12867 9077
rect 11329 9072 12867 9074
rect 11329 9016 11334 9072
rect 11390 9016 12806 9072
rect 12862 9016 12867 9072
rect 11329 9014 12867 9016
rect 11329 9011 11395 9014
rect 12801 9011 12867 9014
rect 13261 9074 13327 9077
rect 16297 9074 16363 9077
rect 16665 9074 16731 9077
rect 13261 9072 16731 9074
rect 13261 9016 13266 9072
rect 13322 9016 16302 9072
rect 16358 9016 16670 9072
rect 16726 9016 16731 9072
rect 13261 9014 16731 9016
rect 13261 9011 13327 9014
rect 16297 9011 16363 9014
rect 16665 9011 16731 9014
rect 26877 8938 26943 8941
rect 27521 8938 27587 8941
rect 26877 8936 27587 8938
rect 26877 8880 26882 8936
rect 26938 8880 27526 8936
rect 27582 8880 27587 8936
rect 26877 8878 27587 8880
rect 26877 8875 26943 8878
rect 27521 8875 27587 8878
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 12433 8666 12499 8669
rect 17033 8666 17099 8669
rect 12433 8664 17099 8666
rect 12433 8608 12438 8664
rect 12494 8608 17038 8664
rect 17094 8608 17099 8664
rect 12433 8606 17099 8608
rect 12433 8603 12499 8606
rect 17033 8603 17099 8606
rect 7373 8394 7439 8397
rect 22829 8394 22895 8397
rect 7373 8392 22895 8394
rect 7373 8336 7378 8392
rect 7434 8336 22834 8392
rect 22890 8336 22895 8392
rect 7373 8334 22895 8336
rect 7373 8331 7439 8334
rect 22829 8331 22895 8334
rect 9949 8258 10015 8261
rect 10501 8258 10567 8261
rect 9949 8256 10567 8258
rect 9949 8200 9954 8256
rect 10010 8200 10506 8256
rect 10562 8200 10567 8256
rect 9949 8198 10567 8200
rect 9949 8195 10015 8198
rect 10501 8195 10567 8198
rect 18505 8258 18571 8261
rect 19057 8258 19123 8261
rect 18505 8256 19123 8258
rect 18505 8200 18510 8256
rect 18566 8200 19062 8256
rect 19118 8200 19123 8256
rect 18505 8198 19123 8200
rect 18505 8195 18571 8198
rect 19057 8195 19123 8198
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31213 8127 31529 8128
rect 27061 8122 27127 8125
rect 30741 8122 30807 8125
rect 24810 8120 30807 8122
rect 24810 8064 27066 8120
rect 27122 8064 30746 8120
rect 30802 8064 30807 8120
rect 24810 8062 30807 8064
rect 11789 7850 11855 7853
rect 16573 7850 16639 7853
rect 11789 7848 16639 7850
rect 11789 7792 11794 7848
rect 11850 7792 16578 7848
rect 16634 7792 16639 7848
rect 11789 7790 16639 7792
rect 11789 7787 11855 7790
rect 16573 7787 16639 7790
rect 20529 7850 20595 7853
rect 24810 7850 24870 8062
rect 27061 8059 27127 8062
rect 30741 8059 30807 8062
rect 20529 7848 24870 7850
rect 20529 7792 20534 7848
rect 20590 7792 24870 7848
rect 20529 7790 24870 7792
rect 27521 7850 27587 7853
rect 27981 7850 28047 7853
rect 27521 7848 28047 7850
rect 27521 7792 27526 7848
rect 27582 7792 27986 7848
rect 28042 7792 28047 7848
rect 27521 7790 28047 7792
rect 20529 7787 20595 7790
rect 27521 7787 27587 7790
rect 27981 7787 28047 7790
rect 4246 7648 4562 7649
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 31017 7578 31083 7581
rect 31600 7578 32000 7608
rect 31017 7576 32000 7578
rect 31017 7520 31022 7576
rect 31078 7520 32000 7576
rect 31017 7518 32000 7520
rect 31017 7515 31083 7518
rect 31600 7488 32000 7518
rect 6453 7306 6519 7309
rect 8201 7306 8267 7309
rect 6453 7304 8267 7306
rect 6453 7248 6458 7304
rect 6514 7248 8206 7304
rect 8262 7248 8267 7304
rect 6453 7246 8267 7248
rect 6453 7243 6519 7246
rect 8201 7243 8267 7246
rect 14089 7306 14155 7309
rect 20713 7306 20779 7309
rect 14089 7304 20779 7306
rect 14089 7248 14094 7304
rect 14150 7248 20718 7304
rect 20774 7248 20779 7304
rect 14089 7246 20779 7248
rect 14089 7243 14155 7246
rect 20713 7243 20779 7246
rect 22737 7306 22803 7309
rect 22737 7304 28274 7306
rect 22737 7248 22742 7304
rect 22798 7248 28274 7304
rect 22737 7246 28274 7248
rect 22737 7243 22803 7246
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 15009 6898 15075 6901
rect 27705 6898 27771 6901
rect 15009 6896 27771 6898
rect 15009 6840 15014 6896
rect 15070 6840 27710 6896
rect 27766 6840 27771 6896
rect 15009 6838 27771 6840
rect 28214 6898 28274 7246
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 31600 6898 32000 6928
rect 28214 6838 32000 6898
rect 15009 6835 15075 6838
rect 27705 6835 27771 6838
rect 31600 6808 32000 6838
rect 11697 6762 11763 6765
rect 18689 6762 18755 6765
rect 11697 6760 18755 6762
rect 11697 6704 11702 6760
rect 11758 6704 18694 6760
rect 18750 6704 18755 6760
rect 11697 6702 18755 6704
rect 11697 6699 11763 6702
rect 18689 6699 18755 6702
rect 21725 6762 21791 6765
rect 29361 6762 29427 6765
rect 21725 6760 29427 6762
rect 21725 6704 21730 6760
rect 21786 6704 29366 6760
rect 29422 6704 29427 6760
rect 21725 6702 29427 6704
rect 21725 6699 21791 6702
rect 29361 6699 29427 6702
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 10225 5810 10291 5813
rect 20713 5810 20779 5813
rect 10225 5808 20779 5810
rect 10225 5752 10230 5808
rect 10286 5752 20718 5808
rect 20774 5752 20779 5808
rect 10225 5750 20779 5752
rect 10225 5747 10291 5750
rect 20713 5747 20779 5750
rect 7189 5674 7255 5677
rect 15101 5674 15167 5677
rect 7189 5672 15167 5674
rect 7189 5616 7194 5672
rect 7250 5616 15106 5672
rect 15162 5616 15167 5672
rect 7189 5614 15167 5616
rect 7189 5611 7255 5614
rect 15101 5611 15167 5614
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 27361 5407 27677 5408
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 12249 3498 12315 3501
rect 14641 3498 14707 3501
rect 12249 3496 14707 3498
rect 12249 3440 12254 3496
rect 12310 3440 14646 3496
rect 14702 3440 14707 3496
rect 12249 3438 14707 3440
rect 12249 3435 12315 3438
rect 14641 3435 14707 3438
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11949 12000 12269 13024
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 11949 8736 12269 9760
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 11949 6560 12269 7584
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 15801 15808 16121 16832
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 15801 10368 16121 11392
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15801 4928 16121 5952
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15801 3840 16121 4864
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19654 12000 19974 13024
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19654 7648 19974 8672
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 19654 4384 19974 5408
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 23506 15808 23826 16832
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
use sky130_fd_sc_hd__buf_2  _233_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16560 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _234_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16744 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _235_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16560 0 1 8160
box -38 -48 1418 592
use sky130_fd_sc_hd__clkbuf_4  _236_
timestamp 1701704242
transform 1 0 11960 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _237_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _238_
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _239_
timestamp 1701704242
transform 1 0 16744 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_2  _240_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14628 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _241_
timestamp 1701704242
transform 1 0 12512 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _242_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 30544 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _243_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15272 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _244_
timestamp 1701704242
transform 1 0 13984 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _245_
timestamp 1701704242
transform -1 0 14628 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _246_
timestamp 1701704242
transform 1 0 9936 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _247_
timestamp 1701704242
transform 1 0 24104 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _248_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 26128 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _249_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 19412 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _250_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18216 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _251_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 19596 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _252_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20056 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _253_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9200 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _254_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 24932 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _255_
timestamp 1701704242
transform 1 0 9476 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _256_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 19136 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _257_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20148 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _258_
timestamp 1701704242
transform 1 0 18768 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _259_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 21712 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_4  _260_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 24656 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _261_
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _262_
timestamp 1701704242
transform 1 0 26864 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _263_
timestamp 1701704242
transform 1 0 25300 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _264_
timestamp 1701704242
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1701704242
transform 1 0 21252 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _266_
timestamp 1701704242
transform -1 0 29624 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _267_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 22816 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _268_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 25944 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_4  _269_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 27324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _270_
timestamp 1701704242
transform 1 0 18308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _271_
timestamp 1701704242
transform 1 0 24932 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _272_
timestamp 1701704242
transform -1 0 30176 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _273_
timestamp 1701704242
transform 1 0 25392 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _274_
timestamp 1701704242
transform 1 0 23920 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _275_
timestamp 1701704242
transform 1 0 24656 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _276_
timestamp 1701704242
transform 1 0 25484 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _277_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 26404 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _278_
timestamp 1701704242
transform 1 0 26220 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _279_
timestamp 1701704242
transform 1 0 28704 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _280_
timestamp 1701704242
transform 1 0 20424 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _281_
timestamp 1701704242
transform -1 0 21988 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _282_
timestamp 1701704242
transform 1 0 12420 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _283_
timestamp 1701704242
transform 1 0 19872 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _284_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 21436 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _285_
timestamp 1701704242
transform 1 0 20700 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_4  _286_
timestamp 1701704242
transform -1 0 22816 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _287_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15180 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _288_
timestamp 1701704242
transform 1 0 15180 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _289_
timestamp 1701704242
transform 1 0 14996 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _290_
timestamp 1701704242
transform -1 0 15640 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _291_
timestamp 1701704242
transform -1 0 15916 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _292_
timestamp 1701704242
transform -1 0 16744 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _293_
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _294_
timestamp 1701704242
transform 1 0 14996 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _295_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 17664 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _296_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16560 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _297_
timestamp 1701704242
transform 1 0 10120 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _298_
timestamp 1701704242
transform 1 0 11408 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _299_
timestamp 1701704242
transform 1 0 11040 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _300_
timestamp 1701704242
transform -1 0 12880 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _301_
timestamp 1701704242
transform 1 0 9936 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _302_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 19964 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__a311o_1  _303_
timestamp 1701704242
transform 1 0 18676 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _304_
timestamp 1701704242
transform 1 0 11684 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_4  _305_
timestamp 1701704242
transform -1 0 12696 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _306_
timestamp 1701704242
transform 1 0 10488 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _307_
timestamp 1701704242
transform 1 0 9844 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _308_
timestamp 1701704242
transform 1 0 9568 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _309_
timestamp 1701704242
transform 1 0 10212 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _310_
timestamp 1701704242
transform 1 0 10028 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _311_
timestamp 1701704242
transform 1 0 10120 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _312_
timestamp 1701704242
transform 1 0 9384 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _313_
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _314_
timestamp 1701704242
transform -1 0 6532 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _315_
timestamp 1701704242
transform 1 0 10028 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1701704242
transform -1 0 18400 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1701704242
transform 1 0 18768 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _318_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 19688 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _319_
timestamp 1701704242
transform -1 0 20056 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _320_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20700 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _321_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 21436 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _322_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20056 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _323_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 20792 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _324_
timestamp 1701704242
transform -1 0 21068 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _325_
timestamp 1701704242
transform -1 0 21528 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _326_
timestamp 1701704242
transform 1 0 10764 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _327_
timestamp 1701704242
transform -1 0 11592 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _328_
timestamp 1701704242
transform 1 0 10304 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _329_
timestamp 1701704242
transform -1 0 11684 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _330_
timestamp 1701704242
transform -1 0 11960 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _331_
timestamp 1701704242
transform -1 0 9936 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _332_
timestamp 1701704242
transform -1 0 10488 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _333_
timestamp 1701704242
transform -1 0 9844 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _334_
timestamp 1701704242
transform 1 0 9108 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _335_
timestamp 1701704242
transform 1 0 10212 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _336_
timestamp 1701704242
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _337_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8464 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _338_
timestamp 1701704242
transform 1 0 12788 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _339_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15640 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _340_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15640 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _341_
timestamp 1701704242
transform 1 0 15088 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _342_
timestamp 1701704242
transform 1 0 16560 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _343_
timestamp 1701704242
transform -1 0 16192 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _344_
timestamp 1701704242
transform 1 0 16100 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _345_
timestamp 1701704242
transform -1 0 15088 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _346_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _347_
timestamp 1701704242
transform -1 0 10212 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _348_
timestamp 1701704242
transform 1 0 3404 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _349_
timestamp 1701704242
transform 1 0 5980 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _350_
timestamp 1701704242
transform 1 0 6440 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _351_
timestamp 1701704242
transform -1 0 6716 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _352_
timestamp 1701704242
transform -1 0 4784 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _353_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3680 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _354_
timestamp 1701704242
transform 1 0 4140 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _355_
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _356_
timestamp 1701704242
transform 1 0 20700 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _357_
timestamp 1701704242
transform 1 0 20332 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _358_
timestamp 1701704242
transform 1 0 20608 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _359_
timestamp 1701704242
transform -1 0 20976 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _360_
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _361_
timestamp 1701704242
transform 1 0 21896 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _362_
timestamp 1701704242
transform 1 0 22264 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _363_
timestamp 1701704242
transform 1 0 22540 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _364_
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _365_
timestamp 1701704242
transform -1 0 12512 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _366_
timestamp 1701704242
transform -1 0 11408 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _367_
timestamp 1701704242
transform -1 0 12236 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _368_
timestamp 1701704242
transform -1 0 11684 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _369_
timestamp 1701704242
transform -1 0 11500 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _370_
timestamp 1701704242
transform -1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _371_
timestamp 1701704242
transform 1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _372_
timestamp 1701704242
transform 1 0 9752 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _373_
timestamp 1701704242
transform 1 0 10580 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _374_
timestamp 1701704242
transform 1 0 11040 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _375_
timestamp 1701704242
transform 1 0 9292 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _376_
timestamp 1701704242
transform 1 0 12696 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _377_
timestamp 1701704242
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _378_
timestamp 1701704242
transform 1 0 14904 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _379_
timestamp 1701704242
transform 1 0 13892 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _380_
timestamp 1701704242
transform 1 0 15364 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _381_
timestamp 1701704242
transform -1 0 14996 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _382_
timestamp 1701704242
transform -1 0 14720 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _383_
timestamp 1701704242
transform -1 0 12788 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _384_
timestamp 1701704242
transform -1 0 14996 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _385_
timestamp 1701704242
transform -1 0 10856 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _386_
timestamp 1701704242
transform 1 0 6256 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _387_
timestamp 1701704242
transform -1 0 6164 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _388_
timestamp 1701704242
transform 1 0 5336 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _389_
timestamp 1701704242
transform 1 0 5152 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _390_
timestamp 1701704242
transform -1 0 6072 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _391_
timestamp 1701704242
transform -1 0 6256 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _392_
timestamp 1701704242
transform -1 0 3772 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _393_
timestamp 1701704242
transform 1 0 2484 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _394_
timestamp 1701704242
transform -1 0 14260 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _395_
timestamp 1701704242
transform 1 0 12788 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _396_
timestamp 1701704242
transform -1 0 14168 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _397_
timestamp 1701704242
transform 1 0 13524 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _398_
timestamp 1701704242
transform -1 0 14168 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _399_
timestamp 1701704242
transform 1 0 10672 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _400_
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _401_
timestamp 1701704242
transform 1 0 14168 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1701704242
transform -1 0 5520 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _403_
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_4  _404_
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1701704242
transform 1 0 19044 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1701704242
transform 1 0 21436 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1701704242
transform 1 0 22540 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1701704242
transform 1 0 22724 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1701704242
transform -1 0 12696 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1701704242
transform -1 0 13800 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1701704242
transform 1 0 9016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1701704242
transform -1 0 8096 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1701704242
transform 1 0 14628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1701704242
transform -1 0 18400 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1701704242
transform -1 0 18584 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1701704242
transform -1 0 16376 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1701704242
transform 1 0 4784 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1701704242
transform 1 0 7360 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1701704242
transform 1 0 3864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1701704242
transform -1 0 4140 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _421_
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1701704242
transform 1 0 20056 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1701704242
transform 1 0 23460 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1701704242
transform 1 0 19504 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1701704242
transform 1 0 22816 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1701704242
transform -1 0 18952 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1701704242
transform -1 0 13064 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1701704242
transform 1 0 9016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1701704242
transform -1 0 9200 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1701704242
transform -1 0 15548 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1701704242
transform -1 0 18952 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1701704242
transform -1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1701704242
transform -1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1701704242
transform 1 0 7912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1701704242
transform 1 0 4324 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1701704242
transform -1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1701704242
transform -1 0 4416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _438_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18492 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _439_
timestamp 1701704242
transform -1 0 21620 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _440_
timestamp 1701704242
transform 1 0 24840 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _441_
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _442_
timestamp 1701704242
transform 1 0 11316 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1701704242
transform 1 0 13248 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _444_
timestamp 1701704242
transform 1 0 9844 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _445_
timestamp 1701704242
transform 1 0 8188 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1701704242
transform 1 0 23368 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _449_
timestamp 1701704242
transform 1 0 21620 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp 1701704242
transform 1 0 6164 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1701704242
transform 1 0 7176 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp 1701704242
transform 1 0 4968 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1701704242
transform 1 0 3404 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1701704242
transform 1 0 19596 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp 1701704242
transform 1 0 23828 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1701704242
transform 1 0 24012 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1701704242
transform 1 0 21252 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1701704242
transform 1 0 16192 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1701704242
transform 1 0 7912 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1701704242
transform 1 0 4232 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1701704242
transform 1 0 11684 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1701704242
transform 1 0 17112 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1701704242
transform 1 0 24840 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _465_
timestamp 1701704242
transform 1 0 21712 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _466_
timestamp 1701704242
transform 1 0 19872 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _467_
timestamp 1701704242
transform 1 0 14076 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _468_
timestamp 1701704242
transform 1 0 9384 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _469_
timestamp 1701704242
transform 1 0 6164 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _470_
timestamp 1701704242
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _471_
timestamp 1701704242
transform 1 0 16376 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _472_
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _473_
timestamp 1701704242
transform 1 0 23184 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1701704242
transform -1 0 23736 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _475_
timestamp 1701704242
transform 1 0 13708 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _476_
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _477_
timestamp 1701704242
transform 1 0 7636 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _478_
timestamp 1701704242
transform 1 0 9384 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _479_
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _480_
timestamp 1701704242
transform -1 0 29348 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _481_
timestamp 1701704242
transform -1 0 27876 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1701704242
transform 1 0 18400 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1701704242
transform 1 0 13524 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1701704242
transform 1 0 8648 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1701704242
transform 1 0 5612 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _486_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18676 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _487_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20608 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1701704242
transform 1 0 21620 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1701704242
transform 1 0 21804 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1701704242
transform 1 0 11316 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 1701704242
transform 1 0 11592 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 1701704242
transform -1 0 10212 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1701704242
transform 1 0 6624 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _494_
timestamp 1701704242
transform 1 0 13616 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1701704242
transform 1 0 16284 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1701704242
transform 1 0 17388 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _497_
timestamp 1701704242
transform 1 0 14996 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _498_
timestamp 1701704242
transform 1 0 3772 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _499_
timestamp 1701704242
transform 1 0 6256 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1701704242
transform -1 0 4048 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1701704242
transform -1 0 14260 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1701704242
transform 1 0 23276 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1701704242
transform 1 0 20332 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1701704242
transform 1 0 23460 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1701704242
transform 1 0 24840 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1701704242
transform 1 0 12144 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1701704242
transform 1 0 10028 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1701704242
transform 1 0 8556 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1701704242
transform 1 0 11776 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1701704242
transform 1 0 21804 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1701704242
transform 1 0 18676 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _513_
timestamp 1701704242
transform 1 0 16836 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _514_
timestamp 1701704242
transform 1 0 19412 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _515_
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _516_
timestamp 1701704242
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _517_
timestamp 1701704242
transform 1 0 5060 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _518_
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _519_
timestamp 1701704242
transform 1 0 23092 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _520_
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _521_
timestamp 1701704242
transform 1 0 24288 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _522_
timestamp 1701704242
transform 1 0 20056 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _523_
timestamp 1701704242
transform 1 0 16652 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _524_
timestamp 1701704242
transform 1 0 17112 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _525_
timestamp 1701704242
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _526_
timestamp 1701704242
transform 1 0 11960 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _527_
timestamp 1701704242
transform 1 0 28428 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _528_
timestamp 1701704242
transform 1 0 26588 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _529_
timestamp 1701704242
transform 1 0 28060 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _530_
timestamp 1701704242
transform 1 0 27232 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _531_
timestamp 1701704242
transform 1 0 13248 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _532_
timestamp 1701704242
transform 1 0 18400 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _533_
timestamp 1701704242
transform 1 0 7636 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _534_
timestamp 1701704242
transform 1 0 7268 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _535_
timestamp 1701704242
transform 1 0 24104 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _536_
timestamp 1701704242
transform -1 0 22724 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _537_
timestamp 1701704242
transform 1 0 24012 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _538_
timestamp 1701704242
transform 1 0 24748 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _539_
timestamp 1701704242
transform 1 0 14812 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _540_
timestamp 1701704242
transform 1 0 10764 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _541_
timestamp 1701704242
transform 1 0 8832 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _542_
timestamp 1701704242
transform 1 0 11592 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _543_
timestamp 1701704242
transform 1 0 28980 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _544_
timestamp 1701704242
transform 1 0 28060 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _545_
timestamp 1701704242
transform 1 0 28980 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _546_
timestamp 1701704242
transform 1 0 27324 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _547_
timestamp 1701704242
transform 1 0 15272 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _548_
timestamp 1701704242
transform 1 0 8740 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _549_
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _550_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 19044 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _551_
timestamp 1701704242
transform 1 0 21528 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _552_
timestamp 1701704242
transform 1 0 18584 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _553_
timestamp 1701704242
transform 1 0 21896 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _554_
timestamp 1701704242
transform 1 0 16652 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _555_
timestamp 1701704242
transform 1 0 10948 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _556_
timestamp 1701704242
transform 1 0 8096 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _557_
timestamp 1701704242
transform 1 0 6440 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _558_
timestamp 1701704242
transform 1 0 13340 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _559_
timestamp 1701704242
transform 1 0 16468 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _560_
timestamp 1701704242
transform 1 0 16652 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _561_
timestamp 1701704242
transform 1 0 14720 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _562_
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _563_
timestamp 1701704242
transform 1 0 3312 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _564_
timestamp 1701704242
transform 1 0 3312 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _565_
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _620_
timestamp 1701704242
transform -1 0 3680 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _621_
timestamp 1701704242
transform -1 0 3312 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _622_
timestamp 1701704242
transform -1 0 3128 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _623_
timestamp 1701704242
transform -1 0 4876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 20332 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  fanout7
timestamp 1701704242
transform -1 0 7268 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout8
timestamp 1701704242
transform 1 0 14996 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout9
timestamp 1701704242
transform 1 0 18032 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout10
timestamp 1701704242
transform -1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1701704242
transform -1 0 9568 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1701704242
transform -1 0 15088 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1701704242
transform -1 0 27324 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1701704242
transform 1 0 26588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1701704242
transform -1 0 27876 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1701704242
transform -1 0 3864 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1701704242
transform -1 0 3772 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1701704242
transform 1 0 19228 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1701704242
transform 1 0 13708 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1701704242
transform 1 0 3772 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1701704242
transform -1 0 3404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1701704242
transform -1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1701704242
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1701704242
transform -1 0 10212 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1701704242
transform -1 0 12052 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1701704242
transform 1 0 17296 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1701704242
transform -1 0 17388 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 1701704242
transform -1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1701704242
transform -1 0 24564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1701704242
transform -1 0 23368 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1701704242
transform 1 0 23644 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1701704242
transform -1 0 16928 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 1701704242
transform -1 0 17664 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1701704242
transform 1 0 27324 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1701704242
transform 1 0 26956 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_68
timestamp 1701704242
transform 1 0 6808 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_80 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7912 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1701704242
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_152
timestamp 1701704242
transform 1 0 14536 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_160
timestamp 1701704242
transform 1 0 15272 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15824 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_173
timestamp 1701704242
transform 1 0 16468 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_180
timestamp 1701704242
transform 1 0 17112 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_192
timestamp 1701704242
transform 1 0 18216 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_201
timestamp 1701704242
transform 1 0 19044 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_213
timestamp 1701704242
transform 1 0 20148 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1701704242
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1701704242
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1701704242
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1701704242
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_329
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1701704242
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1701704242
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1701704242
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1701704242
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1701704242
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1701704242
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1701704242
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1701704242
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1701704242
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1701704242
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1701704242
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1701704242
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1701704242
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1701704242
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1701704242
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1701704242
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1701704242
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1701704242
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1701704242
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1701704242
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1701704242
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1701704242
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1701704242
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1701704242
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_91
timestamp 1701704242
transform 1 0 8924 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_95
timestamp 1701704242
transform 1 0 9292 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_107
timestamp 1701704242
transform 1 0 10396 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1701704242
transform 1 0 13064 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_165
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_173
timestamp 1701704242
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_200
timestamp 1701704242
transform 1 0 18952 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_215
timestamp 1701704242
transform 1 0 20332 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_226
timestamp 1701704242
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_238
timestamp 1701704242
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1701704242
transform 1 0 23552 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1701704242
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1701704242
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1701704242
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1701704242
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1701704242
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1701704242
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_329
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_102
timestamp 1701704242
transform 1 0 9936 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1701704242
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_121
timestamp 1701704242
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_127
timestamp 1701704242
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_131
timestamp 1701704242
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_163
timestamp 1701704242
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_176
timestamp 1701704242
transform 1 0 16744 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_188
timestamp 1701704242
transform 1 0 17848 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_196
timestamp 1701704242
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21252 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_252
timestamp 1701704242
transform 1 0 23736 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_264
timestamp 1701704242
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_276
timestamp 1701704242
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1701704242
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1701704242
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1701704242
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1701704242
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_61
timestamp 1701704242
transform 1 0 6164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_94
timestamp 1701704242
transform 1 0 9200 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_103
timestamp 1701704242
transform 1 0 10028 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_119
timestamp 1701704242
transform 1 0 11500 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1701704242
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1701704242
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_153
timestamp 1701704242
transform 1 0 14628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_166
timestamp 1701704242
transform 1 0 15824 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_172
timestamp 1701704242
transform 1 0 16376 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1701704242
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_200
timestamp 1701704242
transform 1 0 18952 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_222
timestamp 1701704242
transform 1 0 20976 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_230
timestamp 1701704242
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_253
timestamp 1701704242
transform 1 0 23828 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_261
timestamp 1701704242
transform 1 0 24564 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_280
timestamp 1701704242
transform 1 0 26312 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_292
timestamp 1701704242
transform 1 0 27416 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_304
timestamp 1701704242
transform 1 0 28520 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1701704242
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_329
timestamp 1701704242
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_44
timestamp 1701704242
transform 1 0 4600 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_98
timestamp 1701704242
transform 1 0 9568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_118
timestamp 1701704242
transform 1 0 11408 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_142
timestamp 1701704242
transform 1 0 13616 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_157
timestamp 1701704242
transform 1 0 14996 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_195
timestamp 1701704242
transform 1 0 18492 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_216
timestamp 1701704242
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1701704242
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_245
timestamp 1701704242
transform 1 0 23092 0 -1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_265
timestamp 1701704242
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1701704242
transform 1 0 26036 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1701704242
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1701704242
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_329
timestamp 1701704242
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_50
timestamp 1701704242
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_61
timestamp 1701704242
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_73
timestamp 1701704242
transform 1 0 7268 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_79
timestamp 1701704242
transform 1 0 7820 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_119
timestamp 1701704242
transform 1 0 11500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1701704242
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_141
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_174
timestamp 1701704242
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_186
timestamp 1701704242
transform 1 0 17664 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_190
timestamp 1701704242
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_213
timestamp 1701704242
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_231
timestamp 1701704242
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_243
timestamp 1701704242
transform 1 0 22908 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1701704242
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1701704242
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1701704242
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_277
timestamp 1701704242
transform 1 0 26036 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_298
timestamp 1701704242
transform 1 0 27968 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_306
timestamp 1701704242
transform 1 0 28704 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 1701704242
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_329
timestamp 1701704242
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_31
timestamp 1701704242
transform 1 0 3404 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_35
timestamp 1701704242
transform 1 0 3772 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_47
timestamp 1701704242
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_62
timestamp 1701704242
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_74
timestamp 1701704242
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_86
timestamp 1701704242
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_98
timestamp 1701704242
transform 1 0 9568 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1701704242
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_125
timestamp 1701704242
transform 1 0 12052 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_149
timestamp 1701704242
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1701704242
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1701704242
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_172
timestamp 1701704242
transform 1 0 16376 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_176
timestamp 1701704242
transform 1 0 16744 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1701704242
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1701704242
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_225
timestamp 1701704242
transform 1 0 21252 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1701704242
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_281
timestamp 1701704242
transform 1 0 26404 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_287
timestamp 1701704242
transform 1 0 26956 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_307
timestamp 1701704242
transform 1 0 28796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_319
timestamp 1701704242
transform 1 0 29900 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_331
timestamp 1701704242
transform 1 0 31004 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_60
timestamp 1701704242
transform 1 0 6072 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_105
timestamp 1701704242
transform 1 0 10212 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_134
timestamp 1701704242
transform 1 0 12880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_144
timestamp 1701704242
transform 1 0 13800 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_155
timestamp 1701704242
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_176
timestamp 1701704242
transform 1 0 16744 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_188
timestamp 1701704242
transform 1 0 17848 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_205
timestamp 1701704242
transform 1 0 19412 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_211
timestamp 1701704242
transform 1 0 19964 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_228
timestamp 1701704242
transform 1 0 21528 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_236
timestamp 1701704242
transform 1 0 22264 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_263
timestamp 1701704242
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_275
timestamp 1701704242
transform 1 0 25852 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_292
timestamp 1701704242
transform 1 0 27416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_304
timestamp 1701704242
transform 1 0 28520 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_321
timestamp 1701704242
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 1701704242
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_42
timestamp 1701704242
transform 1 0 4416 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1701704242
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_73
timestamp 1701704242
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_92
timestamp 1701704242
transform 1 0 9016 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_104
timestamp 1701704242
transform 1 0 10120 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_119
timestamp 1701704242
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_126
timestamp 1701704242
transform 1 0 12144 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_137
timestamp 1701704242
transform 1 0 13156 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1701704242
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1701704242
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_177
timestamp 1701704242
transform 1 0 16836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_210
timestamp 1701704242
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_215
timestamp 1701704242
transform 1 0 20332 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_225
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_229
timestamp 1701704242
transform 1 0 21620 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_253
timestamp 1701704242
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_271
timestamp 1701704242
transform 1 0 25484 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_281
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_314
timestamp 1701704242
transform 1 0 29440 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_326
timestamp 1701704242
transform 1 0 30544 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_15
timestamp 1701704242
transform 1 0 1932 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_65
timestamp 1701704242
transform 1 0 6532 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_72
timestamp 1701704242
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1701704242
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_114
timestamp 1701704242
transform 1 0 11040 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_118
timestamp 1701704242
transform 1 0 11408 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_125
timestamp 1701704242
transform 1 0 12052 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_137
timestamp 1701704242
transform 1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_149
timestamp 1701704242
transform 1 0 14260 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_171
timestamp 1701704242
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1701704242
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_200
timestamp 1701704242
transform 1 0 18952 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_212
timestamp 1701704242
transform 1 0 20056 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_224
timestamp 1701704242
transform 1 0 21160 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1701704242
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_245
timestamp 1701704242
transform 1 0 23092 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1701704242
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_260
timestamp 1701704242
transform 1 0 24472 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_264
timestamp 1701704242
transform 1 0 24840 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_273
timestamp 1701704242
transform 1 0 25668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_287
timestamp 1701704242
transform 1 0 26956 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_303
timestamp 1701704242
transform 1 0 28428 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1701704242
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_325
timestamp 1701704242
transform 1 0 30452 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_331
timestamp 1701704242
transform 1 0 31004 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1701704242
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_39
timestamp 1701704242
transform 1 0 4140 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_47
timestamp 1701704242
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1701704242
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_75
timestamp 1701704242
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_93
timestamp 1701704242
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_97
timestamp 1701704242
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1701704242
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_123
timestamp 1701704242
transform 1 0 11868 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_148
timestamp 1701704242
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_156
timestamp 1701704242
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1701704242
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_189
timestamp 1701704242
transform 1 0 17940 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_219
timestamp 1701704242
transform 1 0 20700 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1701704242
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_241
timestamp 1701704242
transform 1 0 22724 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_274
timestamp 1701704242
transform 1 0 25760 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_45
timestamp 1701704242
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_51
timestamp 1701704242
transform 1 0 5244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_76
timestamp 1701704242
transform 1 0 7544 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_89
timestamp 1701704242
transform 1 0 8740 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_106
timestamp 1701704242
transform 1 0 10304 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1701704242
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1701704242
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_152
timestamp 1701704242
transform 1 0 14536 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_158
timestamp 1701704242
transform 1 0 15088 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_178
timestamp 1701704242
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_205
timestamp 1701704242
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_212
timestamp 1701704242
transform 1 0 20056 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_220
timestamp 1701704242
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_225
timestamp 1701704242
transform 1 0 21252 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_237
timestamp 1701704242
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1701704242
transform 1 0 23552 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_260
timestamp 1701704242
transform 1 0 24472 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_268
timestamp 1701704242
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_277
timestamp 1701704242
transform 1 0 26036 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_304
timestamp 1701704242
transform 1 0 28520 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_325
timestamp 1701704242
transform 1 0 30452 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_331
timestamp 1701704242
transform 1 0 31004 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_23
timestamp 1701704242
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_34
timestamp 1701704242
transform 1 0 3680 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_65
timestamp 1701704242
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_89
timestamp 1701704242
transform 1 0 8740 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_95
timestamp 1701704242
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_99
timestamp 1701704242
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1701704242
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_119
timestamp 1701704242
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_131
timestamp 1701704242
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_140
timestamp 1701704242
transform 1 0 13432 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_163
timestamp 1701704242
transform 1 0 15548 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1701704242
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_189
timestamp 1701704242
transform 1 0 17940 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_211
timestamp 1701704242
transform 1 0 19964 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_218
timestamp 1701704242
transform 1 0 20608 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_241
timestamp 1701704242
transform 1 0 22724 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_246
timestamp 1701704242
transform 1 0 23184 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1701704242
transform 1 0 26128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_281
timestamp 1701704242
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_301
timestamp 1701704242
transform 1 0 28244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_326
timestamp 1701704242
transform 1 0 30544 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_54
timestamp 1701704242
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_65
timestamp 1701704242
transform 1 0 6532 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_74
timestamp 1701704242
transform 1 0 7360 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1701704242
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_93
timestamp 1701704242
transform 1 0 9108 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_117
timestamp 1701704242
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1701704242
transform 1 0 13064 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_155
timestamp 1701704242
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_159
timestamp 1701704242
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_174
timestamp 1701704242
transform 1 0 16560 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1701704242
transform 1 0 18124 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1701704242
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1701704242
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_209
timestamp 1701704242
transform 1 0 19780 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_218
timestamp 1701704242
transform 1 0 20608 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_226
timestamp 1701704242
transform 1 0 21344 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_242
timestamp 1701704242
transform 1 0 22816 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 1701704242
transform 1 0 23368 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1701704242
transform 1 0 23828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_265
timestamp 1701704242
transform 1 0 24932 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_273
timestamp 1701704242
transform 1 0 25668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_281
timestamp 1701704242
transform 1 0 26404 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_291
timestamp 1701704242
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_295
timestamp 1701704242
transform 1 0 27692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_300
timestamp 1701704242
transform 1 0 28152 0 1 9248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_316
timestamp 1701704242
transform 1 0 29624 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_328
timestamp 1701704242
transform 1 0 30728 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_31
timestamp 1701704242
transform 1 0 3404 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_39
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_93
timestamp 1701704242
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1701704242
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_118
timestamp 1701704242
transform 1 0 11408 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_136
timestamp 1701704242
transform 1 0 13064 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_144
timestamp 1701704242
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_152
timestamp 1701704242
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_160
timestamp 1701704242
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_195
timestamp 1701704242
transform 1 0 18492 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_201
timestamp 1701704242
transform 1 0 19044 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_210
timestamp 1701704242
transform 1 0 19872 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_214
timestamp 1701704242
transform 1 0 20240 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_217
timestamp 1701704242
transform 1 0 20516 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_241
timestamp 1701704242
transform 1 0 22724 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_261
timestamp 1701704242
transform 1 0 24564 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1701704242
transform 1 0 26128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_315
timestamp 1701704242
transform 1 0 29532 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_327
timestamp 1701704242
transform 1 0 30636 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_331
timestamp 1701704242
transform 1 0 31004 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_6
timestamp 1701704242
transform 1 0 1104 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_18
timestamp 1701704242
transform 1 0 2208 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1701704242
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_47
timestamp 1701704242
transform 1 0 4876 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_51
timestamp 1701704242
transform 1 0 5244 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_71
timestamp 1701704242
transform 1 0 7084 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_77
timestamp 1701704242
transform 1 0 7636 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1701704242
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_97
timestamp 1701704242
transform 1 0 9476 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_108
timestamp 1701704242
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_117
timestamp 1701704242
transform 1 0 11316 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1701704242
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_153
timestamp 1701704242
transform 1 0 14628 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_168
timestamp 1701704242
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_173
timestamp 1701704242
transform 1 0 16468 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_185
timestamp 1701704242
transform 1 0 17572 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1701704242
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_213
timestamp 1701704242
transform 1 0 20148 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_222
timestamp 1701704242
transform 1 0 20976 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_233
timestamp 1701704242
transform 1 0 21988 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_265
timestamp 1701704242
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_281
timestamp 1701704242
transform 1 0 26404 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_293
timestamp 1701704242
transform 1 0 27508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1701704242
transform 1 0 28612 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_321
timestamp 1701704242
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_329
timestamp 1701704242
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_38
timestamp 1701704242
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_46
timestamp 1701704242
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1701704242
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1701704242
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_60
timestamp 1701704242
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_72
timestamp 1701704242
transform 1 0 7176 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_92
timestamp 1701704242
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_120
timestamp 1701704242
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_125
timestamp 1701704242
transform 1 0 12052 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_129
timestamp 1701704242
transform 1 0 12420 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_136
timestamp 1701704242
transform 1 0 13064 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1701704242
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1701704242
transform 1 0 16100 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_187
timestamp 1701704242
transform 1 0 17756 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_213
timestamp 1701704242
transform 1 0 20148 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1701704242
transform 1 0 20516 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1701704242
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_225
timestamp 1701704242
transform 1 0 21252 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_233
timestamp 1701704242
transform 1 0 21988 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_248
timestamp 1701704242
transform 1 0 23368 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1701704242
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_297
timestamp 1701704242
transform 1 0 27876 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_309
timestamp 1701704242
transform 1 0 28980 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_321
timestamp 1701704242
transform 1 0 30084 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_329
timestamp 1701704242
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1701704242
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_39
timestamp 1701704242
transform 1 0 4140 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_43
timestamp 1701704242
transform 1 0 4508 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_63
timestamp 1701704242
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_70
timestamp 1701704242
transform 1 0 6992 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_74
timestamp 1701704242
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_91
timestamp 1701704242
transform 1 0 8924 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_103
timestamp 1701704242
transform 1 0 10028 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_111
timestamp 1701704242
transform 1 0 10764 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_126
timestamp 1701704242
transform 1 0 12144 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_130
timestamp 1701704242
transform 1 0 12512 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_148
timestamp 1701704242
transform 1 0 14168 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_156
timestamp 1701704242
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1701704242
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_177
timestamp 1701704242
transform 1 0 16836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_181
timestamp 1701704242
transform 1 0 17204 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_190
timestamp 1701704242
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1701704242
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_200
timestamp 1701704242
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_205
timestamp 1701704242
transform 1 0 19412 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_229
timestamp 1701704242
transform 1 0 21620 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1701704242
transform 1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_256
timestamp 1701704242
transform 1 0 24104 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_268
timestamp 1701704242
transform 1 0 25208 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_291
timestamp 1701704242
transform 1 0 27324 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_296
timestamp 1701704242
transform 1 0 27784 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1701704242
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_329
timestamp 1701704242
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_43
timestamp 1701704242
transform 1 0 4508 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1701704242
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_61
timestamp 1701704242
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_116
timestamp 1701704242
transform 1 0 11224 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_136
timestamp 1701704242
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_146
timestamp 1701704242
transform 1 0 13984 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_163
timestamp 1701704242
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_180
timestamp 1701704242
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_194
timestamp 1701704242
transform 1 0 18400 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_206
timestamp 1701704242
transform 1 0 19504 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_212
timestamp 1701704242
transform 1 0 20056 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_236
timestamp 1701704242
transform 1 0 22264 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_252
timestamp 1701704242
transform 1 0 23736 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_313
timestamp 1701704242
transform 1 0 29348 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_325
timestamp 1701704242
transform 1 0 30452 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_331
timestamp 1701704242
transform 1 0 31004 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_23
timestamp 1701704242
transform 1 0 2668 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_49
timestamp 1701704242
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_60
timestamp 1701704242
transform 1 0 6072 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1701704242
transform 1 0 7912 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_90
timestamp 1701704242
transform 1 0 8832 0 1 12512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_101
timestamp 1701704242
transform 1 0 9844 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_113
timestamp 1701704242
transform 1 0 10948 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_117
timestamp 1701704242
transform 1 0 11316 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_126
timestamp 1701704242
transform 1 0 12144 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1701704242
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1701704242
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_149
timestamp 1701704242
transform 1 0 14260 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_156
timestamp 1701704242
transform 1 0 14904 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_178
timestamp 1701704242
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_197
timestamp 1701704242
transform 1 0 18676 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_203
timestamp 1701704242
transform 1 0 19228 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_233
timestamp 1701704242
transform 1 0 21988 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_239
timestamp 1701704242
transform 1 0 22540 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_243
timestamp 1701704242
transform 1 0 22908 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1701704242
transform 1 0 23552 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_253
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_261
timestamp 1701704242
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_266
timestamp 1701704242
transform 1 0 25024 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_278
timestamp 1701704242
transform 1 0 26128 0 1 12512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_294
timestamp 1701704242
transform 1 0 27600 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_306
timestamp 1701704242
transform 1 0 28704 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 1701704242
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_15
timestamp 1701704242
transform 1 0 1932 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_23
timestamp 1701704242
transform 1 0 2668 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_27
timestamp 1701704242
transform 1 0 3036 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_42
timestamp 1701704242
transform 1 0 4416 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_50
timestamp 1701704242
transform 1 0 5152 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1701704242
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_60
timestamp 1701704242
transform 1 0 6072 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_69
timestamp 1701704242
transform 1 0 6900 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1701704242
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_139
timestamp 1701704242
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_164
timestamp 1701704242
transform 1 0 15640 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_188
timestamp 1701704242
transform 1 0 17848 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_196
timestamp 1701704242
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_205
timestamp 1701704242
transform 1 0 19412 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_221
timestamp 1701704242
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_225
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_229
timestamp 1701704242
transform 1 0 21620 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_262
timestamp 1701704242
transform 1 0 24656 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_288
timestamp 1701704242
transform 1 0 27048 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_300
timestamp 1701704242
transform 1 0 28152 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_312
timestamp 1701704242
transform 1 0 29256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_324
timestamp 1701704242
transform 1 0 30360 0 -1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1701704242
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_46
timestamp 1701704242
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_70
timestamp 1701704242
transform 1 0 6992 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1701704242
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1701704242
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_97
timestamp 1701704242
transform 1 0 9476 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_117
timestamp 1701704242
transform 1 0 11316 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_129
timestamp 1701704242
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1701704242
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_177
timestamp 1701704242
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1701704242
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1701704242
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1701704242
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_253
timestamp 1701704242
transform 1 0 23828 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_261
timestamp 1701704242
transform 1 0 24564 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_270
timestamp 1701704242
transform 1 0 25392 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_282
timestamp 1701704242
transform 1 0 26496 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_294
timestamp 1701704242
transform 1 0 27600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1701704242
transform 1 0 28704 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 1701704242
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_329
timestamp 1701704242
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_6
timestamp 1701704242
transform 1 0 1104 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_18
timestamp 1701704242
transform 1 0 2208 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_29
timestamp 1701704242
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_38
timestamp 1701704242
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_49
timestamp 1701704242
transform 1 0 5060 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_82
timestamp 1701704242
transform 1 0 8096 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_99
timestamp 1701704242
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1701704242
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1701704242
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_133
timestamp 1701704242
transform 1 0 12788 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_137
timestamp 1701704242
transform 1 0 13156 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_154
timestamp 1701704242
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1701704242
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_176
timestamp 1701704242
transform 1 0 16744 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_203
timestamp 1701704242
transform 1 0 19228 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_215
timestamp 1701704242
transform 1 0 20332 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1701704242
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1701704242
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_237
timestamp 1701704242
transform 1 0 22356 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_242
timestamp 1701704242
transform 1 0 22816 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1701704242
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1701704242
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1701704242
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_329
timestamp 1701704242
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1701704242
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1701704242
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_56
timestamp 1701704242
transform 1 0 5704 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_60
timestamp 1701704242
transform 1 0 6072 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_67
timestamp 1701704242
transform 1 0 6716 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1701704242
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_114
timestamp 1701704242
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_144
timestamp 1701704242
transform 1 0 13800 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_152
timestamp 1701704242
transform 1 0 14536 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_170
timestamp 1701704242
transform 1 0 16192 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_185
timestamp 1701704242
transform 1 0 17572 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_207
timestamp 1701704242
transform 1 0 19596 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_227
timestamp 1701704242
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 1701704242
transform 1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_269
timestamp 1701704242
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_281
timestamp 1701704242
transform 1 0 26404 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_293
timestamp 1701704242
transform 1 0 27508 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_305
timestamp 1701704242
transform 1 0 28612 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1701704242
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1701704242
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_65
timestamp 1701704242
transform 1 0 6532 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_94
timestamp 1701704242
transform 1 0 9200 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_102
timestamp 1701704242
transform 1 0 9936 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_124
timestamp 1701704242
transform 1 0 11960 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_136
timestamp 1701704242
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_148
timestamp 1701704242
transform 1 0 14168 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_152
timestamp 1701704242
transform 1 0 14536 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_156
timestamp 1701704242
transform 1 0 14904 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1701704242
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 1701704242
transform 1 0 17204 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_189
timestamp 1701704242
transform 1 0 17940 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_194
timestamp 1701704242
transform 1 0 18400 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_200
timestamp 1701704242
transform 1 0 18952 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_204
timestamp 1701704242
transform 1 0 19320 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_215
timestamp 1701704242
transform 1 0 20332 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_228
timestamp 1701704242
transform 1 0 21528 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_255
timestamp 1701704242
transform 1 0 24012 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_267
timestamp 1701704242
transform 1 0 25116 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1701704242
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1701704242
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1701704242
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1701704242
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1701704242
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_329
timestamp 1701704242
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1701704242
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1701704242
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1701704242
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1701704242
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_108
timestamp 1701704242
transform 1 0 10488 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_118
timestamp 1701704242
transform 1 0 11408 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_126
timestamp 1701704242
transform 1 0 12144 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_132
timestamp 1701704242
transform 1 0 12696 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_163
timestamp 1701704242
transform 1 0 15548 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1701704242
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_238
timestamp 1701704242
transform 1 0 22448 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_244
timestamp 1701704242
transform 1 0 23000 0 1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1701704242
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1701704242
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1701704242
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1701704242
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1701704242
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1701704242
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1701704242
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1701704242
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1701704242
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1701704242
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1701704242
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1701704242
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1701704242
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_81
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_89
timestamp 1701704242
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_95
timestamp 1701704242
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_101
timestamp 1701704242
transform 1 0 9844 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1701704242
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_189
timestamp 1701704242
transform 1 0 17940 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_194
timestamp 1701704242
transform 1 0 18400 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_206
timestamp 1701704242
transform 1 0 19504 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_218
timestamp 1701704242
transform 1 0 20608 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_225
timestamp 1701704242
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_230
timestamp 1701704242
transform 1 0 21712 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_242
timestamp 1701704242
transform 1 0 22816 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_254
timestamp 1701704242
transform 1 0 23920 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_266
timestamp 1701704242
transform 1 0 25024 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1701704242
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1701704242
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1701704242
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1701704242
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1701704242
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1701704242
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1701704242
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1701704242
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1701704242
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1701704242
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1701704242
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1701704242
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1701704242
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1701704242
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1701704242
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1701704242
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1701704242
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1701704242
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1701704242
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1701704242
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1701704242
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1701704242
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1701704242
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1701704242
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1701704242
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1701704242
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1701704242
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1701704242
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1701704242
transform 1 0 20516 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1701704242
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1701704242
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1701704242
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1701704242
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1701704242
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1701704242
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1701704242
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1701704242
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1701704242
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1701704242
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1701704242
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1701704242
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1701704242
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1701704242
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1701704242
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1701704242
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1701704242
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1701704242
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1701704242
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_105
timestamp 1701704242
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 1701704242
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_117
timestamp 1701704242
transform 1 0 11316 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_131
timestamp 1701704242
transform 1 0 12604 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_138
timestamp 1701704242
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_153
timestamp 1701704242
transform 1 0 14628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_173
timestamp 1701704242
transform 1 0 16468 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_185
timestamp 1701704242
transform 1 0 17572 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_194
timestamp 1701704242
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_201
timestamp 1701704242
transform 1 0 19044 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_208
timestamp 1701704242
transform 1 0 19688 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_215
timestamp 1701704242
transform 1 0 20332 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1701704242
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_229
timestamp 1701704242
transform 1 0 21620 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_236
timestamp 1701704242
transform 1 0 22264 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_248
timestamp 1701704242
transform 1 0 23368 0 -1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1701704242
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1701704242
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_305
timestamp 1701704242
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 31096 0 -1 8160
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1701704242
transform -1 0 17112 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1701704242
transform 1 0 16192 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1701704242
transform 1 0 15548 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap11
timestamp 1701704242
transform 1 0 5244 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap12
timestamp 1701704242
transform 1 0 19228 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap13
timestamp 1701704242
transform -1 0 8096 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap14
timestamp 1701704242
transform 1 0 12512 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap25
timestamp 1701704242
transform -1 0 16008 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  tdc0.g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[0\].dly_stp
timestamp 1701704242
transform -1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[1\].dly_stp
timestamp 1701704242
transform -1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[2\].dly_stp
timestamp 1701704242
transform -1 0 3036 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[3\].dly_stp
timestamp 1701704242
transform -1 0 3128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[4\].dly_stp
timestamp 1701704242
transform -1 0 3404 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[1\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 19596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[1\].stg01
timestamp 1701704242
transform 1 0 16560 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[1\].stg02 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16192 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[2\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 24104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[2\].stg01
timestamp 1701704242
transform -1 0 22540 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[2\].stg02
timestamp 1701704242
transform -1 0 22816 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[3\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 24012 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[3\].stg01
timestamp 1701704242
transform 1 0 23184 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[3\].stg02
timestamp 1701704242
transform 1 0 22724 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[4\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 20976 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[4\].stg01
timestamp 1701704242
transform 1 0 23092 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[4\].stg02
timestamp 1701704242
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[5\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 16468 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[5\].stg01
timestamp 1701704242
transform 1 0 17204 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[5\].stg02
timestamp 1701704242
transform 1 0 16192 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[6\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[6\].stg01
timestamp 1701704242
transform 1 0 11776 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[6\].stg02
timestamp 1701704242
transform -1 0 12144 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[7\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 4968 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[7\].stg01
timestamp 1701704242
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[7\].stg02
timestamp 1701704242
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[8\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[8\].stg01
timestamp 1701704242
transform -1 0 9016 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[8\].stg02
timestamp 1701704242
transform 1 0 8004 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[9\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 17848 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[9\].stg01
timestamp 1701704242
transform -1 0 13064 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[9\].stg02
timestamp 1701704242
transform -1 0 17664 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[10\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 25024 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[10\].stg01
timestamp 1701704242
transform -1 0 18400 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[10\].stg02
timestamp 1701704242
transform -1 0 19228 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[11\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 21988 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[11\].stg01
timestamp 1701704242
transform -1 0 21160 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[11\].stg02
timestamp 1701704242
transform -1 0 21620 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[12\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 20148 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[12\].stg01
timestamp 1701704242
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[12\].stg02
timestamp 1701704242
transform 1 0 19688 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[13\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 14628 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[13\].stg01
timestamp 1701704242
transform 1 0 19136 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[13\].stg02
timestamp 1701704242
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[14\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 9568 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[14\].stg01
timestamp 1701704242
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[14\].stg02
timestamp 1701704242
transform 1 0 12696 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[15\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 6716 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[15\].stg01
timestamp 1701704242
transform 1 0 7636 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[15\].stg02
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[16\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[16\].stg01
timestamp 1701704242
transform -1 0 6900 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring1\[16\].stg02_42 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[16\].stg02
timestamp 1701704242
transform 1 0 4876 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[16\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 4968 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[16\].stg01_43
timestamp 1701704242
transform -1 0 6900 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[16\].stg01
timestamp 1701704242
transform -1 0 6624 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[16\].stg02
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[17\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 15732 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[17\].stg01_44
timestamp 1701704242
transform -1 0 5520 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[17\].stg01
timestamp 1701704242
transform -1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[17\].stg02
timestamp 1701704242
transform -1 0 16376 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[18\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 26312 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[18\].stg01_45
timestamp 1701704242
transform 1 0 15732 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[18\].stg01
timestamp 1701704242
transform -1 0 17112 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[18\].stg02
timestamp 1701704242
transform -1 0 23184 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[19\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 23552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[19\].stg01_46
timestamp 1701704242
transform 1 0 23000 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[19\].stg01
timestamp 1701704242
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[19\].stg02
timestamp 1701704242
transform 1 0 23092 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[20\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 23092 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[20\].stg01
timestamp 1701704242
transform 1 0 22448 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[20\].stg01_47
timestamp 1701704242
transform 1 0 22172 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[20\].stg02
timestamp 1701704242
transform -1 0 22816 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[21\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 13708 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[21\].stg01_48
timestamp 1701704242
transform -1 0 17756 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[21\].stg01
timestamp 1701704242
transform 1 0 16928 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[21\].stg02
timestamp 1701704242
transform 1 0 16560 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[22\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 11224 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[22\].stg01_49
timestamp 1701704242
transform -1 0 13432 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[22\].stg01
timestamp 1701704242
transform 1 0 12512 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[22\].stg02
timestamp 1701704242
transform 1 0 11224 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[23\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[23\].stg01_50
timestamp 1701704242
transform -1 0 10028 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[23\].stg01
timestamp 1701704242
transform 1 0 9476 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[23\].stg02
timestamp 1701704242
transform 1 0 7636 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[24\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 9384 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[24\].stg01_51
timestamp 1701704242
transform -1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[24\].stg01
timestamp 1701704242
transform -1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[24\].stg02
timestamp 1701704242
transform -1 0 8740 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[25\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 18124 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[25\].stg01_52
timestamp 1701704242
transform -1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[25\].stg01
timestamp 1701704242
transform -1 0 12880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[25\].stg02
timestamp 1701704242
transform -1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[26\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 27784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[26\].stg01
timestamp 1701704242
transform -1 0 18400 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[26\].stg01_53
timestamp 1701704242
transform -1 0 18952 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[26\].stg02
timestamp 1701704242
transform -1 0 18860 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[27\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 26220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[27\].stg01
timestamp 1701704242
transform 1 0 21988 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[27\].stg01_54
timestamp 1701704242
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[27\].stg02
timestamp 1701704242
transform 1 0 21620 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[28\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 18400 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[28\].stg01_55
timestamp 1701704242
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[28\].stg01
timestamp 1701704242
transform 1 0 20240 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[28\].stg02
timestamp 1701704242
transform 1 0 19504 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[29\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 14352 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[29\].stg01_56
timestamp 1701704242
transform -1 0 17848 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[29\].stg01
timestamp 1701704242
transform 1 0 17296 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[29\].stg02
timestamp 1701704242
transform 1 0 13616 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[30\].g_buf1.ctr_buf
timestamp 1701704242
transform -1 0 8832 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[30\].stg01_57
timestamp 1701704242
transform -1 0 13340 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[30\].stg01
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[30\].stg02
timestamp 1701704242
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[31\].g_buf1.ctr_buf
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[31\].stg01_58
timestamp 1701704242
transform -1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[31\].stg01
timestamp 1701704242
transform -1 0 7728 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[31\].stg02
timestamp 1701704242
transform 1 0 7268 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tdc0.stg01_59
timestamp 1701704242
transform -1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.stg01
timestamp 1701704242
transform 1 0 5520 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.stg02
timestamp 1701704242
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  tdc1.g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 5520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[0\].dly_stp
timestamp 1701704242
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[1\].dly_stp
timestamp 1701704242
transform -1 0 27140 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[2\].dly_stp
timestamp 1701704242
transform 1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[3\].dly_stp
timestamp 1701704242
transform -1 0 27416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  tdc1.g_dly_stp\[4\].dly_stp
timestamp 1701704242
transform -1 0 27968 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[1\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[1\].stg01
timestamp 1701704242
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[1\].stg02
timestamp 1701704242
transform -1 0 23184 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[2\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 21252 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[2\].stg01
timestamp 1701704242
transform -1 0 23184 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[2\].stg02
timestamp 1701704242
transform -1 0 23552 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[3\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 24472 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[3\].stg01
timestamp 1701704242
transform 1 0 23736 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[3\].stg02
timestamp 1701704242
transform 1 0 23276 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[4\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 20332 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[4\].stg01
timestamp 1701704242
transform 1 0 23552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[4\].stg02
timestamp 1701704242
transform 1 0 22816 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[5\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 17664 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[5\].stg01
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[5\].stg02
timestamp 1701704242
transform 1 0 17756 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[6\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[6\].stg01
timestamp 1701704242
transform -1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[6\].stg02
timestamp 1701704242
transform 1 0 16744 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[7\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 4968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[7\].stg01
timestamp 1701704242
transform 1 0 16468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[7\].stg02
timestamp 1701704242
transform 1 0 11500 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[8\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 12512 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[8\].stg01
timestamp 1701704242
transform -1 0 11224 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[8\].stg02
timestamp 1701704242
transform -1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[9\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 28152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[9\].stg01
timestamp 1701704242
transform -1 0 14536 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[9\].stg02
timestamp 1701704242
transform -1 0 27232 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[10\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 26772 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[10\].stg01
timestamp 1701704242
transform -1 0 27324 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[10\].stg02
timestamp 1701704242
transform -1 0 27600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[11\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 28152 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[11\].stg01
timestamp 1701704242
transform 1 0 26680 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[11\].stg02
timestamp 1701704242
transform -1 0 27692 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[12\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[12\].stg01
timestamp 1701704242
transform 1 0 26956 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[12\].stg02
timestamp 1701704242
transform 1 0 26588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[13\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[13\].stg01
timestamp 1701704242
transform 1 0 25668 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[13\].stg02
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[14\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 18400 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[14\].stg01
timestamp 1701704242
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[14\].stg02
timestamp 1701704242
transform 1 0 12788 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[15\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 7820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[15\].stg01
timestamp 1701704242
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[15\].stg02
timestamp 1701704242
transform 1 0 7452 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[16\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[16\].stg01
timestamp 1701704242
transform 1 0 6900 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  tdc1.g_ring1\[16\].stg02 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring1\[16\].stg02_60
timestamp 1701704242
transform 1 0 6256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[16\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 7360 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[16\].stg01_61
timestamp 1701704242
transform -1 0 6256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[16\].stg01
timestamp 1701704242
transform -1 0 5428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  tdc1.g_ring3\[16\].stg02
timestamp 1701704242
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[17\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 24104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[17\].stg01_62
timestamp 1701704242
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[17\].stg01
timestamp 1701704242
transform -1 0 7544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[17\].stg02
timestamp 1701704242
transform -1 0 23184 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[18\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 23184 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[18\].stg01_63
timestamp 1701704242
transform 1 0 23552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[18\].stg01
timestamp 1701704242
transform 1 0 24196 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[18\].stg02
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[19\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 24104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[19\].stg01
timestamp 1701704242
transform -1 0 24288 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[19\].stg01_64
timestamp 1701704242
transform 1 0 23460 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[19\].stg02
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[20\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 23184 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[20\].stg01_65
timestamp 1701704242
transform 1 0 23184 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[20\].stg01
timestamp 1701704242
transform 1 0 23460 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[20\].stg02
timestamp 1701704242
transform 1 0 23184 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[21\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[21\].stg01
timestamp 1701704242
transform 1 0 22632 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[21\].stg01_66
timestamp 1701704242
transform 1 0 22356 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[21\].stg02
timestamp 1701704242
transform 1 0 17388 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[22\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[22\].stg01_67
timestamp 1701704242
transform -1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[22\].stg01
timestamp 1701704242
transform 1 0 17112 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[22\].stg02
timestamp 1701704242
transform -1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[23\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 9384 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[23\].stg01
timestamp 1701704242
transform 1 0 11776 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[23\].stg01_68
timestamp 1701704242
transform 1 0 11500 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[23\].stg02
timestamp 1701704242
transform 1 0 11132 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[24\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[24\].stg01_69
timestamp 1701704242
transform -1 0 11500 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[24\].stg01
timestamp 1701704242
transform -1 0 10948 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[24\].stg02
timestamp 1701704242
transform -1 0 12236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[25\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 28520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[25\].stg01_70
timestamp 1701704242
transform 1 0 12052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[25\].stg01
timestamp 1701704242
transform 1 0 12236 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[25\].stg02
timestamp 1701704242
transform -1 0 26864 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[26\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 27692 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[26\].stg01_71
timestamp 1701704242
transform -1 0 28244 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[26\].stg01
timestamp 1701704242
transform -1 0 27968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[26\].stg02
timestamp 1701704242
transform 1 0 27600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[27\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 28428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[27\].stg01_72
timestamp 1701704242
transform -1 0 28244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[27\].stg01
timestamp 1701704242
transform -1 0 26680 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[27\].stg02
timestamp 1701704242
transform -1 0 28060 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[28\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 27324 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[28\].stg01_73
timestamp 1701704242
transform -1 0 26588 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[28\].stg01
timestamp 1701704242
transform 1 0 26036 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[28\].stg02
timestamp 1701704242
transform -1 0 26312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[29\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 15272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[29\].stg01_74
timestamp 1701704242
transform -1 0 27140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[29\].stg01
timestamp 1701704242
transform 1 0 25944 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[29\].stg02
timestamp 1701704242
transform 1 0 19044 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[30\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 8740 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[30\].stg01_75
timestamp 1701704242
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[30\].stg01
timestamp 1701704242
transform -1 0 14444 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[30\].stg02
timestamp 1701704242
transform -1 0 14812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[31\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[31\].stg01_76
timestamp 1701704242
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[31\].stg01
timestamp 1701704242
transform 1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[31\].stg02
timestamp 1701704242
transform 1 0 7820 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tdc1.stg01_77
timestamp 1701704242
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.stg01
timestamp 1701704242
transform 1 0 6624 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  tdc1.stg02
timestamp 1701704242
transform 1 0 6716 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_78
timestamp 1701704242
transform -1 0 20332 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_79
timestamp 1701704242
transform -1 0 19688 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_80
timestamp 1701704242
transform -1 0 19044 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_81
timestamp 1701704242
transform -1 0 16468 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_82
timestamp 1701704242
transform -1 0 22264 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_83
timestamp 1701704242
transform -1 0 20976 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_84
timestamp 1701704242
transform -1 0 19044 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_85
timestamp 1701704242
transform -1 0 12604 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_86
timestamp 1701704242
transform -1 0 10672 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_87
timestamp 1701704242
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_88
timestamp 1701704242
transform -1 0 11316 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_89
timestamp 1701704242
transform -1 0 13248 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_90
timestamp 1701704242
transform -1 0 6808 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_91
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_92
timestamp 1701704242
transform -1 0 14536 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_93
timestamp 1701704242
transform -1 0 18400 0 -1 19040
box -38 -48 314 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 662 0 718 400 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 1306 0 1362 400 0 FreeSans 224 90 0 0 ena
port 3 nsew signal input
flabel metal2 s 1950 0 2006 400 0 FreeSans 224 90 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 31600 7488 32000 7608 0 FreeSans 480 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 14288 400 14408 0 FreeSans 480 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 10208 400 10328 0 FreeSans 480 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal2 s 2594 0 2650 400 0 FreeSans 224 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal2 s 3238 0 3294 400 0 FreeSans 224 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal2 s 3882 0 3938 400 0 FreeSans 224 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal2 s 4526 0 4582 400 0 FreeSans 224 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal2 s 5170 0 5226 400 0 FreeSans 224 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal2 s 5814 0 5870 400 0 FreeSans 224 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal2 s 7102 0 7158 400 0 FreeSans 224 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal2 s 18 0 74 400 0 FreeSans 224 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal2 s 8390 0 8446 400 0 FreeSans 224 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal2 s 16118 19600 16174 20000 0 FreeSans 224 90 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal2 s 21914 19600 21970 20000 0 FreeSans 224 90 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal2 s 20626 19600 20682 20000 0 FreeSans 224 90 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal2 s 12254 19600 12310 20000 0 FreeSans 224 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal2 s 10322 19600 10378 20000 0 FreeSans 224 90 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal2 s 21270 19600 21326 20000 0 FreeSans 224 90 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal2 s 10966 19600 11022 20000 0 FreeSans 224 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal2 s 12898 19600 12954 20000 0 FreeSans 224 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal2 s 6458 0 6514 400 0 FreeSans 224 90 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal3 s 31600 18368 32000 18488 0 FreeSans 480 0 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal3 s 31600 12248 32000 12368 0 FreeSans 480 0 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal3 s 31600 6808 32000 6928 0 FreeSans 480 0 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal2 s 15474 19600 15530 20000 0 FreeSans 224 90 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal2 s 11610 19600 11666 20000 0 FreeSans 224 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal1 18630 15674 18630 15674 0 _000_
rlabel metal1 17710 14552 17710 14552 0 _001_
rlabel metal2 15318 14076 15318 14076 0 _002_
rlabel metal1 4048 14382 4048 14382 0 _003_
rlabel metal1 6578 14552 6578 14552 0 _004_
rlabel metal1 3864 12818 3864 12818 0 _005_
rlabel metal1 3772 11254 3772 11254 0 _006_
rlabel metal1 20608 15402 20608 15402 0 _007_
rlabel metal1 21620 14858 21620 14858 0 _008_
rlabel metal1 22126 15640 22126 15640 0 _009_
rlabel metal1 11500 16218 11500 16218 0 _010_
rlabel metal1 11868 14858 11868 14858 0 _011_
rlabel metal1 9844 16082 9844 16082 0 _012_
rlabel metal1 7728 15470 7728 15470 0 _013_
rlabel metal1 13662 16082 13662 16082 0 _014_
rlabel metal1 16366 16218 16366 16218 0 _015_
rlabel metal1 19136 3638 19136 3638 0 _016_
rlabel metal1 16238 4522 16238 4522 0 _017_
rlabel metal2 15042 5372 15042 5372 0 _018_
rlabel metal1 7222 4760 7222 4760 0 _019_
rlabel metal1 4416 4726 4416 4726 0 _020_
rlabel metal2 3634 6018 3634 6018 0 _021_
rlabel metal1 3312 7378 3312 7378 0 _022_
rlabel metal1 21574 3162 21574 3162 0 _023_
rlabel metal1 20884 4250 20884 4250 0 _024_
rlabel metal1 22402 4114 22402 4114 0 _025_
rlabel metal2 16974 3128 16974 3128 0 _026_
rlabel metal1 11454 3026 11454 3026 0 _027_
rlabel metal1 8924 3502 8924 3502 0 _028_
rlabel metal1 8832 3910 8832 3910 0 _029_
rlabel metal1 13386 3434 13386 3434 0 _030_
rlabel metal1 15502 3944 15502 3944 0 _031_
rlabel metal1 19320 15674 19320 15674 0 _032_
rlabel metal2 21574 16184 21574 16184 0 _033_
rlabel metal2 22678 14722 22678 14722 0 _034_
rlabel metal2 22862 15742 22862 15742 0 _035_
rlabel metal1 12604 16218 12604 16218 0 _036_
rlabel metal1 13393 14858 13393 14858 0 _037_
rlabel metal2 9154 16184 9154 16184 0 _038_
rlabel metal2 7958 15368 7958 15368 0 _039_
rlabel metal1 14720 15674 14720 15674 0 _040_
rlabel metal1 18039 15946 18039 15946 0 _041_
rlabel metal2 18446 14654 18446 14654 0 _042_
rlabel metal1 15962 13226 15962 13226 0 _043_
rlabel metal1 4876 14586 4876 14586 0 _044_
rlabel metal1 7544 14042 7544 14042 0 _045_
rlabel metal1 4094 12410 4094 12410 0 _046_
rlabel metal1 3411 11254 3411 11254 0 _047_
rlabel metal1 20148 3162 20148 3162 0 _048_
rlabel metal1 23329 3638 23329 3638 0 _049_
rlabel metal1 19596 4250 19596 4250 0 _050_
rlabel metal2 22954 4216 22954 4216 0 _051_
rlabel metal1 18499 2890 18499 2890 0 _052_
rlabel metal1 12703 2890 12703 2890 0 _053_
rlabel metal2 9154 3400 9154 3400 0 _054_
rlabel metal1 7866 4087 7866 4087 0 _055_
rlabel metal1 15141 3638 15141 3638 0 _056_
rlabel metal1 18407 3978 18407 3978 0 _057_
rlabel metal1 17940 4998 17940 4998 0 _058_
rlabel metal1 16199 5134 16199 5134 0 _059_
rlabel metal2 7958 4862 7958 4862 0 _060_
rlabel metal1 4416 4794 4416 4794 0 _061_
rlabel metal1 5067 6154 5067 6154 0 _062_
rlabel metal2 4278 7106 4278 7106 0 _063_
rlabel metal1 19826 8058 19826 8058 0 _064_
rlabel metal1 19826 7922 19826 7922 0 _065_
rlabel metal2 21758 7786 21758 7786 0 _066_
rlabel metal2 13018 7650 13018 7650 0 _067_
rlabel metal1 11132 10574 11132 10574 0 _068_
rlabel metal1 11362 9078 11362 9078 0 _069_
rlabel metal2 14766 9554 14766 9554 0 _070_
rlabel metal1 15042 9146 15042 9146 0 _071_
rlabel metal2 12742 10880 12742 10880 0 _072_
rlabel metal1 26082 8942 26082 8942 0 _073_
rlabel metal1 15640 10506 15640 10506 0 _074_
rlabel metal1 13386 6154 13386 6154 0 _075_
rlabel metal1 13892 8874 13892 8874 0 _076_
rlabel metal2 20746 6307 20746 6307 0 _077_
rlabel metal2 25254 7684 25254 7684 0 _078_
rlabel metal2 25622 9588 25622 9588 0 _079_
rlabel viali 21761 9418 21761 9418 0 _080_
rlabel metal1 21758 9486 21758 9486 0 _081_
rlabel metal1 20056 8602 20056 8602 0 _082_
rlabel metal1 21252 12682 21252 12682 0 _083_
rlabel metal1 22310 9486 22310 9486 0 _084_
rlabel metal1 25162 9690 25162 9690 0 _085_
rlabel metal1 10442 9350 10442 9350 0 _086_
rlabel metal2 20194 12891 20194 12891 0 _087_
rlabel metal1 21206 12784 21206 12784 0 _088_
rlabel metal1 20884 12750 20884 12750 0 _089_
rlabel metal1 23966 12648 23966 12648 0 _090_
rlabel metal2 26910 12954 26910 12954 0 _091_
rlabel metal2 26266 12138 26266 12138 0 _092_
rlabel metal1 26404 11662 26404 11662 0 _093_
rlabel metal1 20976 7310 20976 7310 0 _094_
rlabel metal1 24058 7480 24058 7480 0 _095_
rlabel metal1 27600 9622 27600 9622 0 _096_
rlabel metal2 24334 9503 24334 9503 0 _097_
rlabel metal1 26542 9690 26542 9690 0 _098_
rlabel metal1 21390 7752 21390 7752 0 _099_
rlabel metal1 25760 7514 25760 7514 0 _100_
rlabel metal1 27784 8058 27784 8058 0 _101_
rlabel metal1 25392 8602 25392 8602 0 _102_
rlabel metal2 24518 13396 24518 13396 0 _103_
rlabel metal1 25484 13702 25484 13702 0 _104_
rlabel metal1 25944 10574 25944 10574 0 _105_
rlabel metal1 27784 6358 27784 6358 0 _106_
rlabel via2 21758 6749 21758 6749 0 _107_
rlabel metal1 21942 6766 21942 6766 0 _108_
rlabel metal1 21160 10098 21160 10098 0 _109_
rlabel metal2 20378 10455 20378 10455 0 _110_
rlabel metal1 21988 9486 21988 9486 0 _111_
rlabel metal1 21114 9690 21114 9690 0 _112_
rlabel metal2 22310 8330 22310 8330 0 _113_
rlabel metal1 15456 10642 15456 10642 0 _114_
rlabel metal1 15686 10778 15686 10778 0 _115_
rlabel metal1 15272 10574 15272 10574 0 _116_
rlabel metal2 15502 9962 15502 9962 0 _117_
rlabel metal1 15364 7922 15364 7922 0 _118_
rlabel metal1 15686 7718 15686 7718 0 _119_
rlabel metal1 14628 7514 14628 7514 0 _120_
rlabel metal2 15410 8772 15410 8772 0 _121_
rlabel metal1 16238 9486 16238 9486 0 _122_
rlabel metal1 11086 12750 11086 12750 0 _123_
rlabel metal1 11638 12308 11638 12308 0 _124_
rlabel metal1 11776 11866 11776 11866 0 _125_
rlabel metal1 12052 6426 12052 6426 0 _126_
rlabel metal1 11132 5882 11132 5882 0 _127_
rlabel metal1 19182 8058 19182 8058 0 _128_
rlabel metal2 18722 7497 18722 7497 0 _129_
rlabel metal1 12006 6630 12006 6630 0 _130_
rlabel metal2 10534 7684 10534 7684 0 _131_
rlabel metal2 10442 7616 10442 7616 0 _132_
rlabel metal1 10206 7928 10206 7928 0 _133_
rlabel metal1 10856 8058 10856 8058 0 _134_
rlabel metal1 11086 10132 11086 10132 0 _135_
rlabel metal1 10856 9894 10856 9894 0 _136_
rlabel metal1 10902 10098 10902 10098 0 _137_
rlabel metal1 10948 9554 10948 9554 0 _138_
rlabel metal1 10718 9520 10718 9520 0 _139_
rlabel metal1 21068 14926 21068 14926 0 _140_
rlabel metal1 21068 15130 21068 15130 0 _141_
rlabel metal2 20654 15334 20654 15334 0 _142_
rlabel metal1 19274 15606 19274 15606 0 _143_
rlabel metal1 21436 15538 21436 15538 0 _144_
rlabel metal1 10810 15130 10810 15130 0 _145_
rlabel metal1 10580 15674 10580 15674 0 _146_
rlabel metal1 11914 15504 11914 15504 0 _147_
rlabel metal1 9568 15334 9568 15334 0 _148_
rlabel metal1 10396 16218 10396 16218 0 _149_
rlabel metal1 9706 14858 9706 14858 0 _150_
rlabel metal1 10718 14858 10718 14858 0 _151_
rlabel metal1 12926 16014 12926 16014 0 _152_
rlabel metal1 15732 15674 15732 15674 0 _153_
rlabel metal1 16698 15028 16698 15028 0 _154_
rlabel metal1 15640 14382 15640 14382 0 _155_
rlabel metal1 15042 15028 15042 15028 0 _156_
rlabel metal1 9062 15096 9062 15096 0 _157_
rlabel metal1 6992 13838 6992 13838 0 _158_
rlabel metal1 6256 14586 6256 14586 0 _159_
rlabel metal2 6486 14416 6486 14416 0 _160_
rlabel metal1 4554 13362 4554 13362 0 _161_
rlabel metal2 4186 13515 4186 13515 0 _162_
rlabel metal1 20746 4080 20746 4080 0 _163_
rlabel metal1 21564 4522 21564 4522 0 _164_
rlabel metal1 21942 4658 21942 4658 0 _165_
rlabel metal1 11316 4250 11316 4250 0 _166_
rlabel metal1 22586 4624 22586 4624 0 _167_
rlabel metal1 10810 4216 10810 4216 0 _168_
rlabel metal1 10672 3638 10672 3638 0 _169_
rlabel metal1 11638 3536 11638 3536 0 _170_
rlabel metal1 9798 3978 9798 3978 0 _171_
rlabel metal1 10442 3536 10442 3536 0 _172_
rlabel metal1 10350 4658 10350 4658 0 _173_
rlabel metal1 11086 4250 11086 4250 0 _174_
rlabel metal1 13992 4794 13992 4794 0 _175_
rlabel metal1 15548 4182 15548 4182 0 _176_
rlabel metal1 14306 4556 14306 4556 0 _177_
rlabel metal1 14490 4794 14490 4794 0 _178_
rlabel metal2 13294 4896 13294 4896 0 _179_
rlabel metal1 13386 4250 13386 4250 0 _180_
rlabel metal1 6578 5236 6578 5236 0 _181_
rlabel metal1 5750 4658 5750 4658 0 _182_
rlabel metal1 5382 4726 5382 4726 0 _183_
rlabel metal1 3174 5746 3174 5746 0 _184_
rlabel metal1 3726 5712 3726 5712 0 _185_
rlabel metal1 13800 8602 13800 8602 0 _186_
rlabel metal1 13478 8806 13478 8806 0 _187_
rlabel metal1 13524 8058 13524 8058 0 _188_
rlabel metal1 14260 9146 14260 9146 0 _189_
rlabel metal2 14306 11084 14306 11084 0 _190_
rlabel metal1 12742 10778 12742 10778 0 _191_
rlabel metal1 14168 10574 14168 10574 0 _192_
rlabel metal2 14674 9962 14674 9962 0 _193_
rlabel metal1 9430 9452 9430 9452 0 _194_
rlabel metal1 21482 16592 21482 16592 0 _195_
rlabel metal1 9062 2890 9062 2890 0 _196_
rlabel metal2 16882 12580 16882 12580 0 net1
rlabel metal1 21574 14994 21574 14994 0 net10
rlabel metal2 5474 12461 5474 12461 0 net11
rlabel metal1 22402 12274 22402 12274 0 net12
rlabel metal1 7130 7344 7130 7344 0 net13
rlabel metal2 14674 6154 14674 6154 0 net14
rlabel metal1 8694 4046 8694 4046 0 net15
rlabel metal2 9430 4828 9430 4828 0 net16
rlabel metal1 23966 8398 23966 8398 0 net17
rlabel metal1 26450 6834 26450 6834 0 net18
rlabel metal1 19136 6222 19136 6222 0 net19
rlabel metal1 506 14144 506 14144 0 net2
rlabel metal1 6992 12274 6992 12274 0 net20
rlabel metal1 3634 12342 3634 12342 0 net21
rlabel metal1 18722 14858 18722 14858 0 net22
rlabel metal1 16330 13396 16330 13396 0 net23
rlabel via2 4094 13243 4094 13243 0 net24
rlabel metal1 14858 10166 14858 10166 0 net25
rlabel metal2 6854 5780 6854 5780 0 net26
rlabel metal1 2392 13838 2392 13838 0 net27
rlabel metal1 2990 14450 2990 14450 0 net28
rlabel metal1 13432 13906 13432 13906 0 net29
rlabel metal1 1909 10778 1909 10778 0 net3
rlabel metal1 14214 5610 14214 5610 0 net30
rlabel metal1 20102 6324 20102 6324 0 net31
rlabel metal2 18722 13940 18722 13940 0 net32
rlabel metal1 21528 13294 21528 13294 0 net33
rlabel metal2 24058 6290 24058 6290 0 net34
rlabel metal1 23690 10540 23690 10540 0 net35
rlabel metal1 26634 5236 26634 5236 0 net36
rlabel metal1 2622 14484 2622 14484 0 net37
rlabel metal1 9016 11186 9016 11186 0 net38
rlabel metal1 14444 8398 14444 8398 0 net39
rlabel metal1 16744 8398 16744 8398 0 net4
rlabel metal1 23138 7956 23138 7956 0 net40
rlabel metal1 18722 7344 18722 7344 0 net41
rlabel metal1 5014 12308 5014 12308 0 net42
rlabel metal2 6670 12789 6670 12789 0 net43
rlabel metal1 5060 13158 5060 13158 0 net44
rlabel metal1 16514 12886 16514 12886 0 net45
rlabel metal1 23552 12886 23552 12886 0 net46
rlabel metal1 22448 11662 22448 11662 0 net47
rlabel metal1 17158 11050 17158 11050 0 net48
rlabel metal1 12558 11254 12558 11254 0 net49
rlabel metal1 16698 7990 16698 7990 0 net5
rlabel metal1 9522 11696 9522 11696 0 net50
rlabel metal1 7958 11696 7958 11696 0 net51
rlabel metal1 12880 11662 12880 11662 0 net52
rlabel metal1 18538 11662 18538 11662 0 net53
rlabel metal1 21804 11866 21804 11866 0 net54
rlabel metal1 20286 11220 20286 11220 0 net55
rlabel metal1 17480 12206 17480 12206 0 net56
rlabel metal1 12834 12784 12834 12784 0 net57
rlabel metal2 7682 12206 7682 12206 0 net58
rlabel metal1 5566 12784 5566 12784 0 net59
rlabel metal1 16560 9010 16560 9010 0 net6
rlabel metal1 6578 7922 6578 7922 0 net60
rlabel metal1 5704 7922 5704 7922 0 net61
rlabel metal1 7498 8432 7498 8432 0 net62
rlabel metal1 24242 8432 24242 8432 0 net63
rlabel metal1 23966 7854 23966 7854 0 net64
rlabel metal1 23460 6222 23460 6222 0 net65
rlabel metal1 22632 6222 22632 6222 0 net66
rlabel metal1 17158 6800 17158 6800 0 net67
rlabel metal1 11776 7310 11776 7310 0 net68
rlabel metal1 10902 8432 10902 8432 0 net69
rlabel metal1 10994 3094 10994 3094 0 net7
rlabel metal1 12328 8398 12328 8398 0 net70
rlabel metal2 27922 8602 27922 8602 0 net71
rlabel metal1 26634 8432 26634 8432 0 net72
rlabel metal1 26082 7344 26082 7344 0 net73
rlabel metal2 25990 6324 25990 6324 0 net74
rlabel metal1 14398 6256 14398 6256 0 net75
rlabel metal1 8418 6868 8418 6868 0 net76
rlabel metal1 6440 7310 6440 7310 0 net77
rlabel metal1 20056 18802 20056 18802 0 net78
rlabel metal1 19412 18802 19412 18802 0 net79
rlabel metal1 15456 5542 15456 5542 0 net8
rlabel metal1 18768 18802 18768 18802 0 net80
rlabel metal2 16238 19023 16238 19023 0 net81
rlabel metal1 21988 18802 21988 18802 0 net82
rlabel metal1 20700 18802 20700 18802 0 net83
rlabel metal2 18722 415 18722 415 0 net84
rlabel metal1 12328 18802 12328 18802 0 net85
rlabel metal1 10396 18802 10396 18802 0 net86
rlabel metal1 21344 18802 21344 18802 0 net87
rlabel metal1 11040 18802 11040 18802 0 net88
rlabel metal1 12972 18802 12972 18802 0 net89
rlabel metal1 18492 16082 18492 16082 0 net9
rlabel metal2 6486 415 6486 415 0 net90
rlabel metal3 31380 18428 31380 18428 0 net91
rlabel metal2 14214 415 14214 415 0 net92
rlabel metal1 18124 18802 18124 18802 0 net93
rlabel metal1 14306 10506 14306 10506 0 tdc0.r_dly_store_ctr\[0\]
rlabel metal2 25530 13260 25530 13260 0 tdc0.r_dly_store_ctr\[10\]
rlabel viali 24794 13838 24794 13838 0 tdc0.r_dly_store_ctr\[11\]
rlabel metal2 11638 13124 11638 13124 0 tdc0.r_dly_store_ctr\[12\]
rlabel metal2 10626 13328 10626 13328 0 tdc0.r_dly_store_ctr\[13\]
rlabel metal1 10166 13396 10166 13396 0 tdc0.r_dly_store_ctr\[14\]
rlabel metal2 10166 10438 10166 10438 0 tdc0.r_dly_store_ctr\[15\]
rlabel metal2 20562 13532 20562 13532 0 tdc0.r_dly_store_ctr\[1\]
rlabel metal1 26496 13430 26496 13430 0 tdc0.r_dly_store_ctr\[2\]
rlabel metal2 25070 14314 25070 14314 0 tdc0.r_dly_store_ctr\[3\]
rlabel metal2 12742 13838 12742 13838 0 tdc0.r_dly_store_ctr\[4\]
rlabel metal1 14950 14314 14950 14314 0 tdc0.r_dly_store_ctr\[5\]
rlabel via1 11546 12750 11546 12750 0 tdc0.r_dly_store_ctr\[6\]
rlabel metal1 9706 14246 9706 14246 0 tdc0.r_dly_store_ctr\[7\]
rlabel metal2 13892 12716 13892 12716 0 tdc0.r_dly_store_ctr\[8\]
rlabel via1 20286 13362 20286 13362 0 tdc0.r_dly_store_ctr\[9\]
rlabel metal1 4876 9418 4876 9418 0 tdc0.r_dly_store_ring\[0\]
rlabel metal1 26358 13362 26358 13362 0 tdc0.r_dly_store_ring\[10\]
rlabel metal1 23966 12784 23966 12784 0 tdc0.r_dly_store_ring\[11\]
rlabel metal1 21896 10574 21896 10574 0 tdc0.r_dly_store_ring\[12\]
rlabel metal1 15548 11662 15548 11662 0 tdc0.r_dly_store_ring\[13\]
rlabel metal1 11454 11696 11454 11696 0 tdc0.r_dly_store_ring\[14\]
rlabel viali 9522 10098 9522 10098 0 tdc0.r_dly_store_ring\[15\]
rlabel metal1 10718 10540 10718 10540 0 tdc0.r_dly_store_ring\[16\]
rlabel metal1 19090 13328 19090 13328 0 tdc0.r_dly_store_ring\[17\]
rlabel metal1 27462 12070 27462 12070 0 tdc0.r_dly_store_ring\[18\]
rlabel metal1 24242 12784 24242 12784 0 tdc0.r_dly_store_ring\[19\]
rlabel metal1 21344 12750 21344 12750 0 tdc0.r_dly_store_ring\[1\]
rlabel metal1 21666 10472 21666 10472 0 tdc0.r_dly_store_ring\[20\]
rlabel metal1 15318 11254 15318 11254 0 tdc0.r_dly_store_ring\[21\]
rlabel metal1 11822 12784 11822 12784 0 tdc0.r_dly_store_ring\[22\]
rlabel metal1 10442 10064 10442 10064 0 tdc0.r_dly_store_ring\[23\]
rlabel metal1 10902 10574 10902 10574 0 tdc0.r_dly_store_ring\[24\]
rlabel metal1 19780 10234 19780 10234 0 tdc0.r_dly_store_ring\[25\]
rlabel metal1 27600 12410 27600 12410 0 tdc0.r_dly_store_ring\[26\]
rlabel metal1 25898 11288 25898 11288 0 tdc0.r_dly_store_ring\[27\]
rlabel metal1 20298 9554 20298 9554 0 tdc0.r_dly_store_ring\[28\]
rlabel metal1 15134 13430 15134 13430 0 tdc0.r_dly_store_ring\[29\]
rlabel metal1 25714 12376 25714 12376 0 tdc0.r_dly_store_ring\[2\]
rlabel metal1 10350 13362 10350 13362 0 tdc0.r_dly_store_ring\[30\]
rlabel metal1 10074 10676 10074 10676 0 tdc0.r_dly_store_ring\[31\]
rlabel viali 25622 11186 25622 11186 0 tdc0.r_dly_store_ring\[3\]
rlabel via1 21850 9435 21850 9435 0 tdc0.r_dly_store_ring\[4\]
rlabel metal1 17848 10234 17848 10234 0 tdc0.r_dly_store_ring\[5\]
rlabel viali 11178 11662 11178 11662 0 tdc0.r_dly_store_ring\[6\]
rlabel metal1 5888 9486 5888 9486 0 tdc0.r_dly_store_ring\[7\]
rlabel metal1 13340 10574 13340 10574 0 tdc0.r_dly_store_ring\[8\]
rlabel metal1 18676 12954 18676 12954 0 tdc0.r_dly_store_ring\[9\]
rlabel metal1 18262 15538 18262 15538 0 tdc0.r_ring_ctr\[0\]
rlabel metal1 23497 14416 23497 14416 0 tdc0.r_ring_ctr\[10\]
rlabel metal1 16790 13872 16790 13872 0 tdc0.r_ring_ctr\[11\]
rlabel metal2 6854 13226 6854 13226 0 tdc0.r_ring_ctr\[12\]
rlabel metal1 7585 13430 7585 13430 0 tdc0.r_ring_ctr\[13\]
rlabel metal1 5136 13770 5136 13770 0 tdc0.r_ring_ctr\[14\]
rlabel metal1 3496 11662 3496 11662 0 tdc0.r_ring_ctr\[15\]
rlabel metal1 20930 15096 20930 15096 0 tdc0.r_ring_ctr\[1\]
rlabel metal1 23644 14790 23644 14790 0 tdc0.r_ring_ctr\[2\]
rlabel metal1 23874 15334 23874 15334 0 tdc0.r_ring_ctr\[3\]
rlabel metal2 11454 16048 11454 16048 0 tdc0.r_ring_ctr\[4\]
rlabel metal1 13462 14518 13462 14518 0 tdc0.r_ring_ctr\[5\]
rlabel metal1 9108 14926 9108 14926 0 tdc0.r_ring_ctr\[6\]
rlabel metal1 9108 15538 9108 15538 0 tdc0.r_ring_ctr\[7\]
rlabel metal1 14214 16218 14214 16218 0 tdc0.r_ring_ctr\[8\]
rlabel metal1 18216 15878 18216 15878 0 tdc0.r_ring_ctr\[9\]
rlabel metal1 2576 13838 2576 13838 0 tdc0.w_dly_stop\[1\]
rlabel metal1 2806 13430 2806 13430 0 tdc0.w_dly_stop\[2\]
rlabel metal1 2944 13498 2944 13498 0 tdc0.w_dly_stop\[3\]
rlabel metal1 3128 13362 3128 13362 0 tdc0.w_dly_stop\[4\]
rlabel metal1 3634 13430 3634 13430 0 tdc0.w_dly_stop\[5\]
rlabel metal2 15134 15538 15134 15538 0 tdc0.w_ring_buf\[0\]
rlabel metal1 25070 12954 25070 12954 0 tdc0.w_ring_buf\[10\]
rlabel metal1 21988 12954 21988 12954 0 tdc0.w_ring_buf\[11\]
rlabel metal1 20148 11322 20148 11322 0 tdc0.w_ring_buf\[12\]
rlabel metal1 14531 12342 14531 12342 0 tdc0.w_ring_buf\[13\]
rlabel metal1 9660 12614 9660 12614 0 tdc0.w_ring_buf\[14\]
rlabel metal1 6619 10166 6619 10166 0 tdc0.w_ring_buf\[15\]
rlabel via1 4998 11594 4998 11594 0 tdc0.w_ring_buf\[16\]
rlabel metal1 16100 12954 16100 12954 0 tdc0.w_ring_buf\[17\]
rlabel metal1 26480 12342 26480 12342 0 tdc0.w_ring_buf\[18\]
rlabel metal2 23506 13158 23506 13158 0 tdc0.w_ring_buf\[19\]
rlabel metal1 19887 12648 19887 12648 0 tdc0.w_ring_buf\[1\]
rlabel metal1 23234 10574 23234 10574 0 tdc0.w_ring_buf\[20\]
rlabel metal1 13830 11254 13830 11254 0 tdc0.w_ring_buf\[21\]
rlabel via1 11265 13362 11265 13362 0 tdc0.w_ring_buf\[22\]
rlabel via1 7953 10098 7953 10098 0 tdc0.w_ring_buf\[23\]
rlabel metal1 9506 11254 9506 11254 0 tdc0.w_ring_buf\[24\]
rlabel metal1 18896 10574 18896 10574 0 tdc0.w_ring_buf\[25\]
rlabel metal2 27738 12070 27738 12070 0 tdc0.w_ring_buf\[26\]
rlabel metal1 26868 11254 26868 11254 0 tdc0.w_ring_buf\[27\]
rlabel metal1 18522 11254 18522 11254 0 tdc0.w_ring_buf\[28\]
rlabel metal1 14260 12614 14260 12614 0 tdc0.w_ring_buf\[29\]
rlabel metal1 24104 11866 24104 11866 0 tdc0.w_ring_buf\[2\]
rlabel metal2 8786 13158 8786 13158 0 tdc0.w_ring_buf\[30\]
rlabel via1 5929 10574 5929 10574 0 tdc0.w_ring_buf\[31\]
rlabel metal1 24134 11254 24134 11254 0 tdc0.w_ring_buf\[3\]
rlabel metal1 21236 10166 21236 10166 0 tdc0.w_ring_buf\[4\]
rlabel metal1 16458 10098 16458 10098 0 tdc0.w_ring_buf\[5\]
rlabel metal2 8694 12070 8694 12070 0 tdc0.w_ring_buf\[6\]
rlabel metal1 4779 10166 4779 10166 0 tdc0.w_ring_buf\[7\]
rlabel metal1 11806 10506 11806 10506 0 tdc0.w_ring_buf\[8\]
rlabel metal1 17659 12682 17659 12682 0 tdc0.w_ring_buf\[9\]
rlabel metal2 5612 12342 5612 12342 0 tdc0.w_ring_int_norsz\[0\]
rlabel metal1 18584 12342 18584 12342 0 tdc0.w_ring_int_norsz\[10\]
rlabel metal1 21160 12206 21160 12206 0 tdc0.w_ring_int_norsz\[11\]
rlabel metal1 20194 12206 20194 12206 0 tdc0.w_ring_int_norsz\[12\]
rlabel via2 19182 11883 19182 11883 0 tdc0.w_ring_int_norsz\[13\]
rlabel metal1 13110 12342 13110 12342 0 tdc0.w_ring_int_norsz\[14\]
rlabel metal1 7498 12342 7498 12342 0 tdc0.w_ring_int_norsz\[15\]
rlabel metal2 6118 12036 6118 12036 0 tdc0.w_ring_int_norsz\[16\]
rlabel metal2 15778 12716 15778 12716 0 tdc0.w_ring_int_norsz\[17\]
rlabel metal1 21850 12274 21850 12274 0 tdc0.w_ring_int_norsz\[18\]
rlabel metal1 23460 11730 23460 11730 0 tdc0.w_ring_int_norsz\[19\]
rlabel metal1 16606 12206 16606 12206 0 tdc0.w_ring_int_norsz\[1\]
rlabel metal1 22540 11254 22540 11254 0 tdc0.w_ring_int_norsz\[20\]
rlabel metal1 16974 11118 16974 11118 0 tdc0.w_ring_int_norsz\[21\]
rlabel metal1 12098 11118 12098 11118 0 tdc0.w_ring_int_norsz\[22\]
rlabel metal2 7958 11322 7958 11322 0 tdc0.w_ring_int_norsz\[23\]
rlabel metal1 8464 11118 8464 11118 0 tdc0.w_ring_int_norsz\[24\]
rlabel metal1 16836 11730 16836 11730 0 tdc0.w_ring_int_norsz\[25\]
rlabel metal1 18446 11866 18446 11866 0 tdc0.w_ring_int_norsz\[26\]
rlabel metal1 22034 12172 22034 12172 0 tdc0.w_ring_int_norsz\[27\]
rlabel metal1 20332 11322 20332 11322 0 tdc0.w_ring_int_norsz\[28\]
rlabel metal1 14582 12274 14582 12274 0 tdc0.w_ring_int_norsz\[29\]
rlabel metal1 22448 12342 22448 12342 0 tdc0.w_ring_int_norsz\[2\]
rlabel metal1 12834 12682 12834 12682 0 tdc0.w_ring_int_norsz\[30\]
rlabel metal1 7636 11866 7636 11866 0 tdc0.w_ring_int_norsz\[31\]
rlabel metal1 23138 11730 23138 11730 0 tdc0.w_ring_int_norsz\[3\]
rlabel metal1 22724 11118 22724 11118 0 tdc0.w_ring_int_norsz\[4\]
rlabel metal2 16514 11118 16514 11118 0 tdc0.w_ring_int_norsz\[5\]
rlabel metal1 11868 11322 11868 11322 0 tdc0.w_ring_int_norsz\[6\]
rlabel metal2 7590 11390 7590 11390 0 tdc0.w_ring_int_norsz\[7\]
rlabel metal1 8740 11254 8740 11254 0 tdc0.w_ring_int_norsz\[8\]
rlabel metal1 13386 11050 13386 11050 0 tdc0.w_ring_int_norsz\[9\]
rlabel metal2 5290 12580 5290 12580 0 tdc0.w_ring_norsz\[0\]
rlabel metal1 18722 12104 18722 12104 0 tdc0.w_ring_norsz\[10\]
rlabel metal1 21668 12138 21668 12138 0 tdc0.w_ring_norsz\[11\]
rlabel metal1 19596 11798 19596 11798 0 tdc0.w_ring_norsz\[12\]
rlabel metal1 13294 12784 13294 12784 0 tdc0.w_ring_norsz\[13\]
rlabel metal1 7866 12648 7866 12648 0 tdc0.w_ring_norsz\[14\]
rlabel metal1 7130 12104 7130 12104 0 tdc0.w_ring_norsz\[15\]
rlabel metal1 5566 12138 5566 12138 0 tdc0.w_ring_norsz\[16\]
rlabel metal1 15916 12614 15916 12614 0 tdc0.w_ring_norsz\[17\]
rlabel metal1 23828 12274 23828 12274 0 tdc0.w_ring_norsz\[18\]
rlabel metal1 22954 11798 22954 11798 0 tdc0.w_ring_norsz\[19\]
rlabel metal1 16744 12818 16744 12818 0 tdc0.w_ring_norsz\[1\]
rlabel metal2 22218 11424 22218 11424 0 tdc0.w_ring_norsz\[20\]
rlabel metal1 13478 11220 13478 11220 0 tdc0.w_ring_norsz\[21\]
rlabel metal1 10856 12274 10856 12274 0 tdc0.w_ring_norsz\[22\]
rlabel metal1 7728 11322 7728 11322 0 tdc0.w_ring_norsz\[23\]
rlabel metal1 9154 11220 9154 11220 0 tdc0.w_ring_norsz\[24\]
rlabel metal1 17756 11798 17756 11798 0 tdc0.w_ring_norsz\[25\]
rlabel metal1 18952 12138 18952 12138 0 tdc0.w_ring_norsz\[26\]
rlabel metal1 22356 12070 22356 12070 0 tdc0.w_ring_norsz\[27\]
rlabel metal1 18078 11186 18078 11186 0 tdc0.w_ring_norsz\[28\]
rlabel metal1 13708 12410 13708 12410 0 tdc0.w_ring_norsz\[29\]
rlabel metal1 23414 12240 23414 12240 0 tdc0.w_ring_norsz\[2\]
rlabel metal2 12834 12580 12834 12580 0 tdc0.w_ring_norsz\[30\]
rlabel metal1 6532 12138 6532 12138 0 tdc0.w_ring_norsz\[31\]
rlabel metal1 23322 11220 23322 11220 0 tdc0.w_ring_norsz\[3\]
rlabel metal1 20792 10574 20792 10574 0 tdc0.w_ring_norsz\[4\]
rlabel metal1 15042 11322 15042 11322 0 tdc0.w_ring_norsz\[5\]
rlabel metal1 11362 11220 11362 11220 0 tdc0.w_ring_norsz\[6\]
rlabel metal1 6256 11050 6256 11050 0 tdc0.w_ring_norsz\[7\]
rlabel metal1 8924 11050 8924 11050 0 tdc0.w_ring_norsz\[8\]
rlabel metal1 17894 11628 17894 11628 0 tdc0.w_ring_norsz\[9\]
rlabel metal2 12834 7106 12834 7106 0 tdc1.r_dly_store_ctr\[0\]
rlabel metal1 20298 7922 20298 7922 0 tdc1.r_dly_store_ctr\[10\]
rlabel metal2 18262 6902 18262 6902 0 tdc1.r_dly_store_ctr\[11\]
rlabel metal1 20746 5882 20746 5882 0 tdc1.r_dly_store_ctr\[12\]
rlabel metal2 13662 6528 13662 6528 0 tdc1.r_dly_store_ctr\[13\]
rlabel metal1 9292 5746 9292 5746 0 tdc1.r_dly_store_ctr\[14\]
rlabel metal1 8510 7344 8510 7344 0 tdc1.r_dly_store_ctr\[15\]
rlabel metal1 24564 5882 24564 5882 0 tdc1.r_dly_store_ctr\[1\]
rlabel via1 21464 7310 21464 7310 0 tdc1.r_dly_store_ctr\[2\]
rlabel metal1 24978 4794 24978 4794 0 tdc1.r_dly_store_ctr\[3\]
rlabel metal2 26266 5066 26266 5066 0 tdc1.r_dly_store_ctr\[4\]
rlabel metal1 13662 4794 13662 4794 0 tdc1.r_dly_store_ctr\[5\]
rlabel metal1 12788 6222 12788 6222 0 tdc1.r_dly_store_ctr\[6\]
rlabel metal2 9982 6324 9982 6324 0 tdc1.r_dly_store_ctr\[7\]
rlabel metal2 13202 6596 13202 6596 0 tdc1.r_dly_store_ctr\[8\]
rlabel metal1 23690 5882 23690 5882 0 tdc1.r_dly_store_ctr\[9\]
rlabel metal1 4738 8602 4738 8602 0 tdc1.r_dly_store_ring\[0\]
rlabel metal1 29578 9588 29578 9588 0 tdc1.r_dly_store_ring\[10\]
rlabel metal1 30130 7854 30130 7854 0 tdc1.r_dly_store_ring\[11\]
rlabel viali 28842 6834 28842 6834 0 tdc1.r_dly_store_ring\[12\]
rlabel metal1 14674 6732 14674 6732 0 tdc1.r_dly_store_ring\[13\]
rlabel metal1 19688 6970 19688 6970 0 tdc1.r_dly_store_ring\[14\]
rlabel metal1 9338 7922 9338 7922 0 tdc1.r_dly_store_ring\[15\]
rlabel metal2 11362 9095 11362 9095 0 tdc1.r_dly_store_ring\[16\]
rlabel metal1 25760 9146 25760 9146 0 tdc1.r_dly_store_ring\[17\]
rlabel metal1 21666 7344 21666 7344 0 tdc1.r_dly_store_ring\[18\]
rlabel metal1 25392 6970 25392 6970 0 tdc1.r_dly_store_ring\[19\]
rlabel metal1 24610 9894 24610 9894 0 tdc1.r_dly_store_ring\[1\]
rlabel metal1 26358 5882 26358 5882 0 tdc1.r_dly_store_ring\[20\]
rlabel metal1 16698 7888 16698 7888 0 tdc1.r_dly_store_ring\[21\]
rlabel metal1 12190 6120 12190 6120 0 tdc1.r_dly_store_ring\[22\]
rlabel metal1 9982 7990 9982 7990 0 tdc1.r_dly_store_ring\[23\]
rlabel metal2 13110 9214 13110 9214 0 tdc1.r_dly_store_ring\[24\]
rlabel metal1 30314 8602 30314 8602 0 tdc1.r_dly_store_ring\[25\]
rlabel metal1 29394 9486 29394 9486 0 tdc1.r_dly_store_ring\[26\]
rlabel metal2 30406 7752 30406 7752 0 tdc1.r_dly_store_ring\[27\]
rlabel metal1 28934 5882 28934 5882 0 tdc1.r_dly_store_ring\[28\]
rlabel metal1 16560 6426 16560 6426 0 tdc1.r_dly_store_ring\[29\]
rlabel metal1 22540 9146 22540 9146 0 tdc1.r_dly_store_ring\[2\]
rlabel metal1 10258 5848 10258 5848 0 tdc1.r_dly_store_ring\[30\]
rlabel metal1 10350 7174 10350 7174 0 tdc1.r_dly_store_ring\[31\]
rlabel metal2 25714 8228 25714 8228 0 tdc1.r_dly_store_ring\[3\]
rlabel metal1 21160 6426 21160 6426 0 tdc1.r_dly_store_ring\[4\]
rlabel metal1 18124 9690 18124 9690 0 tdc1.r_dly_store_ring\[5\]
rlabel metal2 19090 8313 19090 8313 0 tdc1.r_dly_store_ring\[6\]
rlabel metal1 5842 9146 5842 9146 0 tdc1.r_dly_store_ring\[7\]
rlabel metal1 13570 7990 13570 7990 0 tdc1.r_dly_store_ring\[8\]
rlabel metal1 30498 8942 30498 8942 0 tdc1.r_dly_store_ring\[9\]
rlabel metal1 16606 5746 16606 5746 0 tdc1.r_ring_ctr\[0\]
rlabel metal1 14490 5066 14490 5066 0 tdc1.r_ring_ctr\[10\]
rlabel metal1 17056 5746 17056 5746 0 tdc1.r_ring_ctr\[11\]
rlabel metal1 14214 5236 14214 5236 0 tdc1.r_ring_ctr\[12\]
rlabel metal1 5888 6086 5888 6086 0 tdc1.r_ring_ctr\[13\]
rlabel metal1 5934 6222 5934 6222 0 tdc1.r_ring_ctr\[14\]
rlabel metal1 2714 7242 2714 7242 0 tdc1.r_ring_ctr\[15\]
rlabel metal1 23777 5746 23777 5746 0 tdc1.r_ring_ctr\[1\]
rlabel metal1 21222 4726 21222 4726 0 tdc1.r_ring_ctr\[2\]
rlabel metal1 22494 4726 22494 4726 0 tdc1.r_ring_ctr\[3\]
rlabel metal1 21160 3094 21160 3094 0 tdc1.r_ring_ctr\[4\]
rlabel via1 12461 4658 12461 4658 0 tdc1.r_ring_ctr\[5\]
rlabel metal2 10166 3468 10166 3468 0 tdc1.r_ring_ctr\[6\]
rlabel metal1 8822 5134 8822 5134 0 tdc1.r_ring_ctr\[7\]
rlabel metal2 13938 4896 13938 4896 0 tdc1.r_ring_ctr\[8\]
rlabel metal1 14950 4658 14950 4658 0 tdc1.r_ring_ctr\[9\]
rlabel metal1 26864 5134 26864 5134 0 tdc1.w_dly_stop\[1\]
rlabel metal1 27646 5168 27646 5168 0 tdc1.w_dly_stop\[2\]
rlabel metal1 27324 5134 27324 5134 0 tdc1.w_dly_stop\[3\]
rlabel metal1 27922 5202 27922 5202 0 tdc1.w_dly_stop\[4\]
rlabel via2 15042 6851 15042 6851 0 tdc1.w_dly_stop\[5\]
rlabel metal2 15134 5695 15134 5695 0 tdc1.w_ring_buf\[0\]
rlabel metal1 26864 9690 26864 9690 0 tdc1.w_ring_buf\[10\]
rlabel metal1 28152 7514 28152 7514 0 tdc1.w_ring_buf\[11\]
rlabel metal1 27324 6426 27324 6426 0 tdc1.w_ring_buf\[12\]
rlabel metal2 13570 6630 13570 6630 0 tdc1.w_ring_buf\[13\]
rlabel metal1 18528 6834 18528 6834 0 tdc1.w_ring_buf\[14\]
rlabel metal2 7774 7718 7774 7718 0 tdc1.w_ring_buf\[15\]
rlabel metal1 7436 9078 7436 9078 0 tdc1.w_ring_buf\[16\]
rlabel metal1 24226 9078 24226 9078 0 tdc1.w_ring_buf\[17\]
rlabel metal1 22642 7922 22642 7922 0 tdc1.w_ring_buf\[18\]
rlabel metal1 24104 6426 24104 6426 0 tdc1.w_ring_buf\[19\]
rlabel metal1 23368 9690 23368 9690 0 tdc1.w_ring_buf\[1\]
rlabel metal1 23138 5848 23138 5848 0 tdc1.w_ring_buf\[20\]
rlabel metal1 15727 7310 15727 7310 0 tdc1.w_ring_buf\[21\]
rlabel via1 11081 6222 11081 6222 0 tdc1.w_ring_buf\[22\]
rlabel metal1 9287 8398 9287 8398 0 tdc1.w_ring_buf\[23\]
rlabel metal1 12328 8874 12328 8874 0 tdc1.w_ring_buf\[24\]
rlabel metal1 28872 8330 28872 8330 0 tdc1.w_ring_buf\[25\]
rlabel metal1 27784 9690 27784 9690 0 tdc1.w_ring_buf\[26\]
rlabel metal1 28826 7242 28826 7242 0 tdc1.w_ring_buf\[27\]
rlabel metal1 27446 5814 27446 5814 0 tdc1.w_ring_buf\[28\]
rlabel metal1 15394 6154 15394 6154 0 tdc1.w_ring_buf\[29\]
rlabel metal2 21206 8806 21206 8806 0 tdc1.w_ring_buf\[2\]
rlabel metal1 8862 6154 8862 6154 0 tdc1.w_ring_buf\[30\]
rlabel metal1 8172 7242 8172 7242 0 tdc1.w_ring_buf\[31\]
rlabel metal2 24426 7718 24426 7718 0 tdc1.w_ring_buf\[3\]
rlabel via1 20373 6222 20373 6222 0 tdc1.w_ring_buf\[4\]
rlabel metal2 17710 9282 17710 9282 0 tdc1.w_ring_buf\[5\]
rlabel metal2 17710 8194 17710 8194 0 tdc1.w_ring_buf\[6\]
rlabel metal2 5014 8806 5014 8806 0 tdc1.w_ring_buf\[7\]
rlabel metal2 12558 8126 12558 8126 0 tdc1.w_ring_buf\[8\]
rlabel metal1 28412 9078 28412 9078 0 tdc1.w_ring_buf\[9\]
rlabel metal1 6716 7514 6716 7514 0 tdc1.w_ring_int_norsz\[0\]
rlabel metal1 27186 9078 27186 9078 0 tdc1.w_ring_int_norsz\[10\]
rlabel metal1 27094 7990 27094 7990 0 tdc1.w_ring_int_norsz\[11\]
rlabel metal1 27002 6766 27002 6766 0 tdc1.w_ring_int_norsz\[12\]
rlabel metal1 19366 6664 19366 6664 0 tdc1.w_ring_int_norsz\[13\]
rlabel metal1 13156 6426 13156 6426 0 tdc1.w_ring_int_norsz\[14\]
rlabel metal1 7912 6766 7912 6766 0 tdc1.w_ring_int_norsz\[15\]
rlabel metal1 6578 8364 6578 8364 0 tdc1.w_ring_int_norsz\[16\]
rlabel via2 7406 8347 7406 8347 0 tdc1.w_ring_int_norsz\[17\]
rlabel metal1 24242 8330 24242 8330 0 tdc1.w_ring_int_norsz\[18\]
rlabel metal1 24104 7378 24104 7378 0 tdc1.w_ring_int_norsz\[19\]
rlabel metal1 22770 8330 22770 8330 0 tdc1.w_ring_int_norsz\[1\]
rlabel metal2 23506 6596 23506 6596 0 tdc1.w_ring_int_norsz\[20\]
rlabel metal1 19274 6188 19274 6188 0 tdc1.w_ring_int_norsz\[21\]
rlabel metal1 17204 6970 17204 6970 0 tdc1.w_ring_int_norsz\[22\]
rlabel metal1 11638 7514 11638 7514 0 tdc1.w_ring_int_norsz\[23\]
rlabel metal1 11914 8500 11914 8500 0 tdc1.w_ring_int_norsz\[24\]
rlabel metal1 23966 9044 23966 9044 0 tdc1.w_ring_int_norsz\[25\]
rlabel metal1 27876 8602 27876 8602 0 tdc1.w_ring_int_norsz\[26\]
rlabel metal1 27738 7956 27738 7956 0 tdc1.w_ring_int_norsz\[27\]
rlabel metal1 26082 6902 26082 6902 0 tdc1.w_ring_int_norsz\[28\]
rlabel metal1 24058 6120 24058 6120 0 tdc1.w_ring_int_norsz\[29\]
rlabel metal1 23138 8058 23138 8058 0 tdc1.w_ring_int_norsz\[2\]
rlabel metal1 14398 6154 14398 6154 0 tdc1.w_ring_int_norsz\[30\]
rlabel metal1 8510 6766 8510 6766 0 tdc1.w_ring_int_norsz\[31\]
rlabel metal1 23690 7378 23690 7378 0 tdc1.w_ring_int_norsz\[3\]
rlabel metal1 23276 6766 23276 6766 0 tdc1.w_ring_int_norsz\[4\]
rlabel metal1 18446 6902 18446 6902 0 tdc1.w_ring_int_norsz\[5\]
rlabel metal1 17480 7378 17480 7378 0 tdc1.w_ring_int_norsz\[6\]
rlabel metal1 16560 7514 16560 7514 0 tdc1.w_ring_int_norsz\[7\]
rlabel metal1 11316 8330 11316 8330 0 tdc1.w_ring_int_norsz\[8\]
rlabel metal1 19734 8364 19734 8364 0 tdc1.w_ring_int_norsz\[9\]
rlabel metal1 13294 8840 13294 8840 0 tdc1.w_ring_norsz\[0\]
rlabel metal2 26910 8942 26910 8942 0 tdc1.w_ring_norsz\[10\]
rlabel metal1 27324 7718 27324 7718 0 tdc1.w_ring_norsz\[11\]
rlabel metal1 27002 6630 27002 6630 0 tdc1.w_ring_norsz\[12\]
rlabel metal1 18952 6358 18952 6358 0 tdc1.w_ring_norsz\[13\]
rlabel metal1 12834 6732 12834 6732 0 tdc1.w_ring_norsz\[14\]
rlabel metal1 8004 6834 8004 6834 0 tdc1.w_ring_norsz\[15\]
rlabel metal1 6762 9044 6762 9044 0 tdc1.w_ring_norsz\[16\]
rlabel metal1 23874 8908 23874 8908 0 tdc1.w_ring_norsz\[17\]
rlabel metal2 24058 8092 24058 8092 0 tdc1.w_ring_norsz\[18\]
rlabel metal1 23644 7446 23644 7446 0 tdc1.w_ring_norsz\[19\]
rlabel metal2 23046 9248 23046 9248 0 tdc1.w_ring_norsz\[1\]
rlabel metal1 23092 6698 23092 6698 0 tdc1.w_ring_norsz\[20\]
rlabel metal1 17572 6970 17572 6970 0 tdc1.w_ring_norsz\[21\]
rlabel metal1 16882 7242 16882 7242 0 tdc1.w_ring_norsz\[22\]
rlabel metal1 10350 8398 10350 8398 0 tdc1.w_ring_norsz\[23\]
rlabel metal1 12512 8398 12512 8398 0 tdc1.w_ring_norsz\[24\]
rlabel metal1 26956 8874 26956 8874 0 tdc1.w_ring_norsz\[25\]
rlabel metal1 27462 8840 27462 8840 0 tdc1.w_ring_norsz\[26\]
rlabel metal1 26910 7786 26910 7786 0 tdc1.w_ring_norsz\[27\]
rlabel metal2 26726 6222 26726 6222 0 tdc1.w_ring_norsz\[28\]
rlabel metal1 18814 6188 18814 6188 0 tdc1.w_ring_norsz\[29\]
rlabel metal1 21022 8432 21022 8432 0 tdc1.w_ring_norsz\[2\]
rlabel metal1 13662 6392 13662 6392 0 tdc1.w_ring_norsz\[30\]
rlabel metal1 7728 6698 7728 6698 0 tdc1.w_ring_norsz\[31\]
rlabel metal1 24242 7276 24242 7276 0 tdc1.w_ring_norsz\[3\]
rlabel metal1 20102 6800 20102 6800 0 tdc1.w_ring_norsz\[4\]
rlabel metal2 17802 8160 17802 8160 0 tdc1.w_ring_norsz\[5\]
rlabel metal1 17434 7514 17434 7514 0 tdc1.w_ring_norsz\[6\]
rlabel metal1 10994 8364 10994 8364 0 tdc1.w_ring_norsz\[7\]
rlabel metal1 12742 8432 12742 8432 0 tdc1.w_ring_norsz\[8\]
rlabel metal1 27094 9520 27094 9520 0 tdc1.w_ring_norsz\[9\]
rlabel metal2 31050 7701 31050 7701 0 ui_in[0]
rlabel metal3 590 14348 590 14348 0 ui_in[1]
rlabel metal3 590 10268 590 10268 0 ui_in[2]
rlabel metal2 16790 568 16790 568 0 ui_in[3]
rlabel metal2 16245 340 16245 340 0 ui_in[4]
rlabel metal2 15502 415 15502 415 0 ui_in[5]
rlabel metal2 13570 9146 13570 9146 0 uo_out[0]
rlabel metal3 28804 9588 28804 9588 0 uo_out[1]
rlabel metal2 27278 11985 27278 11985 0 uo_out[2]
rlabel via2 31702 10268 31702 10268 0 uo_out[3]
rlabel metal2 22770 7021 22770 7021 0 uo_out[4]
rlabel metal1 15962 9622 15962 9622 0 uo_out[5]
rlabel metal2 12650 14008 12650 14008 0 uo_out[6]
rlabel metal2 10074 9537 10074 9537 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
