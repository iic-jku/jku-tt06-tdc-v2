magic
tech sky130A
magscale 1 2
timestamp 1711751087
<< viali >>
rect 14657 12393 14691 12427
rect 14933 12393 14967 12427
rect 17877 12393 17911 12427
rect 20085 12393 20119 12427
rect 20545 12393 20579 12427
rect 12449 12325 12483 12359
rect 14841 12325 14875 12359
rect 20269 12325 20303 12359
rect 13533 12257 13567 12291
rect 18337 12257 18371 12291
rect 18961 12257 18995 12291
rect 13277 12189 13311 12223
rect 16129 12189 16163 12223
rect 16405 12189 16439 12223
rect 18245 12189 18279 12223
rect 18705 12189 18739 12223
rect 17969 12121 18003 12155
rect 12541 12053 12575 12087
rect 12265 11849 12299 11883
rect 13829 11849 13863 11883
rect 16681 11849 16715 11883
rect 18153 11849 18187 11883
rect 18797 11849 18831 11883
rect 14657 11713 14691 11747
rect 16405 11713 16439 11747
rect 17509 11713 17543 11747
rect 17969 11713 18003 11747
rect 11345 11645 11379 11679
rect 11621 11645 11655 11679
rect 12725 11645 12759 11679
rect 13093 11645 13127 11679
rect 14105 11645 14139 11679
rect 16589 11645 16623 11679
rect 17325 11645 17359 11679
rect 17785 11645 17819 11679
rect 18061 11645 18095 11679
rect 18245 11645 18279 11679
rect 19073 11645 19107 11679
rect 19441 11645 19475 11679
rect 11989 11577 12023 11611
rect 14933 11577 14967 11611
rect 17141 11577 17175 11611
rect 19686 11577 19720 11611
rect 21005 11577 21039 11611
rect 21373 11577 21407 11611
rect 11529 11509 11563 11543
rect 11805 11509 11839 11543
rect 17601 11509 17635 11543
rect 20821 11509 20855 11543
rect 14013 11305 14047 11339
rect 14289 11305 14323 11339
rect 15025 11305 15059 11339
rect 15669 11305 15703 11339
rect 19717 11305 19751 11339
rect 14197 11237 14231 11271
rect 18245 11237 18279 11271
rect 19625 11237 19659 11271
rect 10977 11169 11011 11203
rect 11244 11169 11278 11203
rect 12633 11169 12667 11203
rect 12900 11169 12934 11203
rect 15209 11169 15243 11203
rect 15577 11169 15611 11203
rect 16681 11169 16715 11203
rect 17141 11169 17175 11203
rect 18613 11169 18647 11203
rect 20085 11169 20119 11203
rect 12357 10965 12391 10999
rect 16773 10965 16807 10999
rect 17049 10965 17083 10999
rect 10885 10761 10919 10795
rect 11345 10761 11379 10795
rect 11897 10761 11931 10795
rect 12909 10761 12943 10795
rect 13737 10761 13771 10795
rect 20361 10761 20395 10795
rect 15945 10625 15979 10659
rect 16221 10625 16255 10659
rect 17693 10625 17727 10659
rect 11161 10557 11195 10591
rect 11529 10557 11563 10591
rect 12173 10557 12207 10591
rect 12725 10557 12759 10591
rect 13185 10557 13219 10591
rect 13921 10557 13955 10591
rect 14013 10557 14047 10591
rect 18705 10557 18739 10591
rect 18961 10557 18995 10591
rect 20269 10489 20303 10523
rect 12541 10421 12575 10455
rect 20085 10421 20119 10455
rect 10793 10217 10827 10251
rect 11161 10217 11195 10251
rect 12265 10217 12299 10251
rect 13277 10217 13311 10251
rect 14289 10217 14323 10251
rect 15761 10217 15795 10251
rect 16313 10217 16347 10251
rect 18061 10217 18095 10251
rect 18337 10217 18371 10251
rect 20729 10217 20763 10251
rect 11069 10149 11103 10183
rect 14626 10149 14660 10183
rect 16221 10149 16255 10183
rect 18245 10149 18279 10183
rect 21373 10149 21407 10183
rect 9413 10081 9447 10115
rect 9680 10081 9714 10115
rect 11621 10081 11655 10115
rect 11805 10081 11839 10115
rect 12449 10081 12483 10115
rect 12817 10081 12851 10115
rect 13185 10081 13219 10115
rect 13461 10081 13495 10115
rect 14105 10081 14139 10115
rect 16937 10081 16971 10115
rect 19605 10081 19639 10115
rect 21741 10081 21775 10115
rect 12541 10013 12575 10047
rect 12725 10013 12759 10047
rect 12909 10013 12943 10047
rect 14381 10013 14415 10047
rect 16681 10013 16715 10047
rect 19349 10013 19383 10047
rect 11805 9945 11839 9979
rect 12081 9945 12115 9979
rect 13093 9945 13127 9979
rect 13185 9945 13219 9979
rect 12817 9877 12851 9911
rect 14013 9877 14047 9911
rect 10333 9673 10367 9707
rect 11621 9673 11655 9707
rect 11897 9673 11931 9707
rect 12357 9673 12391 9707
rect 12725 9673 12759 9707
rect 13001 9673 13035 9707
rect 16037 9673 16071 9707
rect 16681 9673 16715 9707
rect 14013 9605 14047 9639
rect 14105 9605 14139 9639
rect 14289 9605 14323 9639
rect 16221 9605 16255 9639
rect 17049 9605 17083 9639
rect 19073 9605 19107 9639
rect 11989 9537 12023 9571
rect 12449 9537 12483 9571
rect 12633 9537 12667 9571
rect 9781 9469 9815 9503
rect 10149 9469 10183 9503
rect 10517 9469 10551 9503
rect 11437 9469 11471 9503
rect 11621 9469 11655 9503
rect 11719 9469 11753 9503
rect 11897 9469 11931 9503
rect 12541 9469 12575 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 13001 9469 13035 9503
rect 13185 9469 13219 9503
rect 13553 9469 13587 9503
rect 13737 9469 13771 9503
rect 14105 9469 14139 9503
rect 14197 9469 14231 9503
rect 14657 9469 14691 9503
rect 15209 9469 15243 9503
rect 15393 9469 15427 9503
rect 15669 9469 15703 9503
rect 15945 9469 15979 9503
rect 16037 9469 16071 9503
rect 16129 9469 16163 9503
rect 16405 9469 16439 9503
rect 16497 9469 16531 9503
rect 17325 9469 17359 9503
rect 17509 9469 17543 9503
rect 17785 9469 17819 9503
rect 18889 9469 18923 9503
rect 19533 9469 19567 9503
rect 19901 9469 19935 9503
rect 12265 9401 12299 9435
rect 13645 9401 13679 9435
rect 13829 9401 13863 9435
rect 14473 9401 14507 9435
rect 15301 9401 15335 9435
rect 15761 9401 15795 9435
rect 16865 9401 16899 9435
rect 17417 9401 17451 9435
rect 20085 9401 20119 9435
rect 20453 9401 20487 9435
rect 14197 9333 14231 9367
rect 14749 9333 14783 9367
rect 16129 9333 16163 9367
rect 17969 9333 18003 9367
rect 9321 9129 9355 9163
rect 10793 9129 10827 9163
rect 12357 9129 12391 9163
rect 12449 9129 12483 9163
rect 14381 9129 14415 9163
rect 19717 9129 19751 9163
rect 9658 9061 9692 9095
rect 11069 9061 11103 9095
rect 15853 9061 15887 9095
rect 16497 9061 16531 9095
rect 17877 9061 17911 9095
rect 18582 9061 18616 9095
rect 9137 8993 9171 9027
rect 9413 8993 9447 9027
rect 11805 8993 11839 9027
rect 11989 8993 12023 9027
rect 12357 8993 12391 9027
rect 12449 8993 12483 9027
rect 12817 8993 12851 9027
rect 13001 8993 13035 9027
rect 13093 8993 13127 9027
rect 14289 8993 14323 9027
rect 14473 8993 14507 9027
rect 15761 8993 15795 9027
rect 15945 8993 15979 9027
rect 16129 8993 16163 9027
rect 16221 8993 16255 9027
rect 16681 8993 16715 9027
rect 16773 8993 16807 9027
rect 17049 8993 17083 9027
rect 17141 8993 17175 9027
rect 17325 8993 17359 9027
rect 17417 8993 17451 9027
rect 21373 8993 21407 9027
rect 11897 8925 11931 8959
rect 12081 8925 12115 8959
rect 12725 8925 12759 8959
rect 12909 8925 12943 8959
rect 16405 8925 16439 8959
rect 17233 8925 17267 8959
rect 18337 8925 18371 8959
rect 12265 8857 12299 8891
rect 12541 8857 12575 8891
rect 16773 8857 16807 8891
rect 11161 8789 11195 8823
rect 13461 8789 13495 8823
rect 15025 8789 15059 8823
rect 16313 8789 16347 8823
rect 17601 8789 17635 8823
rect 18153 8789 18187 8823
rect 21649 8789 21683 8823
rect 9597 8585 9631 8619
rect 13093 8585 13127 8619
rect 13553 8585 13587 8619
rect 13921 8585 13955 8619
rect 15025 8585 15059 8619
rect 20821 8585 20855 8619
rect 15117 8517 15151 8551
rect 13185 8449 13219 8483
rect 13829 8449 13863 8483
rect 14657 8449 14691 8483
rect 19441 8449 19475 8483
rect 9781 8381 9815 8415
rect 10057 8381 10091 8415
rect 10701 8381 10735 8415
rect 11897 8381 11931 8415
rect 13093 8381 13127 8415
rect 13553 8381 13587 8415
rect 13645 8381 13679 8415
rect 13927 8381 13961 8415
rect 14105 8381 14139 8415
rect 14289 8381 14323 8415
rect 14473 8381 14507 8415
rect 14565 8381 14599 8415
rect 14841 8381 14875 8415
rect 15209 8381 15243 8415
rect 15301 8381 15335 8415
rect 15485 8381 15519 8415
rect 16405 8381 16439 8415
rect 18337 8381 18371 8415
rect 18705 8381 18739 8415
rect 10425 8313 10459 8347
rect 13369 8313 13403 8347
rect 14381 8313 14415 8347
rect 14933 8313 14967 8347
rect 17969 8313 18003 8347
rect 19686 8313 19720 8347
rect 10517 8245 10551 8279
rect 11713 8245 11747 8279
rect 14565 8245 14599 8279
rect 15393 8245 15427 8279
rect 16589 8245 16623 8279
rect 18889 8245 18923 8279
rect 12633 8041 12667 8075
rect 13461 8041 13495 8075
rect 14933 8041 14967 8075
rect 18153 8041 18187 8075
rect 20177 8041 20211 8075
rect 9680 7973 9714 8007
rect 11520 7973 11554 8007
rect 12817 7973 12851 8007
rect 15209 7973 15243 8007
rect 17018 7973 17052 8007
rect 18337 7973 18371 8007
rect 19042 7973 19076 8007
rect 20361 7973 20395 8007
rect 9413 7905 9447 7939
rect 11253 7905 11287 7939
rect 13369 7905 13403 7939
rect 13553 7905 13587 7939
rect 13645 7905 13679 7939
rect 14749 7905 14783 7939
rect 15669 7905 15703 7939
rect 18797 7905 18831 7939
rect 16773 7837 16807 7871
rect 15853 7769 15887 7803
rect 10793 7701 10827 7735
rect 12909 7701 12943 7735
rect 13829 7701 13863 7735
rect 15485 7701 15519 7735
rect 18429 7701 18463 7735
rect 20637 7701 20671 7735
rect 9781 7497 9815 7531
rect 15025 7361 15059 7395
rect 10057 7293 10091 7327
rect 10793 7293 10827 7327
rect 11713 7293 11747 7327
rect 13553 7293 13587 7327
rect 13820 7293 13854 7327
rect 15292 7293 15326 7327
rect 16957 7293 16991 7327
rect 18981 7293 19015 7327
rect 19349 7225 19383 7259
rect 10885 7157 10919 7191
rect 11805 7157 11839 7191
rect 14933 7157 14967 7191
rect 16405 7157 16439 7191
rect 17049 7157 17083 7191
rect 13829 6885 13863 6919
rect 14933 6885 14967 6919
rect 16589 6885 16623 6919
rect 13921 6613 13955 6647
rect 15025 6613 15059 6647
rect 16681 6613 16715 6647
rect 12633 901 12667 935
rect 10057 833 10091 867
rect 9781 765 9815 799
rect 12449 697 12483 731
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12393 14703 12427
rect 14645 12387 14703 12393
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 14660 12356 14688 12387
rect 14918 12384 14924 12436
rect 14976 12384 14982 12436
rect 17865 12427 17923 12433
rect 17865 12393 17877 12427
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20533 12427 20591 12433
rect 20119 12396 20300 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 14829 12359 14887 12365
rect 14829 12356 14841 12359
rect 12492 12328 13676 12356
rect 14660 12328 14841 12356
rect 12492 12316 12498 12328
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 13521 12291 13579 12297
rect 13521 12288 13533 12291
rect 13412 12260 13533 12288
rect 13412 12248 13418 12260
rect 13521 12257 13533 12260
rect 13567 12257 13579 12291
rect 13648 12288 13676 12328
rect 14829 12325 14841 12328
rect 14875 12325 14887 12359
rect 14829 12319 14887 12325
rect 15470 12316 15476 12368
rect 15528 12316 15534 12368
rect 16850 12316 16856 12368
rect 16908 12316 16914 12368
rect 15488 12288 15516 12316
rect 13648 12260 15516 12288
rect 17880 12288 17908 12387
rect 20272 12365 20300 12396
rect 20533 12393 20545 12427
rect 20579 12424 20591 12427
rect 20622 12424 20628 12436
rect 20579 12396 20628 12424
rect 20579 12393 20591 12396
rect 20533 12387 20591 12393
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 20257 12359 20315 12365
rect 20257 12325 20269 12359
rect 20303 12325 20315 12359
rect 20257 12319 20315 12325
rect 18966 12297 18972 12300
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 17880 12260 18337 12288
rect 13521 12251 13579 12257
rect 18325 12257 18337 12260
rect 18371 12288 18383 12291
rect 18949 12291 18972 12297
rect 18949 12288 18961 12291
rect 18371 12260 18961 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 18949 12257 18961 12260
rect 18949 12251 18972 12257
rect 18966 12248 18972 12251
rect 19024 12248 19030 12300
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12768 12192 13277 12220
rect 12768 12180 12774 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 16114 12180 16120 12232
rect 16172 12180 16178 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16439 12192 18000 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 17972 12161 18000 12192
rect 18230 12180 18236 12232
rect 18288 12180 18294 12232
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 17957 12155 18015 12161
rect 17957 12121 17969 12155
rect 18003 12121 18015 12155
rect 17957 12115 18015 12121
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12618 12084 12624 12096
rect 12575 12056 12624 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 18708 12084 18736 12183
rect 19058 12084 19064 12096
rect 18708 12056 19064 12084
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12434 11880 12440 11892
rect 12299 11852 12440 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13817 11883 13875 11889
rect 13817 11880 13829 11883
rect 13596 11852 13829 11880
rect 13596 11840 13602 11852
rect 13817 11849 13829 11852
rect 13863 11849 13875 11883
rect 13817 11843 13875 11849
rect 16669 11883 16727 11889
rect 16669 11849 16681 11883
rect 16715 11880 16727 11883
rect 16850 11880 16856 11892
rect 16715 11852 16856 11880
rect 16715 11849 16727 11852
rect 16669 11843 16727 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11880 18199 11883
rect 18230 11880 18236 11892
rect 18187 11852 18236 11880
rect 18187 11849 18199 11852
rect 18141 11843 18199 11849
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 18782 11840 18788 11892
rect 18840 11840 18846 11892
rect 18966 11840 18972 11892
rect 19024 11840 19030 11892
rect 17328 11784 18920 11812
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11744 14703 11747
rect 16114 11744 16120 11756
rect 14691 11716 16120 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11645 11391 11679
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 11333 11639 11391 11645
rect 11532 11648 11621 11676
rect 11348 11552 11376 11639
rect 11330 11500 11336 11552
rect 11388 11500 11394 11552
rect 11532 11549 11560 11648
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 12676 11648 12725 11676
rect 12676 11636 12682 11648
rect 12713 11645 12725 11648
rect 12759 11676 12771 11679
rect 13081 11679 13139 11685
rect 13081 11676 13093 11679
rect 12759 11648 13093 11676
rect 12759 11645 12771 11648
rect 12713 11639 12771 11645
rect 13081 11645 13093 11648
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 11977 11611 12035 11617
rect 11977 11577 11989 11611
rect 12023 11577 12035 11611
rect 11977 11571 12035 11577
rect 11517 11543 11575 11549
rect 11517 11509 11529 11543
rect 11563 11509 11575 11543
rect 11517 11503 11575 11509
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 11992 11540 12020 11571
rect 11839 11512 12020 11540
rect 13096 11540 13124 11639
rect 13354 11636 13360 11688
rect 13412 11676 13418 11688
rect 13722 11676 13728 11688
rect 13412 11648 13728 11676
rect 13412 11636 13418 11648
rect 13722 11636 13728 11648
rect 13780 11676 13786 11688
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 13780 11648 14105 11676
rect 13780 11636 13786 11648
rect 14093 11645 14105 11648
rect 14139 11676 14151 11679
rect 14660 11676 14688 11707
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11744 16451 11747
rect 17328 11744 17356 11784
rect 16439 11716 17356 11744
rect 16439 11713 16451 11716
rect 16393 11707 16451 11713
rect 14139 11648 14688 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 16574 11636 16580 11688
rect 16632 11636 16638 11688
rect 17328 11685 17356 11716
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11744 17555 11747
rect 17957 11747 18015 11753
rect 17957 11744 17969 11747
rect 17543 11716 17969 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 17957 11713 17969 11716
rect 18003 11713 18015 11747
rect 17957 11707 18015 11713
rect 18064 11685 18092 11784
rect 17313 11679 17371 11685
rect 17313 11645 17325 11679
rect 17359 11645 17371 11679
rect 17313 11639 17371 11645
rect 17773 11679 17831 11685
rect 17773 11645 17785 11679
rect 17819 11645 17831 11679
rect 17773 11639 17831 11645
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 14918 11568 14924 11620
rect 14976 11568 14982 11620
rect 15654 11568 15660 11620
rect 15712 11568 15718 11620
rect 16592 11608 16620 11636
rect 16224 11580 16620 11608
rect 16224 11540 16252 11580
rect 17126 11568 17132 11620
rect 17184 11568 17190 11620
rect 17788 11608 17816 11639
rect 18138 11636 18144 11688
rect 18196 11636 18202 11688
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18279 11648 18828 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18156 11608 18184 11636
rect 17788 11580 18184 11608
rect 18800 11552 18828 11648
rect 18892 11608 18920 11784
rect 18984 11676 19012 11840
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 18984 11648 19073 11676
rect 19061 11645 19073 11648
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 19300 11648 19441 11676
rect 19300 11636 19306 11648
rect 19429 11645 19441 11648
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 19610 11608 19616 11620
rect 18892 11580 19616 11608
rect 19610 11568 19616 11580
rect 19668 11617 19674 11620
rect 19668 11611 19732 11617
rect 19668 11577 19686 11611
rect 19720 11577 19732 11611
rect 20993 11611 21051 11617
rect 20993 11608 21005 11611
rect 19668 11571 19732 11577
rect 20824 11580 21005 11608
rect 19668 11568 19674 11571
rect 13096 11512 16252 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 17586 11500 17592 11552
rect 17644 11500 17650 11552
rect 18782 11500 18788 11552
rect 18840 11500 18846 11552
rect 20824 11549 20852 11580
rect 20993 11577 21005 11580
rect 21039 11577 21051 11611
rect 20993 11571 21051 11577
rect 21361 11611 21419 11617
rect 21361 11577 21373 11611
rect 21407 11608 21419 11611
rect 28258 11608 28264 11620
rect 21407 11580 28264 11608
rect 21407 11577 21419 11580
rect 21361 11571 21419 11577
rect 28258 11568 28264 11580
rect 28316 11568 28322 11620
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11509 20867 11543
rect 20809 11503 20867 11509
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 14001 11339 14059 11345
rect 14001 11305 14013 11339
rect 14047 11305 14059 11339
rect 14001 11299 14059 11305
rect 11330 11268 11336 11280
rect 10980 11240 11336 11268
rect 10980 11209 11008 11240
rect 11330 11228 11336 11240
rect 11388 11268 11394 11280
rect 14016 11268 14044 11299
rect 14274 11296 14280 11348
rect 14332 11296 14338 11348
rect 14918 11296 14924 11348
rect 14976 11336 14982 11348
rect 15013 11339 15071 11345
rect 15013 11336 15025 11339
rect 14976 11308 15025 11336
rect 14976 11296 14982 11308
rect 15013 11305 15025 11308
rect 15059 11305 15071 11339
rect 15013 11299 15071 11305
rect 15654 11296 15660 11348
rect 15712 11296 15718 11348
rect 17586 11296 17592 11348
rect 17644 11296 17650 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19392 11308 19717 11336
rect 19392 11296 19398 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 14185 11271 14243 11277
rect 14185 11268 14197 11271
rect 11388 11240 12434 11268
rect 14016 11240 14197 11268
rect 11388 11228 11394 11240
rect 11238 11209 11244 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11232 11163 11244 11209
rect 10980 11064 11008 11163
rect 11238 11160 11244 11163
rect 11296 11160 11302 11212
rect 12406 11200 12434 11240
rect 14185 11237 14197 11240
rect 14231 11237 14243 11271
rect 17604 11268 17632 11296
rect 14185 11231 14243 11237
rect 15212 11240 17632 11268
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12406 11172 12633 11200
rect 12621 11169 12633 11172
rect 12667 11200 12679 11203
rect 12710 11200 12716 11212
rect 12667 11172 12716 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 12888 11203 12946 11209
rect 12888 11169 12900 11203
rect 12934 11200 12946 11203
rect 13170 11200 13176 11212
rect 12934 11172 13176 11200
rect 12934 11169 12946 11172
rect 12888 11163 12946 11169
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 15212 11209 15240 11240
rect 17678 11228 17684 11280
rect 17736 11268 17742 11280
rect 18233 11271 18291 11277
rect 18233 11268 18245 11271
rect 17736 11240 18245 11268
rect 17736 11228 17742 11240
rect 18233 11237 18245 11240
rect 18279 11237 18291 11271
rect 18233 11231 18291 11237
rect 19610 11228 19616 11280
rect 19668 11228 19674 11280
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11169 15255 11203
rect 15197 11163 15255 11169
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 16574 11200 16580 11212
rect 15611 11172 16580 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 16684 11132 16712 11163
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 17184 11172 18613 11200
rect 17184 11160 17190 11172
rect 18601 11169 18613 11172
rect 18647 11200 18659 11203
rect 18647 11172 18828 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 16592 11104 16712 11132
rect 16592 11076 16620 11104
rect 9600 11036 11008 11064
rect 9600 11008 9628 11036
rect 16574 11024 16580 11076
rect 16632 11024 16638 11076
rect 18800 11008 18828 11172
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 20073 11203 20131 11209
rect 20073 11200 20085 11203
rect 19392 11172 20085 11200
rect 19392 11160 19398 11172
rect 20073 11169 20085 11172
rect 20119 11169 20131 11203
rect 20073 11163 20131 11169
rect 9582 10956 9588 11008
rect 9640 10956 9646 11008
rect 12342 10956 12348 11008
rect 12400 10956 12406 11008
rect 16758 10956 16764 11008
rect 16816 10956 16822 11008
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 17037 10999 17095 11005
rect 17037 10996 17049 10999
rect 16908 10968 17049 10996
rect 16908 10956 16914 10968
rect 17037 10965 17049 10968
rect 17083 10965 17095 10999
rect 17037 10959 17095 10965
rect 18782 10956 18788 11008
rect 18840 10956 18846 11008
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 10870 10752 10876 10804
rect 10928 10752 10934 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 11296 10764 11345 10792
rect 11296 10752 11302 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11480 10764 11897 10792
rect 11480 10752 11486 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 12894 10752 12900 10804
rect 12952 10752 12958 10804
rect 13722 10752 13728 10804
rect 13780 10752 13786 10804
rect 16206 10792 16212 10804
rect 15948 10764 16212 10792
rect 11149 10591 11207 10597
rect 11149 10557 11161 10591
rect 11195 10588 11207 10591
rect 11256 10588 11284 10752
rect 14550 10656 14556 10668
rect 12452 10628 14556 10656
rect 12452 10600 12480 10628
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 15948 10665 15976 10764
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 19978 10752 19984 10804
rect 20036 10792 20042 10804
rect 20349 10795 20407 10801
rect 20349 10792 20361 10795
rect 20036 10764 20361 10792
rect 20036 10752 20042 10764
rect 20349 10761 20361 10764
rect 20395 10761 20407 10795
rect 20349 10755 20407 10761
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16209 10659 16267 10665
rect 16209 10625 16221 10659
rect 16255 10656 16267 10659
rect 16850 10656 16856 10668
rect 16255 10628 16856 10656
rect 16255 10625 16267 10628
rect 16209 10619 16267 10625
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10656 17739 10659
rect 17727 10628 18828 10656
rect 17727 10625 17739 10628
rect 17681 10619 17739 10625
rect 18800 10600 18828 10628
rect 11195 10560 11284 10588
rect 11517 10591 11575 10597
rect 11195 10557 11207 10560
rect 11149 10551 11207 10557
rect 11517 10557 11529 10591
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12342 10588 12348 10600
rect 12207 10560 12348 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 11532 10520 11560 10551
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12434 10548 12440 10600
rect 12492 10548 12498 10600
rect 12526 10548 12532 10600
rect 12584 10548 12590 10600
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 12676 10560 12725 10588
rect 12676 10548 12682 10560
rect 12713 10557 12725 10560
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 13170 10548 13176 10600
rect 13228 10548 13234 10600
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13464 10560 13921 10588
rect 12544 10520 12572 10548
rect 13464 10532 13492 10560
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10557 14059 10591
rect 14001 10551 14059 10557
rect 11532 10492 12572 10520
rect 13446 10480 13452 10532
rect 13504 10480 13510 10532
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12529 10455 12587 10461
rect 12529 10452 12541 10455
rect 12492 10424 12541 10452
rect 12492 10412 12498 10424
rect 12529 10421 12541 10424
rect 12575 10421 12587 10455
rect 12529 10415 12587 10421
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 14016 10452 14044 10551
rect 18690 10548 18696 10600
rect 18748 10548 18754 10600
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 18949 10591 19007 10597
rect 18949 10588 18961 10591
rect 18840 10560 18961 10588
rect 18840 10548 18846 10560
rect 18949 10557 18961 10560
rect 18995 10557 19007 10591
rect 18949 10551 19007 10557
rect 16758 10480 16764 10532
rect 16816 10480 16822 10532
rect 20257 10523 20315 10529
rect 20257 10520 20269 10523
rect 20088 10492 20269 10520
rect 20088 10461 20116 10492
rect 20257 10489 20269 10492
rect 20303 10489 20315 10523
rect 20257 10483 20315 10489
rect 13044 10424 14044 10452
rect 20073 10455 20131 10461
rect 13044 10412 13050 10424
rect 20073 10421 20085 10455
rect 20119 10421 20131 10455
rect 20073 10415 20131 10421
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 10781 10251 10839 10257
rect 10781 10217 10793 10251
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 9582 10140 9588 10192
rect 9640 10140 9646 10192
rect 10796 10180 10824 10211
rect 11146 10208 11152 10260
rect 11204 10208 11210 10260
rect 12253 10251 12311 10257
rect 12253 10217 12265 10251
rect 12299 10248 12311 10251
rect 12299 10220 13124 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 11057 10183 11115 10189
rect 11057 10180 11069 10183
rect 10796 10152 11069 10180
rect 11057 10149 11069 10152
rect 11103 10149 11115 10183
rect 12986 10180 12992 10192
rect 11057 10143 11115 10149
rect 11808 10152 12992 10180
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 9600 10112 9628 10140
rect 9456 10084 9628 10112
rect 9668 10115 9726 10121
rect 9456 10072 9462 10084
rect 9668 10081 9680 10115
rect 9714 10112 9726 10115
rect 10042 10112 10048 10124
rect 9714 10084 10048 10112
rect 9714 10081 9726 10084
rect 9668 10075 9726 10081
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 11808 10121 11836 10152
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 13096 10124 13124 10220
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 13265 10251 13323 10257
rect 13265 10248 13277 10251
rect 13228 10220 13277 10248
rect 13228 10208 13234 10220
rect 13265 10217 13277 10220
rect 13311 10217 13323 10251
rect 13265 10211 13323 10217
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 15749 10251 15807 10257
rect 15749 10217 15761 10251
rect 15795 10217 15807 10251
rect 15749 10211 15807 10217
rect 14292 10180 14320 10211
rect 14642 10189 14648 10192
rect 14614 10183 14648 10189
rect 14614 10180 14626 10183
rect 14292 10152 14626 10180
rect 14614 10149 14626 10152
rect 14614 10143 14648 10149
rect 14642 10140 14648 10143
rect 14700 10140 14706 10192
rect 15764 10180 15792 10211
rect 16298 10208 16304 10260
rect 16356 10208 16362 10260
rect 18049 10251 18107 10257
rect 18049 10217 18061 10251
rect 18095 10217 18107 10251
rect 18049 10211 18107 10217
rect 16209 10183 16267 10189
rect 16209 10180 16221 10183
rect 15764 10152 16221 10180
rect 16209 10149 16221 10152
rect 16255 10149 16267 10183
rect 18064 10180 18092 10211
rect 18322 10208 18328 10260
rect 18380 10208 18386 10260
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 20763 10220 21404 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 21376 10189 21404 10220
rect 18233 10183 18291 10189
rect 18233 10180 18245 10183
rect 18064 10152 18245 10180
rect 16209 10143 16267 10149
rect 18233 10149 18245 10152
rect 18279 10149 18291 10183
rect 18233 10143 18291 10149
rect 21361 10183 21419 10189
rect 21361 10149 21373 10183
rect 21407 10149 21419 10183
rect 21361 10143 21419 10149
rect 11609 10115 11667 10121
rect 11609 10081 11621 10115
rect 11655 10081 11667 10115
rect 11609 10075 11667 10081
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 11624 9908 11652 10075
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12492 10084 12817 10112
rect 12492 10072 12498 10084
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 13136 10084 13185 10112
rect 13136 10072 13142 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10081 13507 10115
rect 13998 10112 14004 10124
rect 13449 10075 13507 10081
rect 13556 10084 14004 10112
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 11808 10016 12541 10044
rect 11808 9985 11836 10016
rect 12529 10013 12541 10016
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 12710 10004 12716 10056
rect 12768 10004 12774 10056
rect 12894 10004 12900 10056
rect 12952 10004 12958 10056
rect 13464 10044 13492 10075
rect 13096 10016 13492 10044
rect 11793 9979 11851 9985
rect 11793 9945 11805 9979
rect 11839 9945 11851 9979
rect 11793 9939 11851 9945
rect 12069 9979 12127 9985
rect 12069 9945 12081 9979
rect 12115 9976 12127 9979
rect 12636 9976 12664 10004
rect 13096 9985 13124 10016
rect 13081 9979 13139 9985
rect 13081 9976 13093 9979
rect 12115 9948 12664 9976
rect 12728 9948 13093 9976
rect 12115 9945 12127 9948
rect 12069 9939 12127 9945
rect 12342 9908 12348 9920
rect 11624 9880 12348 9908
rect 12342 9868 12348 9880
rect 12400 9908 12406 9920
rect 12728 9908 12756 9948
rect 13081 9945 13093 9948
rect 13127 9945 13139 9979
rect 13081 9939 13139 9945
rect 13173 9979 13231 9985
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 13556 9976 13584 10084
rect 13998 10072 14004 10084
rect 14056 10112 14062 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 14056 10084 14105 10112
rect 14056 10072 14062 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 16758 10072 16764 10124
rect 16816 10112 16822 10124
rect 16925 10115 16983 10121
rect 16925 10112 16937 10115
rect 16816 10084 16937 10112
rect 16816 10072 16822 10084
rect 16925 10081 16937 10084
rect 16971 10081 16983 10115
rect 16925 10075 16983 10081
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19593 10115 19651 10121
rect 19593 10112 19605 10115
rect 19484 10084 19605 10112
rect 19484 10072 19490 10084
rect 19593 10081 19605 10084
rect 19639 10081 19651 10115
rect 19593 10075 19651 10081
rect 21729 10115 21787 10121
rect 21729 10081 21741 10115
rect 21775 10112 21787 10115
rect 31662 10112 31668 10124
rect 21775 10084 31668 10112
rect 21775 10081 21787 10084
rect 21729 10075 21787 10081
rect 31662 10072 31668 10084
rect 31720 10072 31726 10124
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 13688 10016 14381 10044
rect 13688 10004 13694 10016
rect 14369 10013 14381 10016
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10013 16727 10047
rect 18690 10044 18696 10056
rect 16669 10007 16727 10013
rect 18248 10016 18696 10044
rect 13219 9948 13584 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 12400 9880 12756 9908
rect 12805 9911 12863 9917
rect 12400 9868 12406 9880
rect 12805 9877 12817 9911
rect 12851 9908 12863 9911
rect 13446 9908 13452 9920
rect 12851 9880 13452 9908
rect 12851 9877 12863 9880
rect 12805 9871 12863 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 14001 9911 14059 9917
rect 14001 9877 14013 9911
rect 14047 9908 14059 9911
rect 14366 9908 14372 9920
rect 14047 9880 14372 9908
rect 14047 9877 14059 9880
rect 14001 9871 14059 9877
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 16684 9908 16712 10007
rect 18248 9920 18276 10016
rect 18690 10004 18696 10016
rect 18748 10044 18754 10056
rect 19242 10044 19248 10056
rect 18748 10016 19248 10044
rect 18748 10004 18754 10016
rect 19242 10004 19248 10016
rect 19300 10044 19306 10056
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 19300 10016 19349 10044
rect 19300 10004 19306 10016
rect 19337 10013 19349 10016
rect 19383 10013 19395 10047
rect 19337 10007 19395 10013
rect 18230 9908 18236 9920
rect 16684 9880 18236 9908
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10321 9707 10379 9713
rect 10321 9704 10333 9707
rect 10100 9676 10333 9704
rect 10100 9664 10106 9676
rect 9766 9460 9772 9512
rect 9824 9460 9830 9512
rect 10152 9509 10180 9676
rect 10321 9673 10333 9676
rect 10367 9673 10379 9707
rect 10321 9667 10379 9673
rect 11609 9707 11667 9713
rect 11609 9673 11621 9707
rect 11655 9704 11667 9707
rect 11790 9704 11796 9716
rect 11655 9676 11796 9704
rect 11655 9673 11667 9676
rect 11609 9667 11667 9673
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 11931 9676 12296 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 12268 9636 12296 9676
rect 12342 9664 12348 9716
rect 12400 9664 12406 9716
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 12713 9707 12771 9713
rect 12713 9704 12725 9707
rect 12584 9676 12725 9704
rect 12584 9664 12590 9676
rect 12713 9673 12725 9676
rect 12759 9673 12771 9707
rect 12713 9667 12771 9673
rect 12728 9636 12756 9667
rect 12894 9664 12900 9716
rect 12952 9704 12958 9716
rect 12989 9707 13047 9713
rect 12989 9704 13001 9707
rect 12952 9676 13001 9704
rect 12952 9664 12958 9676
rect 12989 9673 13001 9676
rect 13035 9673 13047 9707
rect 16025 9707 16083 9713
rect 12989 9667 13047 9673
rect 13556 9676 14320 9704
rect 11532 9608 12112 9636
rect 12268 9608 12664 9636
rect 12728 9608 13216 9636
rect 11532 9568 11560 9608
rect 12084 9580 12112 9608
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 10520 9540 11560 9568
rect 10520 9509 10548 9540
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9469 11483 9503
rect 11425 9463 11483 9469
rect 11440 9432 11468 9463
rect 9140 9404 11468 9432
rect 11532 9432 11560 9540
rect 11624 9540 11989 9568
rect 11624 9509 11652 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 12636 9577 12664 9608
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12124 9540 12449 9568
rect 12124 9528 12130 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 11609 9503 11667 9509
rect 11609 9469 11621 9503
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 11707 9503 11765 9509
rect 11707 9469 11719 9503
rect 11753 9469 11765 9503
rect 11707 9463 11765 9469
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 11931 9472 12434 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 11716 9432 11744 9463
rect 12406 9444 12434 9472
rect 12526 9460 12532 9512
rect 12584 9496 12590 9512
rect 12584 9468 12664 9496
rect 12584 9460 12590 9468
rect 11532 9404 11744 9432
rect 9140 9376 9168 9404
rect 9122 9324 9128 9376
rect 9180 9324 9186 9376
rect 11440 9364 11468 9404
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 12253 9435 12311 9441
rect 12253 9432 12265 9435
rect 11848 9404 12265 9432
rect 11848 9392 11854 9404
rect 12253 9401 12265 9404
rect 12299 9401 12311 9435
rect 12406 9404 12440 9444
rect 12253 9395 12311 9401
rect 12434 9392 12440 9404
rect 12492 9392 12498 9444
rect 12636 9432 12664 9468
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 12912 9432 12940 9463
rect 12986 9460 12992 9512
rect 13044 9460 13050 9512
rect 13188 9509 13216 9608
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9469 13231 9503
rect 13173 9463 13231 9469
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 13556 9509 13584 9676
rect 13998 9596 14004 9648
rect 14056 9596 14062 9648
rect 14292 9645 14320 9676
rect 16025 9673 16037 9707
rect 16071 9704 16083 9707
rect 16298 9704 16304 9716
rect 16071 9676 16304 9704
rect 16071 9673 16083 9676
rect 16025 9667 16083 9673
rect 16298 9664 16304 9676
rect 16356 9704 16362 9716
rect 16669 9707 16727 9713
rect 16356 9676 16528 9704
rect 16356 9664 16362 9676
rect 16500 9674 16528 9676
rect 14093 9639 14151 9645
rect 14093 9605 14105 9639
rect 14139 9605 14151 9639
rect 14093 9599 14151 9605
rect 14277 9639 14335 9645
rect 14277 9605 14289 9639
rect 14323 9605 14335 9639
rect 16209 9639 16267 9645
rect 16209 9636 16221 9639
rect 14277 9599 14335 9605
rect 15212 9608 16221 9636
rect 14108 9568 14136 9599
rect 15212 9568 15240 9608
rect 16209 9605 16221 9608
rect 16255 9636 16267 9639
rect 16390 9636 16396 9648
rect 16255 9608 16396 9636
rect 16255 9605 16267 9608
rect 16209 9599 16267 9605
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 16500 9646 16620 9674
rect 16669 9673 16681 9707
rect 16715 9704 16727 9707
rect 16758 9704 16764 9716
rect 16715 9676 16764 9704
rect 16715 9673 16727 9676
rect 16669 9667 16727 9673
rect 16758 9664 16764 9676
rect 16816 9664 16822 9716
rect 16960 9676 17172 9704
rect 16592 9636 16620 9646
rect 16960 9636 16988 9676
rect 16592 9608 16988 9636
rect 17034 9596 17040 9648
rect 17092 9596 17098 9648
rect 17144 9636 17172 9676
rect 19061 9639 19119 9645
rect 17144 9608 17816 9636
rect 14108 9540 15240 9568
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 13504 9472 13553 9500
rect 13504 9460 13510 9472
rect 13541 9469 13553 9472
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 13906 9500 13912 9512
rect 13771 9472 13912 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 13906 9460 13912 9472
rect 13964 9460 13970 9512
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9500 14151 9503
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 14139 9472 14197 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14384 9472 14596 9500
rect 13078 9432 13084 9444
rect 12636 9404 13084 9432
rect 13078 9392 13084 9404
rect 13136 9432 13142 9444
rect 13633 9435 13691 9441
rect 13136 9404 13584 9432
rect 13136 9392 13142 9404
rect 13556 9376 13584 9404
rect 13633 9401 13645 9435
rect 13679 9432 13691 9435
rect 13817 9435 13875 9441
rect 13817 9432 13829 9435
rect 13679 9404 13829 9432
rect 13679 9401 13691 9404
rect 13633 9395 13691 9401
rect 13817 9401 13829 9404
rect 13863 9401 13875 9435
rect 13817 9395 13875 9401
rect 12342 9364 12348 9376
rect 11440 9336 12348 9364
rect 12342 9324 12348 9336
rect 12400 9364 12406 9376
rect 12802 9364 12808 9376
rect 12400 9336 12808 9364
rect 12400 9324 12406 9336
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13538 9324 13544 9376
rect 13596 9364 13602 9376
rect 14108 9364 14136 9463
rect 14384 9432 14412 9472
rect 14200 9404 14412 9432
rect 14200 9373 14228 9404
rect 14458 9392 14464 9444
rect 14516 9392 14522 9444
rect 14568 9432 14596 9472
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 15212 9509 15240 9540
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 16724 9540 17356 9568
rect 16724 9528 16730 9540
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9469 15255 9503
rect 15197 9463 15255 9469
rect 15378 9460 15384 9512
rect 15436 9460 15442 9512
rect 15654 9460 15660 9512
rect 15712 9460 15718 9512
rect 15930 9500 15936 9512
rect 15856 9472 15936 9500
rect 15289 9435 15347 9441
rect 14568 9404 15240 9432
rect 13596 9336 14136 9364
rect 14185 9367 14243 9373
rect 13596 9324 13602 9336
rect 14185 9333 14197 9367
rect 14231 9333 14243 9367
rect 14185 9327 14243 9333
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14332 9336 14749 9364
rect 14332 9324 14338 9336
rect 14737 9333 14749 9336
rect 14783 9333 14795 9367
rect 15212 9364 15240 9404
rect 15289 9401 15301 9435
rect 15335 9432 15347 9435
rect 15749 9435 15807 9441
rect 15749 9432 15761 9435
rect 15335 9404 15761 9432
rect 15335 9401 15347 9404
rect 15289 9395 15347 9401
rect 15749 9401 15761 9404
rect 15795 9401 15807 9435
rect 15749 9395 15807 9401
rect 15856 9364 15884 9472
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9500 16083 9503
rect 16117 9503 16175 9509
rect 16117 9500 16129 9503
rect 16071 9472 16129 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16117 9469 16129 9472
rect 16163 9500 16175 9503
rect 16206 9500 16212 9512
rect 16163 9472 16212 9500
rect 16163 9469 16175 9472
rect 16117 9463 16175 9469
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 16408 9432 16436 9463
rect 16482 9460 16488 9512
rect 16540 9460 16546 9512
rect 17328 9509 17356 9540
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 17313 9503 17371 9509
rect 16684 9472 16988 9500
rect 16684 9432 16712 9472
rect 16408 9404 16712 9432
rect 16850 9392 16856 9444
rect 16908 9392 16914 9444
rect 16960 9432 16988 9472
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 17420 9500 17448 9528
rect 17788 9509 17816 9608
rect 19061 9605 19073 9639
rect 19107 9636 19119 9639
rect 19107 9608 19472 9636
rect 19107 9605 19119 9608
rect 19061 9599 19119 9605
rect 19444 9512 19472 9608
rect 17497 9503 17555 9509
rect 17497 9500 17509 9503
rect 17420 9472 17509 9500
rect 17313 9463 17371 9469
rect 17497 9469 17509 9472
rect 17543 9469 17555 9503
rect 17497 9463 17555 9469
rect 17773 9503 17831 9509
rect 17773 9469 17785 9503
rect 17819 9469 17831 9503
rect 17773 9463 17831 9469
rect 18877 9503 18935 9509
rect 18877 9469 18889 9503
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 16960 9404 17417 9432
rect 17405 9401 17417 9404
rect 17451 9401 17463 9435
rect 17512 9432 17540 9463
rect 18892 9432 18920 9463
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19484 9472 19533 9500
rect 19484 9460 19490 9472
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 28258 9500 28264 9512
rect 19935 9472 28264 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 28258 9460 28264 9472
rect 28316 9460 28322 9512
rect 17512 9404 18920 9432
rect 17405 9395 17463 9401
rect 20070 9392 20076 9444
rect 20128 9392 20134 9444
rect 20441 9435 20499 9441
rect 20441 9401 20453 9435
rect 20487 9432 20499 9435
rect 20487 9404 22094 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 15212 9336 15884 9364
rect 16117 9367 16175 9373
rect 14737 9327 14795 9333
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16666 9364 16672 9376
rect 16163 9336 16672 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 17954 9324 17960 9376
rect 18012 9324 18018 9376
rect 22066 9364 22094 9404
rect 28258 9364 28264 9376
rect 22066 9336 28264 9364
rect 28258 9324 28264 9336
rect 28316 9324 28322 9376
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 9309 9163 9367 9169
rect 9309 9129 9321 9163
rect 9355 9129 9367 9163
rect 9309 9123 9367 9129
rect 10781 9163 10839 9169
rect 10781 9129 10793 9163
rect 10827 9129 10839 9163
rect 12250 9160 12256 9172
rect 10781 9123 10839 9129
rect 11808 9132 12256 9160
rect 9324 9092 9352 9123
rect 9674 9101 9680 9104
rect 9646 9095 9680 9101
rect 9646 9092 9658 9095
rect 9324 9064 9658 9092
rect 9646 9061 9658 9064
rect 9646 9055 9680 9061
rect 9674 9052 9680 9055
rect 9732 9052 9738 9104
rect 10796 9092 10824 9123
rect 11057 9095 11115 9101
rect 11057 9092 11069 9095
rect 10796 9064 11069 9092
rect 11057 9061 11069 9064
rect 11103 9061 11115 9095
rect 11057 9055 11115 9061
rect 9122 8984 9128 9036
rect 9180 8984 9186 9036
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 11808 9033 11836 9132
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12342 9120 12348 9172
rect 12400 9120 12406 9172
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9129 12495 9163
rect 12437 9123 12495 9129
rect 14369 9163 14427 9169
rect 14369 9129 14381 9163
rect 14415 9160 14427 9163
rect 14458 9160 14464 9172
rect 14415 9132 14464 9160
rect 14415 9129 14427 9132
rect 14369 9123 14427 9129
rect 12066 9052 12072 9104
rect 12124 9092 12130 9104
rect 12452 9092 12480 9123
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 16206 9160 16212 9172
rect 14608 9132 16212 9160
rect 14608 9120 14614 9132
rect 16206 9120 16212 9132
rect 16264 9160 16270 9172
rect 16574 9160 16580 9172
rect 16264 9132 16580 9160
rect 16264 9120 16270 9132
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 17954 9120 17960 9172
rect 18012 9120 18018 9172
rect 19705 9163 19763 9169
rect 19705 9129 19717 9163
rect 19751 9160 19763 9163
rect 20070 9160 20076 9172
rect 19751 9132 20076 9160
rect 19751 9129 19763 9132
rect 19705 9123 19763 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 12124 9064 12480 9092
rect 12124 9052 12130 9064
rect 12526 9052 12532 9104
rect 12584 9052 12590 9104
rect 13906 9092 13912 9104
rect 12820 9064 13912 9092
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 10704 8996 11805 9024
rect 10704 8832 10732 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 11974 8984 11980 9036
rect 12032 8984 12038 9036
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 12437 9027 12495 9033
rect 12437 9024 12449 9027
rect 12391 8996 12449 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12437 8993 12449 8996
rect 12483 9024 12495 9027
rect 12544 9024 12572 9052
rect 12483 8996 12572 9024
rect 12483 8993 12495 8996
rect 12437 8987 12495 8993
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 12820 9033 12848 9064
rect 13906 9052 13912 9064
rect 13964 9092 13970 9104
rect 15378 9092 15384 9104
rect 13964 9064 15384 9092
rect 13964 9052 13970 9064
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 15841 9095 15899 9101
rect 15841 9061 15853 9095
rect 15887 9092 15899 9095
rect 16485 9095 16543 9101
rect 16485 9092 16497 9095
rect 15887 9064 16497 9092
rect 15887 9061 15899 9064
rect 15841 9055 15899 9061
rect 16485 9061 16497 9064
rect 16531 9061 16543 9095
rect 16485 9055 16543 9061
rect 16684 9092 16712 9120
rect 17865 9095 17923 9101
rect 16684 9064 17356 9092
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12676 8996 12817 9024
rect 12676 8984 12682 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 11931 8928 12081 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12713 8959 12771 8965
rect 12069 8919 12127 8925
rect 12268 8928 12664 8956
rect 12268 8897 12296 8928
rect 12253 8891 12311 8897
rect 12253 8888 12265 8891
rect 11808 8860 12265 8888
rect 11808 8832 11836 8860
rect 12253 8857 12265 8860
rect 12299 8857 12311 8891
rect 12253 8851 12311 8857
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 12526 8888 12532 8900
rect 12400 8860 12532 8888
rect 12400 8848 12406 8860
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 12636 8888 12664 8928
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 12897 8959 12955 8965
rect 12897 8956 12909 8959
rect 12759 8928 12909 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 12897 8925 12909 8928
rect 12943 8925 12955 8959
rect 13004 8956 13032 8987
rect 13078 8984 13084 9036
rect 13136 8984 13142 9036
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 14056 8996 14289 9024
rect 14056 8984 14062 8996
rect 14277 8993 14289 8996
rect 14323 8993 14335 9027
rect 14277 8987 14335 8993
rect 14366 8984 14372 9036
rect 14424 9024 14430 9036
rect 14461 9027 14519 9033
rect 14461 9024 14473 9027
rect 14424 8996 14473 9024
rect 14424 8984 14430 8996
rect 14461 8993 14473 8996
rect 14507 8993 14519 9027
rect 15396 9024 15424 9052
rect 15749 9027 15807 9033
rect 15749 9024 15761 9027
rect 15396 8996 15761 9024
rect 14461 8987 14519 8993
rect 15749 8993 15761 8996
rect 15795 8993 15807 9027
rect 15749 8987 15807 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 15948 8956 15976 8987
rect 16114 8984 16120 9036
rect 16172 8984 16178 9036
rect 16209 9027 16267 9033
rect 16209 8993 16221 9027
rect 16255 9024 16267 9027
rect 16298 9024 16304 9036
rect 16255 8996 16304 9024
rect 16255 8993 16267 8996
rect 16209 8987 16267 8993
rect 16224 8956 16252 8987
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 16684 9033 16712 9064
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 16758 8984 16764 9036
rect 16816 8984 16822 9036
rect 17328 9033 17356 9064
rect 17865 9061 17877 9095
rect 17911 9092 17923 9095
rect 17972 9092 18000 9120
rect 18570 9095 18628 9101
rect 18570 9092 18582 9095
rect 17911 9064 18582 9092
rect 17911 9061 17923 9064
rect 17865 9055 17923 9061
rect 18570 9061 18582 9064
rect 18616 9061 18628 9095
rect 18570 9055 18628 9061
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 17129 9027 17187 9033
rect 17129 9024 17141 9027
rect 17083 8996 17141 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 17129 8993 17141 8996
rect 17175 8993 17187 9027
rect 17129 8987 17187 8993
rect 17313 9027 17371 9033
rect 17313 8993 17325 9027
rect 17359 9024 17371 9027
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 17359 8996 17417 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 17405 8987 17463 8993
rect 21358 8984 21364 9036
rect 21416 8984 21422 9036
rect 13004 8928 13216 8956
rect 15948 8928 16252 8956
rect 16393 8959 16451 8965
rect 12897 8919 12955 8925
rect 13188 8900 13216 8928
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 16439 8928 17233 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18288 8928 18337 8956
rect 18288 8916 18294 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 13170 8888 13176 8900
rect 12636 8860 13176 8888
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 14642 8848 14648 8900
rect 14700 8888 14706 8900
rect 16761 8891 16819 8897
rect 16761 8888 16773 8891
rect 14700 8860 16773 8888
rect 14700 8848 14706 8860
rect 16761 8857 16773 8860
rect 16807 8888 16819 8891
rect 16807 8860 17724 8888
rect 16807 8857 16819 8860
rect 16761 8851 16819 8857
rect 17696 8832 17724 8860
rect 10686 8780 10692 8832
rect 10744 8780 10750 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 11790 8780 11796 8832
rect 11848 8780 11854 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 15013 8823 15071 8829
rect 15013 8789 15025 8823
rect 15059 8820 15071 8823
rect 15286 8820 15292 8832
rect 15059 8792 15292 8820
rect 15059 8789 15071 8792
rect 15013 8783 15071 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 16298 8780 16304 8832
rect 16356 8780 16362 8832
rect 17586 8780 17592 8832
rect 17644 8780 17650 8832
rect 17678 8780 17684 8832
rect 17736 8780 17742 8832
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18690 8820 18696 8832
rect 18187 8792 18696 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 21637 8823 21695 8829
rect 21637 8789 21649 8823
rect 21683 8820 21695 8823
rect 31662 8820 31668 8832
rect 21683 8792 31668 8820
rect 21683 8789 21695 8792
rect 21637 8783 21695 8789
rect 31662 8780 31668 8792
rect 31720 8780 31726 8832
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9456 8588 9597 8616
rect 9456 8576 9462 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 9674 8576 9680 8628
rect 9732 8576 9738 8628
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12584 8588 13093 8616
rect 12584 8576 12590 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13228 8588 13553 8616
rect 13228 8576 13234 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 13909 8619 13967 8625
rect 13909 8616 13921 8619
rect 13872 8588 13921 8616
rect 13872 8576 13878 8588
rect 13909 8585 13921 8588
rect 13955 8585 13967 8619
rect 15013 8619 15071 8625
rect 15013 8616 15025 8619
rect 13909 8579 13967 8585
rect 14844 8588 15025 8616
rect 9692 8480 9720 8576
rect 14844 8548 14872 8588
rect 15013 8585 15025 8588
rect 15059 8585 15071 8619
rect 15013 8579 15071 8585
rect 16298 8576 16304 8628
rect 16356 8576 16362 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 19334 8616 19340 8628
rect 16448 8588 19340 8616
rect 16448 8576 16454 8588
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 20809 8619 20867 8625
rect 20809 8585 20821 8619
rect 20855 8616 20867 8619
rect 21358 8616 21364 8628
rect 20855 8588 21364 8616
rect 20855 8585 20867 8588
rect 20809 8579 20867 8585
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 13740 8520 14872 8548
rect 15105 8551 15163 8557
rect 13173 8483 13231 8489
rect 9692 8452 10088 8480
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 9950 8412 9956 8424
rect 9815 8384 9956 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10060 8421 10088 8452
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13740 8480 13768 8520
rect 13219 8452 13768 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 14108 8424 14136 8520
rect 15105 8517 15117 8551
rect 15151 8548 15163 8551
rect 15151 8520 15516 8548
rect 15151 8517 15163 8520
rect 15105 8511 15163 8517
rect 14642 8480 14648 8492
rect 14384 8452 14648 8480
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8381 10103 8415
rect 10045 8375 10103 8381
rect 10686 8372 10692 8424
rect 10744 8372 10750 8424
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 11848 8384 11897 8412
rect 11848 8372 11854 8384
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 11885 8375 11943 8381
rect 13081 8415 13139 8421
rect 13081 8381 13093 8415
rect 13127 8412 13139 8415
rect 13538 8412 13544 8424
rect 13127 8384 13544 8412
rect 13127 8381 13139 8384
rect 13081 8375 13139 8381
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8381 13691 8415
rect 13633 8375 13691 8381
rect 10410 8304 10416 8356
rect 10468 8304 10474 8356
rect 13354 8304 13360 8356
rect 13412 8304 13418 8356
rect 10502 8236 10508 8288
rect 10560 8236 10566 8288
rect 11698 8236 11704 8288
rect 11756 8236 11762 8288
rect 13648 8276 13676 8375
rect 13906 8372 13912 8424
rect 13964 8421 13970 8424
rect 13964 8412 13973 8421
rect 13964 8406 14009 8412
rect 13964 8378 14044 8406
rect 13964 8375 13973 8378
rect 13964 8372 13970 8375
rect 14016 8344 14044 8378
rect 14090 8372 14096 8424
rect 14148 8372 14154 8424
rect 14384 8422 14412 8452
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14384 8421 14504 8422
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14384 8415 14519 8421
rect 14384 8394 14473 8415
rect 14277 8375 14335 8381
rect 14461 8381 14473 8394
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 14292 8344 14320 8375
rect 14550 8372 14556 8424
rect 14608 8372 14614 8424
rect 14826 8372 14832 8424
rect 14884 8372 14890 8424
rect 15194 8372 15200 8424
rect 15252 8372 15258 8424
rect 15286 8372 15292 8424
rect 15344 8372 15350 8424
rect 15488 8421 15516 8520
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 16316 8412 16344 8576
rect 17586 8508 17592 8560
rect 17644 8508 17650 8560
rect 18230 8508 18236 8560
rect 18288 8548 18294 8560
rect 18288 8520 19472 8548
rect 18288 8508 18294 8520
rect 16393 8415 16451 8421
rect 16393 8412 16405 8415
rect 15519 8384 16405 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 16393 8381 16405 8384
rect 16439 8381 16451 8415
rect 17604 8412 17632 8508
rect 17678 8440 17684 8492
rect 17736 8480 17742 8492
rect 19444 8489 19472 8520
rect 19429 8483 19487 8489
rect 17736 8452 18736 8480
rect 17736 8440 17742 8452
rect 18708 8421 18736 8452
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 18325 8415 18383 8421
rect 18325 8412 18337 8415
rect 17604 8384 18337 8412
rect 16393 8375 16451 8381
rect 18325 8381 18337 8384
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 14016 8316 14320 8344
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14921 8347 14979 8353
rect 14921 8344 14933 8347
rect 14415 8316 14933 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14921 8313 14933 8316
rect 14967 8313 14979 8347
rect 14921 8307 14979 8313
rect 17402 8304 17408 8356
rect 17460 8344 17466 8356
rect 17957 8347 18015 8353
rect 17957 8344 17969 8347
rect 17460 8316 17969 8344
rect 17460 8304 17466 8316
rect 17957 8313 17969 8316
rect 18003 8313 18015 8347
rect 18340 8344 18368 8375
rect 19674 8347 19732 8353
rect 19674 8344 19686 8347
rect 18340 8316 19686 8344
rect 17957 8307 18015 8313
rect 19674 8313 19686 8316
rect 19720 8313 19732 8347
rect 19674 8307 19732 8313
rect 14550 8276 14556 8288
rect 13648 8248 14556 8276
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 15381 8279 15439 8285
rect 15381 8276 15393 8279
rect 14884 8248 15393 8276
rect 14884 8236 14890 8248
rect 15381 8245 15393 8248
rect 15427 8245 15439 8279
rect 15381 8239 15439 8245
rect 16574 8236 16580 8288
rect 16632 8236 16638 8288
rect 18874 8236 18880 8288
rect 18932 8236 18938 8288
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 12621 8075 12679 8081
rect 10008 8044 12572 8072
rect 10008 8032 10014 8044
rect 9668 8007 9726 8013
rect 9668 7973 9680 8007
rect 9714 8004 9726 8007
rect 10042 8004 10048 8016
rect 9714 7976 10048 8004
rect 9714 7973 9726 7976
rect 9668 7967 9726 7973
rect 10042 7964 10048 7976
rect 10100 8004 10106 8016
rect 10502 8004 10508 8016
rect 10100 7976 10508 8004
rect 10100 7964 10106 7976
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 11508 8007 11566 8013
rect 11508 7973 11520 8007
rect 11554 8004 11566 8007
rect 11698 8004 11704 8016
rect 11554 7976 11704 8004
rect 11554 7973 11566 7976
rect 11508 7967 11566 7973
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 9456 7908 11253 7936
rect 9456 7896 9462 7908
rect 11241 7905 11253 7908
rect 11287 7936 11299 7939
rect 11287 7908 12434 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 12406 7800 12434 7908
rect 12544 7868 12572 8044
rect 12621 8041 12633 8075
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 12636 8004 12664 8035
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 13412 8044 13461 8072
rect 13412 8032 13418 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 14550 8032 14556 8084
rect 14608 8032 14614 8084
rect 14921 8075 14979 8081
rect 14921 8041 14933 8075
rect 14967 8041 14979 8075
rect 14921 8035 14979 8041
rect 18141 8075 18199 8081
rect 18141 8041 18153 8075
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 20165 8075 20223 8081
rect 20165 8041 20177 8075
rect 20211 8072 20223 8075
rect 20211 8044 20392 8072
rect 20211 8041 20223 8044
rect 20165 8035 20223 8041
rect 12805 8007 12863 8013
rect 12805 8004 12817 8007
rect 12636 7976 12817 8004
rect 12805 7973 12817 7976
rect 12851 7973 12863 8007
rect 14568 8004 14596 8032
rect 12805 7967 12863 7973
rect 13556 7976 14596 8004
rect 14936 8004 14964 8035
rect 15197 8007 15255 8013
rect 15197 8004 15209 8007
rect 14936 7976 15209 8004
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7936 13415 7939
rect 13446 7936 13452 7948
rect 13403 7908 13452 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13556 7945 13584 7976
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7905 13599 7939
rect 13541 7899 13599 7905
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 14090 7936 14096 7948
rect 13679 7908 14096 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14568 7936 14596 7976
rect 15197 7973 15209 7976
rect 15243 8004 15255 8007
rect 15286 8004 15292 8016
rect 15243 7976 15292 8004
rect 15243 7973 15255 7976
rect 15197 7967 15255 7973
rect 15286 7964 15292 7976
rect 15344 7964 15350 8016
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 17006 8007 17064 8013
rect 17006 8004 17018 8007
rect 16632 7976 17018 8004
rect 16632 7964 16638 7976
rect 17006 7973 17018 7976
rect 17052 7973 17064 8007
rect 18156 8004 18184 8035
rect 18325 8007 18383 8013
rect 18325 8004 18337 8007
rect 18156 7976 18337 8004
rect 17006 7967 17064 7973
rect 18325 7973 18337 7976
rect 18371 7973 18383 8007
rect 18325 7967 18383 7973
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 20364 8013 20392 8044
rect 19030 8007 19088 8013
rect 19030 8004 19042 8007
rect 18932 7976 19042 8004
rect 18932 7964 18938 7976
rect 19030 7973 19042 7976
rect 19076 7973 19088 8007
rect 19030 7967 19088 7973
rect 20349 8007 20407 8013
rect 20349 7973 20361 8007
rect 20395 7973 20407 8007
rect 20349 7967 20407 7973
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 14568 7908 14749 7936
rect 14737 7905 14749 7908
rect 14783 7905 14795 7939
rect 14737 7899 14795 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7936 15715 7939
rect 16390 7936 16396 7948
rect 15703 7908 16396 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 15672 7868 15700 7899
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 18230 7936 18236 7948
rect 16776 7908 18236 7936
rect 16776 7877 16804 7908
rect 18230 7896 18236 7908
rect 18288 7936 18294 7948
rect 18785 7939 18843 7945
rect 18785 7936 18797 7939
rect 18288 7908 18797 7936
rect 18288 7896 18294 7908
rect 18785 7905 18797 7908
rect 18831 7905 18843 7939
rect 18785 7899 18843 7905
rect 16761 7871 16819 7877
rect 16761 7868 16773 7871
rect 12544 7840 15700 7868
rect 15856 7840 16773 7868
rect 13630 7800 13636 7812
rect 12406 7772 13636 7800
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 15856 7809 15884 7840
rect 16761 7837 16773 7840
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 15841 7803 15899 7809
rect 15841 7800 15853 7803
rect 15028 7772 15853 7800
rect 15028 7744 15056 7772
rect 15841 7769 15853 7772
rect 15887 7769 15899 7803
rect 15841 7763 15899 7769
rect 10778 7692 10784 7744
rect 10836 7692 10842 7744
rect 12894 7692 12900 7744
rect 12952 7692 12958 7744
rect 13814 7692 13820 7744
rect 13872 7692 13878 7744
rect 15010 7692 15016 7744
rect 15068 7692 15074 7744
rect 15470 7692 15476 7744
rect 15528 7692 15534 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 18417 7735 18475 7741
rect 18417 7732 18429 7735
rect 18104 7704 18429 7732
rect 18104 7692 18110 7704
rect 18417 7701 18429 7704
rect 18463 7701 18475 7735
rect 18417 7695 18475 7701
rect 20622 7692 20628 7744
rect 20680 7692 20686 7744
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 9766 7488 9772 7540
rect 9824 7488 9830 7540
rect 10778 7488 10784 7540
rect 10836 7488 10842 7540
rect 10042 7284 10048 7336
rect 10100 7284 10106 7336
rect 10796 7333 10824 7488
rect 15010 7352 15016 7404
rect 15068 7352 15074 7404
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 11698 7284 11704 7336
rect 11756 7284 11762 7336
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7324 13599 7327
rect 13630 7324 13636 7336
rect 13587 7296 13636 7324
rect 13587 7293 13599 7296
rect 13541 7287 13599 7293
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13814 7333 13820 7336
rect 13808 7324 13820 7333
rect 13775 7296 13820 7324
rect 13808 7287 13820 7296
rect 13814 7284 13820 7287
rect 13872 7284 13878 7336
rect 15286 7333 15292 7336
rect 15280 7324 15292 7333
rect 15247 7296 15292 7324
rect 15280 7287 15292 7296
rect 15286 7284 15292 7287
rect 15344 7284 15350 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 16945 7327 17003 7333
rect 16945 7324 16957 7327
rect 16632 7296 16957 7324
rect 16632 7284 16638 7296
rect 16945 7293 16957 7296
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18932 7296 18981 7324
rect 18932 7284 18938 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 19334 7216 19340 7268
rect 19392 7216 19398 7268
rect 10870 7148 10876 7200
rect 10928 7148 10934 7200
rect 11790 7148 11796 7200
rect 11848 7148 11854 7200
rect 14918 7148 14924 7200
rect 14976 7148 14982 7200
rect 16393 7191 16451 7197
rect 16393 7157 16405 7191
rect 16439 7188 16451 7191
rect 16574 7188 16580 7200
rect 16439 7160 16580 7188
rect 16439 7157 16451 7160
rect 16393 7151 16451 7157
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 17037 7191 17095 7197
rect 17037 7188 17049 7191
rect 16816 7160 17049 7188
rect 16816 7148 16822 7160
rect 17037 7157 17049 7160
rect 17083 7157 17095 7191
rect 17037 7151 17095 7157
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 13814 6876 13820 6928
rect 13872 6876 13878 6928
rect 14918 6876 14924 6928
rect 14976 6876 14982 6928
rect 16574 6876 16580 6928
rect 16632 6876 16638 6928
rect 13538 6604 13544 6656
rect 13596 6644 13602 6656
rect 13909 6647 13967 6653
rect 13909 6644 13921 6647
rect 13596 6616 13921 6644
rect 13596 6604 13602 6616
rect 13909 6613 13921 6616
rect 13955 6613 13967 6647
rect 13909 6607 13967 6613
rect 15010 6604 15016 6656
rect 15068 6604 15074 6656
rect 16298 6604 16304 6656
rect 16356 6644 16362 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 16356 6616 16681 6644
rect 16356 6604 16362 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 12618 892 12624 944
rect 12676 892 12682 944
rect 9950 824 9956 876
rect 10008 864 10014 876
rect 10045 867 10103 873
rect 10045 864 10057 867
rect 10008 836 10057 864
rect 10008 824 10014 836
rect 10045 833 10057 836
rect 10091 833 10103 867
rect 10045 827 10103 833
rect 9766 756 9772 808
rect 9824 756 9830 808
rect 12250 688 12256 740
rect 12308 728 12314 740
rect 12437 731 12495 737
rect 12437 728 12449 731
rect 12308 700 12449 728
rect 12308 688 12314 700
rect 12437 697 12449 700
rect 12483 697 12495 731
rect 12437 691 12495 697
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
rect 16022 416 16028 468
rect 16080 456 16086 468
rect 16298 456 16304 468
rect 16080 428 16304 456
rect 16080 416 16086 428
rect 16298 416 16304 428
rect 16356 416 16362 468
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 12440 12359 12492 12368
rect 12440 12325 12449 12359
rect 12449 12325 12483 12359
rect 12483 12325 12492 12359
rect 14924 12427 14976 12436
rect 14924 12393 14933 12427
rect 14933 12393 14967 12427
rect 14967 12393 14976 12427
rect 14924 12384 14976 12393
rect 12440 12316 12492 12325
rect 13360 12248 13412 12300
rect 15476 12316 15528 12368
rect 16856 12316 16908 12368
rect 20628 12384 20680 12436
rect 18972 12291 19024 12300
rect 18972 12257 18995 12291
rect 18995 12257 19024 12291
rect 18972 12248 19024 12257
rect 12716 12180 12768 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 12624 12044 12676 12096
rect 19064 12044 19116 12096
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 12440 11840 12492 11892
rect 13544 11840 13596 11892
rect 16856 11840 16908 11892
rect 18236 11840 18288 11892
rect 18788 11883 18840 11892
rect 18788 11849 18797 11883
rect 18797 11849 18831 11883
rect 18831 11849 18840 11883
rect 18788 11840 18840 11849
rect 18972 11840 19024 11892
rect 11336 11500 11388 11552
rect 12624 11636 12676 11688
rect 13360 11636 13412 11688
rect 13728 11636 13780 11688
rect 16120 11704 16172 11756
rect 16580 11679 16632 11688
rect 16580 11645 16589 11679
rect 16589 11645 16623 11679
rect 16623 11645 16632 11679
rect 16580 11636 16632 11645
rect 14924 11611 14976 11620
rect 14924 11577 14933 11611
rect 14933 11577 14967 11611
rect 14967 11577 14976 11611
rect 14924 11568 14976 11577
rect 15660 11568 15712 11620
rect 17132 11611 17184 11620
rect 17132 11577 17141 11611
rect 17141 11577 17175 11611
rect 17175 11577 17184 11611
rect 17132 11568 17184 11577
rect 18144 11636 18196 11688
rect 19248 11636 19300 11688
rect 19616 11568 19668 11620
rect 17592 11543 17644 11552
rect 17592 11509 17601 11543
rect 17601 11509 17635 11543
rect 17635 11509 17644 11543
rect 17592 11500 17644 11509
rect 18788 11500 18840 11552
rect 28264 11568 28316 11620
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 11336 11228 11388 11280
rect 14280 11339 14332 11348
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 14924 11296 14976 11348
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 17592 11296 17644 11348
rect 19340 11296 19392 11348
rect 11244 11203 11296 11212
rect 11244 11169 11278 11203
rect 11278 11169 11296 11203
rect 11244 11160 11296 11169
rect 12716 11160 12768 11212
rect 13176 11160 13228 11212
rect 17684 11228 17736 11280
rect 19616 11271 19668 11280
rect 19616 11237 19625 11271
rect 19625 11237 19659 11271
rect 19659 11237 19668 11271
rect 19616 11228 19668 11237
rect 16580 11160 16632 11212
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 16580 11024 16632 11076
rect 19340 11160 19392 11212
rect 9588 10956 9640 11008
rect 12348 10999 12400 11008
rect 12348 10965 12357 10999
rect 12357 10965 12391 10999
rect 12391 10965 12400 10999
rect 12348 10956 12400 10965
rect 16764 10999 16816 11008
rect 16764 10965 16773 10999
rect 16773 10965 16807 10999
rect 16807 10965 16816 10999
rect 16764 10956 16816 10965
rect 16856 10956 16908 11008
rect 18788 10956 18840 11008
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 11244 10752 11296 10804
rect 11428 10752 11480 10804
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 14556 10616 14608 10668
rect 16212 10752 16264 10804
rect 19984 10752 20036 10804
rect 16856 10616 16908 10668
rect 12348 10548 12400 10600
rect 12440 10548 12492 10600
rect 12532 10548 12584 10600
rect 12624 10548 12676 10600
rect 13176 10591 13228 10600
rect 13176 10557 13185 10591
rect 13185 10557 13219 10591
rect 13219 10557 13228 10591
rect 13176 10548 13228 10557
rect 13452 10480 13504 10532
rect 12440 10412 12492 10464
rect 12992 10412 13044 10464
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 18788 10548 18840 10600
rect 16764 10480 16816 10532
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 9588 10140 9640 10192
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 9404 10115 9456 10124
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 10048 10072 10100 10124
rect 12992 10140 13044 10192
rect 13176 10208 13228 10260
rect 14648 10183 14700 10192
rect 14648 10149 14660 10183
rect 14660 10149 14700 10183
rect 14648 10140 14700 10149
rect 16304 10251 16356 10260
rect 16304 10217 16313 10251
rect 16313 10217 16347 10251
rect 16347 10217 16356 10251
rect 16304 10208 16356 10217
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 12440 10115 12492 10124
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 13084 10072 13136 10124
rect 12624 10004 12676 10056
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 12348 9868 12400 9920
rect 14004 10072 14056 10124
rect 16764 10072 16816 10124
rect 19432 10072 19484 10124
rect 31668 10072 31720 10124
rect 13636 10004 13688 10056
rect 13452 9868 13504 9920
rect 14372 9868 14424 9920
rect 18696 10004 18748 10056
rect 19248 10004 19300 10056
rect 18236 9868 18288 9920
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 10048 9664 10100 9716
rect 9772 9503 9824 9512
rect 9772 9469 9781 9503
rect 9781 9469 9815 9503
rect 9815 9469 9824 9503
rect 9772 9460 9824 9469
rect 11796 9664 11848 9716
rect 12348 9707 12400 9716
rect 12348 9673 12357 9707
rect 12357 9673 12391 9707
rect 12391 9673 12400 9707
rect 12348 9664 12400 9673
rect 12532 9664 12584 9716
rect 12900 9664 12952 9716
rect 12072 9528 12124 9580
rect 12532 9503 12584 9512
rect 12532 9469 12541 9503
rect 12541 9469 12575 9503
rect 12575 9469 12584 9503
rect 12532 9460 12584 9469
rect 9128 9324 9180 9376
rect 11796 9392 11848 9444
rect 12440 9392 12492 9444
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 13452 9460 13504 9512
rect 14004 9639 14056 9648
rect 14004 9605 14013 9639
rect 14013 9605 14047 9639
rect 14047 9605 14056 9639
rect 14004 9596 14056 9605
rect 16304 9664 16356 9716
rect 16396 9596 16448 9648
rect 16764 9664 16816 9716
rect 17040 9639 17092 9648
rect 17040 9605 17049 9639
rect 17049 9605 17083 9639
rect 17083 9605 17092 9639
rect 17040 9596 17092 9605
rect 13912 9460 13964 9512
rect 13084 9392 13136 9444
rect 12348 9324 12400 9376
rect 12808 9324 12860 9376
rect 13544 9324 13596 9376
rect 14464 9435 14516 9444
rect 14464 9401 14473 9435
rect 14473 9401 14507 9435
rect 14507 9401 14516 9435
rect 14464 9392 14516 9401
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 16672 9528 16724 9580
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 15660 9503 15712 9512
rect 15660 9469 15669 9503
rect 15669 9469 15703 9503
rect 15703 9469 15712 9503
rect 15660 9460 15712 9469
rect 15936 9503 15988 9512
rect 14280 9324 14332 9376
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 16212 9460 16264 9512
rect 16488 9503 16540 9512
rect 16488 9469 16497 9503
rect 16497 9469 16531 9503
rect 16531 9469 16540 9503
rect 16488 9460 16540 9469
rect 17408 9528 17460 9580
rect 16856 9435 16908 9444
rect 16856 9401 16865 9435
rect 16865 9401 16899 9435
rect 16899 9401 16908 9435
rect 16856 9392 16908 9401
rect 19432 9460 19484 9512
rect 28264 9460 28316 9512
rect 20076 9435 20128 9444
rect 20076 9401 20085 9435
rect 20085 9401 20119 9435
rect 20119 9401 20128 9435
rect 20076 9392 20128 9401
rect 16672 9324 16724 9376
rect 17960 9367 18012 9376
rect 17960 9333 17969 9367
rect 17969 9333 18003 9367
rect 18003 9333 18012 9367
rect 17960 9324 18012 9333
rect 28264 9324 28316 9376
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 9680 9095 9732 9104
rect 9680 9061 9692 9095
rect 9692 9061 9732 9095
rect 9680 9052 9732 9061
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 12256 9120 12308 9172
rect 12348 9163 12400 9172
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 12072 9052 12124 9104
rect 14464 9120 14516 9172
rect 14556 9120 14608 9172
rect 16212 9120 16264 9172
rect 16580 9120 16632 9172
rect 16672 9120 16724 9172
rect 17960 9120 18012 9172
rect 20076 9120 20128 9172
rect 12532 9052 12584 9104
rect 11980 9027 12032 9036
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 12624 8984 12676 9036
rect 13912 9052 13964 9104
rect 15384 9052 15436 9104
rect 12348 8848 12400 8900
rect 12532 8891 12584 8900
rect 12532 8857 12541 8891
rect 12541 8857 12575 8891
rect 12575 8857 12584 8891
rect 12532 8848 12584 8857
rect 13084 9027 13136 9036
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 14004 8984 14056 9036
rect 14372 8984 14424 9036
rect 16120 9027 16172 9036
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 16304 8984 16356 9036
rect 16764 9027 16816 9036
rect 16764 8993 16773 9027
rect 16773 8993 16807 9027
rect 16807 8993 16816 9027
rect 16764 8984 16816 8993
rect 21364 9027 21416 9036
rect 21364 8993 21373 9027
rect 21373 8993 21407 9027
rect 21407 8993 21416 9027
rect 21364 8984 21416 8993
rect 18236 8916 18288 8968
rect 13176 8848 13228 8900
rect 14648 8848 14700 8900
rect 10692 8780 10744 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 11796 8780 11848 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 15292 8780 15344 8832
rect 16304 8823 16356 8832
rect 16304 8789 16313 8823
rect 16313 8789 16347 8823
rect 16347 8789 16356 8823
rect 16304 8780 16356 8789
rect 17592 8823 17644 8832
rect 17592 8789 17601 8823
rect 17601 8789 17635 8823
rect 17635 8789 17644 8823
rect 17592 8780 17644 8789
rect 17684 8780 17736 8832
rect 18696 8780 18748 8832
rect 31668 8780 31720 8832
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 9404 8576 9456 8628
rect 9680 8576 9732 8628
rect 12532 8576 12584 8628
rect 13176 8576 13228 8628
rect 13820 8576 13872 8628
rect 16304 8576 16356 8628
rect 16396 8576 16448 8628
rect 19340 8576 19392 8628
rect 21364 8576 21416 8628
rect 9956 8372 10008 8424
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 14648 8483 14700 8492
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 11796 8372 11848 8424
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 10416 8347 10468 8356
rect 10416 8313 10425 8347
rect 10425 8313 10459 8347
rect 10459 8313 10468 8347
rect 10416 8304 10468 8313
rect 13360 8347 13412 8356
rect 13360 8313 13369 8347
rect 13369 8313 13403 8347
rect 13403 8313 13412 8347
rect 13360 8304 13412 8313
rect 10508 8279 10560 8288
rect 10508 8245 10517 8279
rect 10517 8245 10551 8279
rect 10551 8245 10560 8279
rect 10508 8236 10560 8245
rect 11704 8279 11756 8288
rect 11704 8245 11713 8279
rect 11713 8245 11747 8279
rect 11747 8245 11756 8279
rect 11704 8236 11756 8245
rect 13912 8415 13964 8424
rect 13912 8381 13927 8415
rect 13927 8381 13961 8415
rect 13961 8381 13964 8415
rect 13912 8372 13964 8381
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14556 8415 14608 8424
rect 14556 8381 14565 8415
rect 14565 8381 14599 8415
rect 14599 8381 14608 8415
rect 14556 8372 14608 8381
rect 14832 8415 14884 8424
rect 14832 8381 14841 8415
rect 14841 8381 14875 8415
rect 14875 8381 14884 8415
rect 14832 8372 14884 8381
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 17592 8508 17644 8560
rect 18236 8508 18288 8560
rect 17684 8440 17736 8492
rect 17408 8304 17460 8356
rect 14556 8279 14608 8288
rect 14556 8245 14565 8279
rect 14565 8245 14599 8279
rect 14599 8245 14608 8279
rect 14556 8236 14608 8245
rect 14832 8236 14884 8288
rect 16580 8279 16632 8288
rect 16580 8245 16589 8279
rect 16589 8245 16623 8279
rect 16623 8245 16632 8279
rect 16580 8236 16632 8245
rect 18880 8279 18932 8288
rect 18880 8245 18889 8279
rect 18889 8245 18923 8279
rect 18923 8245 18932 8279
rect 18880 8236 18932 8245
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 9956 8032 10008 8084
rect 10048 7964 10100 8016
rect 10508 7964 10560 8016
rect 11704 7964 11756 8016
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 13360 8032 13412 8084
rect 14556 8032 14608 8084
rect 13452 7896 13504 7948
rect 14096 7896 14148 7948
rect 15292 7964 15344 8016
rect 16580 7964 16632 8016
rect 18880 7964 18932 8016
rect 16396 7896 16448 7948
rect 18236 7896 18288 7948
rect 13636 7760 13688 7812
rect 10784 7735 10836 7744
rect 10784 7701 10793 7735
rect 10793 7701 10827 7735
rect 10827 7701 10836 7735
rect 10784 7692 10836 7701
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 15016 7692 15068 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 18052 7692 18104 7744
rect 20628 7735 20680 7744
rect 20628 7701 20637 7735
rect 20637 7701 20671 7735
rect 20671 7701 20680 7735
rect 20628 7692 20680 7701
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10784 7488 10836 7540
rect 10048 7327 10100 7336
rect 10048 7293 10057 7327
rect 10057 7293 10091 7327
rect 10091 7293 10100 7327
rect 10048 7284 10100 7293
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 13636 7284 13688 7336
rect 13820 7327 13872 7336
rect 13820 7293 13854 7327
rect 13854 7293 13872 7327
rect 13820 7284 13872 7293
rect 15292 7327 15344 7336
rect 15292 7293 15326 7327
rect 15326 7293 15344 7327
rect 15292 7284 15344 7293
rect 16580 7284 16632 7336
rect 18880 7284 18932 7336
rect 19340 7259 19392 7268
rect 19340 7225 19349 7259
rect 19349 7225 19383 7259
rect 19383 7225 19392 7259
rect 19340 7216 19392 7225
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 16580 7148 16632 7200
rect 16764 7148 16816 7200
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 13820 6919 13872 6928
rect 13820 6885 13829 6919
rect 13829 6885 13863 6919
rect 13863 6885 13872 6919
rect 13820 6876 13872 6885
rect 14924 6919 14976 6928
rect 14924 6885 14933 6919
rect 14933 6885 14967 6919
rect 14967 6885 14976 6919
rect 14924 6876 14976 6885
rect 16580 6919 16632 6928
rect 16580 6885 16589 6919
rect 16589 6885 16623 6919
rect 16623 6885 16632 6919
rect 16580 6876 16632 6885
rect 13544 6604 13596 6656
rect 15016 6647 15068 6656
rect 15016 6613 15025 6647
rect 15025 6613 15059 6647
rect 15059 6613 15068 6647
rect 15016 6604 15068 6613
rect 16304 6604 16356 6656
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 12624 935 12676 944
rect 12624 901 12633 935
rect 12633 901 12667 935
rect 12667 901 12676 935
rect 12624 892 12676 901
rect 9956 824 10008 876
rect 9772 799 9824 808
rect 9772 765 9781 799
rect 9781 765 9815 799
rect 9815 765 9824 799
rect 9772 756 9824 765
rect 12256 688 12308 740
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
rect 16028 416 16080 468
rect 16304 416 16356 468
<< metal2 >>
rect 12898 19600 12954 20000
rect 13542 19600 13598 20000
rect 14186 19600 14242 20000
rect 14830 19600 14886 20000
rect 15474 19600 15530 20000
rect 16118 19600 16174 20000
rect 16762 19600 16818 20000
rect 16868 19638 17080 19666
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 4250 18459 4558 18468
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 4250 15260 4558 15269
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 12452 11898 12480 12310
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12636 11694 12664 12038
rect 12624 11688 12676 11694
rect 11426 11656 11482 11665
rect 12624 11630 12676 11636
rect 11426 11591 11482 11600
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 11348 11286 11376 11494
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 8102 10299 8410 10308
rect 9600 10198 9628 10950
rect 10874 10840 10930 10849
rect 11256 10810 11284 11154
rect 11440 10810 11468 11591
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11955 10843 12263 10852
rect 10874 10775 10876 10784
rect 10928 10775 10930 10784
rect 11244 10804 11296 10810
rect 10876 10746 10928 10752
rect 11244 10746 11296 10752
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 12360 10606 12388 10950
rect 12636 10606 12664 11630
rect 12728 11218 12756 12174
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12912 10810 12940 19600
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13372 11694 13400 12242
rect 13556 11898 13584 19600
rect 14200 16574 14228 19600
rect 14844 16574 14872 19600
rect 14200 16546 14320 16574
rect 14844 16546 14964 16574
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13188 10606 13216 11154
rect 13740 10810 13768 11630
rect 14292 11354 14320 16546
rect 14936 12442 14964 16546
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 15488 12374 15516 19600
rect 16132 19258 16160 19600
rect 16776 19530 16804 19600
rect 16868 19530 16896 19638
rect 16776 19502 16896 19530
rect 16132 19230 16344 19258
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11762 16160 12174
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11642 16160 11698
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 15660 11620 15712 11626
rect 16132 11614 16252 11642
rect 15660 11562 15712 11568
rect 14936 11354 14964 11562
rect 15672 11354 15700 11562
rect 15807 11452 16115 11461
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15807 11387 16115 11396
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 16224 10810 16252 11614
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12452 10470 12480 10542
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 11150 10296 11206 10305
rect 11150 10231 11152 10240
rect 11204 10231 11206 10240
rect 11152 10202 11204 10208
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 12452 10130 12480 10406
rect 12544 10146 12572 10542
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10198 13032 10406
rect 13188 10266 13216 10542
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12992 10192 13044 10198
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12544 10118 12756 10146
rect 12992 10134 13044 10140
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 9140 9042 9168 9318
rect 9416 9042 9444 10066
rect 10060 9722 10088 10066
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 12360 9722 12388 9862
rect 12544 9722 12572 10118
rect 12728 10062 12756 10118
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12636 9908 12664 9998
rect 12636 9880 12848 9908
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 9770 9616 9826 9625
rect 9770 9551 9826 9560
rect 9784 9518 9812 9551
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 11808 9450 11836 9658
rect 12820 9602 12848 9880
rect 12912 9722 12940 9998
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12452 9574 12664 9602
rect 12820 9574 13032 9602
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 12084 9110 12112 9522
rect 12452 9450 12480 9574
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12440 9444 12492 9450
rect 12440 9386 12492 9392
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 9178 12388 9318
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 9680 9104 9732 9110
rect 12072 9104 12124 9110
rect 9680 9046 9732 9052
rect 11978 9072 12034 9081
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 9416 8634 9444 8978
rect 9692 8634 9720 9046
rect 12072 9046 12124 9052
rect 11978 9007 11980 9016
rect 12032 9007 12034 9016
rect 11980 8978 12032 8984
rect 11150 8936 11206 8945
rect 11150 8871 11206 8880
rect 12268 8888 12296 9114
rect 12544 9110 12572 9454
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12636 9042 12664 9574
rect 13004 9518 13032 9574
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12820 9382 12848 9454
rect 13096 9450 13124 10066
rect 13464 9926 13492 10474
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13464 9518 13492 9862
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13082 9072 13138 9081
rect 12624 9036 12676 9042
rect 13082 9007 13084 9016
rect 12624 8978 12676 8984
rect 13136 9007 13138 9016
rect 13084 8978 13136 8984
rect 12348 8900 12400 8906
rect 11164 8838 11192 8871
rect 12268 8860 12348 8888
rect 12348 8842 12400 8848
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 9416 7954 9444 8570
rect 10704 8430 10732 8774
rect 11808 8430 11836 8774
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 12544 8634 12572 8842
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 9968 8090 9996 8366
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 8129 10456 8298
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 10414 8120 10470 8129
rect 9956 8084 10008 8090
rect 10414 8055 10470 8064
rect 9956 8026 10008 8032
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 9770 7576 9826 7585
rect 9770 7511 9772 7520
rect 9824 7511 9826 7520
rect 9772 7482 9824 7488
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 9968 882 9996 8026
rect 10520 8022 10548 8230
rect 11716 8022 11744 8230
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 10060 7342 10088 7958
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7546 10824 7686
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 11716 7342 11744 7958
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 10888 2774 10916 7142
rect 11808 2774 11836 7142
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11955 6491 12263 6500
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 10888 2746 11008 2774
rect 9956 876 10008 882
rect 9956 818 10008 824
rect 9772 808 9824 814
rect 9772 750 9824 756
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 9784 490 9812 750
rect 9692 462 9812 490
rect 9692 400 9720 462
rect 10980 400 11008 2746
rect 11624 2746 11836 2774
rect 11624 400 11652 2746
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 12636 950 12664 8978
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13188 8634 13216 8842
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13372 8090 13400 8298
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 7954 13492 8774
rect 13556 8430 13584 9318
rect 13544 8424 13596 8430
rect 13542 8392 13544 8401
rect 13596 8392 13598 8401
rect 13542 8327 13598 8336
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13648 7818 13676 9998
rect 14016 9654 14044 10066
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13924 9110 13952 9454
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13832 8498 13860 8570
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13924 8430 13952 9046
rect 14016 9042 14044 9590
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14108 7954 14136 8366
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12624 944 12676 950
rect 12624 886 12676 892
rect 12256 740 12308 746
rect 12256 682 12308 688
rect 12268 400 12296 682
rect 12912 400 12940 7686
rect 13648 7342 13676 7754
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7342 13860 7686
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13832 6934 13860 7278
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 400 13584 6598
rect 14292 2774 14320 9318
rect 14384 9042 14412 9862
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14476 9178 14504 9386
rect 14568 9178 14596 10610
rect 15807 10364 16115 10373
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 16316 10266 16344 19230
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16868 11898 16896 12310
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16592 11218 16620 11630
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14660 9518 14688 10134
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 15934 9616 15990 9625
rect 15934 9551 15990 9560
rect 15948 9518 15976 9551
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 15384 9512 15436 9518
rect 15660 9512 15712 9518
rect 15384 9454 15436 9460
rect 15658 9480 15660 9489
rect 15936 9512 15988 9518
rect 15712 9480 15714 9489
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14568 8430 14596 9114
rect 15396 9110 15424 9454
rect 15936 9454 15988 9460
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 15658 9415 15714 9424
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 16224 9178 16252 9454
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 15384 9104 15436 9110
rect 16224 9058 16252 9114
rect 15384 9046 15436 9052
rect 16132 9042 16252 9058
rect 16316 9042 16344 9658
rect 16396 9648 16448 9654
rect 16448 9608 16528 9636
rect 16396 9590 16448 9596
rect 16500 9518 16528 9608
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16592 9178 16620 11018
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16776 10538 16804 10950
rect 16868 10674 16896 10950
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16776 9722 16804 10066
rect 16764 9716 16816 9722
rect 16816 9676 16896 9704
rect 16764 9658 16816 9664
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16684 9489 16712 9522
rect 16670 9480 16726 9489
rect 16868 9450 16896 9676
rect 17052 9654 17080 19638
rect 17406 19600 17462 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 19338 19600 19394 20000
rect 19982 19600 20038 20000
rect 20626 19600 20682 20000
rect 17420 12434 17448 19600
rect 18064 16574 18092 19600
rect 18708 16574 18736 19600
rect 18064 16546 18368 16574
rect 18708 16546 18828 16574
rect 17420 12406 17724 12434
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17144 11218 17172 11562
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11354 17632 11494
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17696 11286 17724 12406
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18248 11898 18276 12174
rect 18236 11892 18288 11898
rect 18156 11852 18236 11880
rect 18156 11694 18184 11852
rect 18236 11834 18288 11840
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 18340 10266 18368 16546
rect 18800 11898 18828 16546
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11898 19012 12242
rect 19064 12096 19116 12102
rect 19116 12044 19288 12050
rect 19064 12038 19288 12044
rect 19076 12022 19288 12038
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19260 11694 19288 12022
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11014 18828 11494
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10606 18828 10950
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18708 10062 18736 10542
rect 19260 10062 19288 11630
rect 19352 11354 19380 19600
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19628 11286 19656 11562
rect 19616 11280 19668 11286
rect 19616 11222 19668 11228
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17406 9616 17462 9625
rect 17406 9551 17408 9560
rect 17460 9551 17462 9560
rect 17408 9522 17460 9528
rect 16670 9415 16726 9424
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 16684 9178 16712 9318
rect 17972 9178 18000 9318
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 16592 9058 16620 9114
rect 16592 9042 16804 9058
rect 16120 9036 16252 9042
rect 16172 9030 16252 9036
rect 16304 9036 16356 9042
rect 16120 8978 16172 8984
rect 16592 9036 16816 9042
rect 16592 9030 16764 9036
rect 16304 8978 16356 8984
rect 16764 8978 16816 8984
rect 18248 8974 18276 9862
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14660 8498 14688 8842
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 15304 8430 15332 8774
rect 16316 8634 16344 8774
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14832 8424 14884 8430
rect 15200 8424 15252 8430
rect 14832 8366 14884 8372
rect 15198 8392 15200 8401
rect 15292 8424 15344 8430
rect 15252 8392 15254 8401
rect 14844 8294 14872 8366
rect 15292 8366 15344 8372
rect 15198 8327 15254 8336
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14568 8090 14596 8230
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15807 8123 16115 8132
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7410 15056 7686
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15304 7342 15332 7958
rect 16408 7954 16436 8570
rect 17604 8566 17632 8774
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17696 8498 17724 8774
rect 18248 8566 18276 8910
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16592 8022 16620 8230
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14936 6934 14964 7142
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15028 2774 15056 6598
rect 14200 2746 14320 2774
rect 14844 2746 15056 2774
rect 14200 400 14228 2746
rect 14844 400 14872 2746
rect 15488 400 15516 7686
rect 16592 7342 16620 7958
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 16592 6934 16620 7142
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 16316 474 16344 6598
rect 16028 468 16080 474
rect 16304 468 16356 474
rect 16080 428 16160 456
rect 16028 410 16080 416
rect 16132 400 16160 428
rect 16304 410 16356 416
rect 16776 400 16804 7142
rect 17420 400 17448 8298
rect 18248 7954 18276 8502
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 400 18092 7686
rect 18708 400 18736 8774
rect 19352 8634 19380 11154
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 19996 10810 20024 19600
rect 20640 12442 20668 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 31217 19068 31525 19077
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 31217 13628 31525 13637
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 28262 11656 28318 11665
rect 28262 11591 28264 11600
rect 28316 11591 28318 11600
rect 28264 11562 28316 11568
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 27365 10908 27673 10917
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31666 10296 31722 10305
rect 31666 10231 31722 10240
rect 31680 10130 31708 10231
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 31668 10124 31720 10130
rect 31668 10066 31720 10072
rect 19444 9518 19472 10066
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 28262 9616 28318 9625
rect 28262 9551 28318 9560
rect 28276 9518 28304 9551
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 28264 9512 28316 9518
rect 28264 9454 28316 9460
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20088 9178 20116 9386
rect 28264 9376 28316 9382
rect 28264 9318 28316 9324
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 21376 8634 21404 8978
rect 28276 8945 28304 9318
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 31217 9211 31525 9220
rect 28262 8936 28318 8945
rect 28262 8871 28318 8880
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 18880 8288 18932 8294
rect 31680 8265 31708 8774
rect 18880 8230 18932 8236
rect 31666 8256 31722 8265
rect 18892 8022 18920 8230
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 31217 8188 31525 8197
rect 31666 8191 31722 8200
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 31217 8123 31525 8132
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18892 7342 18920 7958
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19352 400 19380 7210
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 20640 400 20668 7686
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 27365 7579 27673 7588
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 27365 5468 27673 5477
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 31217 2748 31525 2757
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 9678 0 9734 400
rect 10966 0 11022 400
rect 11610 0 11666 400
rect 12254 0 12310 400
rect 12898 0 12954 400
rect 13542 0 13598 400
rect 14186 0 14242 400
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16118 0 16174 400
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 18050 0 18106 400
rect 18694 0 18750 400
rect 19338 0 19394 400
rect 20626 0 20682 400
<< via2 >>
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 11426 11600 11482 11656
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 10874 10804 10930 10840
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 10874 10784 10876 10804
rect 10876 10784 10928 10804
rect 10928 10784 10930 10804
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 11150 10260 11206 10296
rect 11150 10240 11152 10260
rect 11152 10240 11204 10260
rect 11204 10240 11206 10260
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 9770 9560 9826 9616
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 11978 9036 12034 9072
rect 11978 9016 11980 9036
rect 11980 9016 12032 9036
rect 12032 9016 12034 9036
rect 11150 8880 11206 8936
rect 13082 9036 13138 9072
rect 13082 9016 13084 9036
rect 13084 9016 13136 9036
rect 13136 9016 13138 9036
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 10414 8064 10470 8120
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 9770 7540 9826 7576
rect 9770 7520 9772 7540
rect 9772 7520 9824 7540
rect 9824 7520 9826 7540
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 13542 8372 13544 8392
rect 13544 8372 13596 8392
rect 13596 8372 13598 8392
rect 13542 8336 13598 8372
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 15934 9560 15990 9616
rect 15658 9460 15660 9480
rect 15660 9460 15712 9480
rect 15712 9460 15714 9480
rect 15658 9424 15714 9460
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 16670 9424 16726 9480
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 17406 9580 17462 9616
rect 17406 9560 17408 9580
rect 17408 9560 17460 9580
rect 17460 9560 17462 9580
rect 15198 8372 15200 8392
rect 15200 8372 15252 8392
rect 15252 8372 15254 8392
rect 15198 8336 15254 8372
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 28262 11620 28318 11656
rect 28262 11600 28264 11620
rect 28264 11600 28316 11620
rect 28316 11600 28318 11620
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10240 31722 10296
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 28262 9560 28318 9616
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 28262 8880 28318 8936
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 31666 8200 31722 8256
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
<< metal3 >>
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31213 19007 31529 19008
rect 4246 18528 4562 18529
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31213 13567 31529 13568
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 0 11658 400 11688
rect 11421 11658 11487 11661
rect 0 11656 11487 11658
rect 0 11600 11426 11656
rect 11482 11600 11487 11656
rect 0 11598 11487 11600
rect 0 11568 400 11598
rect 11421 11595 11487 11598
rect 28257 11658 28323 11661
rect 31600 11658 32000 11688
rect 28257 11656 32000 11658
rect 28257 11600 28262 11656
rect 28318 11600 32000 11656
rect 28257 11598 32000 11600
rect 28257 11595 28323 11598
rect 31600 11568 32000 11598
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 0 10978 400 11008
rect 0 10918 2790 10978
rect 0 10888 400 10918
rect 2730 10706 2790 10918
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 27361 10847 27677 10848
rect 10869 10842 10935 10845
rect 4662 10840 10935 10842
rect 4662 10784 10874 10840
rect 10930 10784 10935 10840
rect 4662 10782 10935 10784
rect 4662 10706 4722 10782
rect 10869 10779 10935 10782
rect 2730 10646 4722 10706
rect 8098 10368 8414 10369
rect 0 10298 400 10328
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 11145 10298 11211 10301
rect 0 10238 2790 10298
rect 0 10208 400 10238
rect 2730 10162 2790 10238
rect 8526 10296 11211 10298
rect 8526 10240 11150 10296
rect 11206 10240 11211 10296
rect 8526 10238 11211 10240
rect 8526 10162 8586 10238
rect 11145 10235 11211 10238
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 2730 10102 8586 10162
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 0 9618 400 9648
rect 9765 9618 9831 9621
rect 0 9616 9831 9618
rect 0 9560 9770 9616
rect 9826 9560 9831 9616
rect 0 9558 9831 9560
rect 0 9528 400 9558
rect 9765 9555 9831 9558
rect 15929 9618 15995 9621
rect 17401 9618 17467 9621
rect 15929 9616 17467 9618
rect 15929 9560 15934 9616
rect 15990 9560 17406 9616
rect 17462 9560 17467 9616
rect 15929 9558 17467 9560
rect 15929 9555 15995 9558
rect 17401 9555 17467 9558
rect 28257 9618 28323 9621
rect 31600 9618 32000 9648
rect 28257 9616 32000 9618
rect 28257 9560 28262 9616
rect 28318 9560 32000 9616
rect 28257 9558 32000 9560
rect 28257 9555 28323 9558
rect 31600 9528 32000 9558
rect 15653 9482 15719 9485
rect 16665 9482 16731 9485
rect 15653 9480 16731 9482
rect 15653 9424 15658 9480
rect 15714 9424 16670 9480
rect 16726 9424 16731 9480
rect 15653 9422 16731 9424
rect 15653 9419 15719 9422
rect 16665 9419 16731 9422
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 11973 9074 12039 9077
rect 13077 9074 13143 9077
rect 11973 9072 13143 9074
rect 11973 9016 11978 9072
rect 12034 9016 13082 9072
rect 13138 9016 13143 9072
rect 11973 9014 13143 9016
rect 11973 9011 12039 9014
rect 13077 9011 13143 9014
rect 0 8938 400 8968
rect 11145 8938 11211 8941
rect 0 8936 11211 8938
rect 0 8880 11150 8936
rect 11206 8880 11211 8936
rect 0 8878 11211 8880
rect 0 8848 400 8878
rect 11145 8875 11211 8878
rect 28257 8938 28323 8941
rect 31600 8938 32000 8968
rect 28257 8936 32000 8938
rect 28257 8880 28262 8936
rect 28318 8880 32000 8936
rect 28257 8878 32000 8880
rect 28257 8875 28323 8878
rect 31600 8848 32000 8878
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 13537 8394 13603 8397
rect 15193 8394 15259 8397
rect 13537 8392 15259 8394
rect 13537 8336 13542 8392
rect 13598 8336 15198 8392
rect 15254 8336 15259 8392
rect 13537 8334 15259 8336
rect 13537 8331 13603 8334
rect 15193 8331 15259 8334
rect 0 8258 400 8288
rect 0 8198 2790 8258
rect 0 8168 400 8198
rect 2730 7986 2790 8198
rect 31600 8256 32000 8288
rect 31600 8200 31666 8256
rect 31722 8200 32000 8256
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31600 8168 32000 8200
rect 31213 8127 31529 8128
rect 10409 8122 10475 8125
rect 10366 8120 10475 8122
rect 10366 8064 10414 8120
rect 10470 8064 10475 8120
rect 10366 8059 10475 8064
rect 10366 7986 10426 8059
rect 2730 7926 10426 7986
rect 4246 7648 4562 7649
rect 0 7578 400 7608
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 9765 7578 9831 7581
rect 0 7518 2790 7578
rect 0 7488 400 7518
rect 2730 7442 2790 7518
rect 4662 7576 9831 7578
rect 4662 7520 9770 7576
rect 9826 7520 9831 7576
rect 4662 7518 9831 7520
rect 4662 7442 4722 7518
rect 9765 7515 9831 7518
rect 2730 7382 4722 7442
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 27361 5407 27677 5408
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11949 12000 12269 13024
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 11949 8736 12269 9760
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 11949 6560 12269 7584
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 15801 15808 16121 16832
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 15801 10368 16121 11392
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15801 4928 16121 5952
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15801 3840 16121 4864
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19654 12000 19974 13024
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19654 7648 19974 8672
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 19654 4384 19974 5408
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 23506 15808 23826 16832
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
use sky130_fd_sc_hd__or2_1  _18_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 17112 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _19_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _20_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18032 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _21_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14996 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _22_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18584 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _23_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17204 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _24_
timestamp 1701704242
transform 1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _25_
timestamp 1701704242
transform 1 0 15548 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _26_
timestamp 1701704242
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _27_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14996 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _28_
timestamp 1701704242
transform 1 0 9384 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _29_
timestamp 1701704242
transform 1 0 9384 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _30_
timestamp 1701704242
transform 1 0 12604 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _31_
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _32_
timestamp 1701704242
transform 1 0 19412 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _33_
timestamp 1701704242
transform 1 0 18676 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _34_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15916 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _35_
timestamp 1701704242
transform 1 0 14628 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _36_
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _37_
timestamp 1701704242
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _38_
timestamp 1701704242
transform 1 0 16652 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _39_
timestamp 1701704242
transform 1 0 18308 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _40_
timestamp 1701704242
transform 1 0 18768 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _41_
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _42_
timestamp 1701704242
transform 1 0 11224 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _43_
timestamp 1701704242
transform 1 0 9384 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _44_
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _45_
timestamp 1701704242
transform 1 0 14352 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _46_
timestamp 1701704242
transform 1 0 19320 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _47_
timestamp 1701704242
transform 1 0 19412 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _48_
timestamp 1701704242
transform 1 0 16744 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _59_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13156 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1701704242
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _61_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18768 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _62_
timestamp 1701704242
transform 1 0 19504 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _63_
timestamp 1701704242
transform -1 0 19228 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _64_
timestamp 1701704242
transform -1 0 14260 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _65_
timestamp 1701704242
transform 1 0 16744 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _66_
timestamp 1701704242
transform 1 0 17756 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _67_
timestamp 1701704242
transform 1 0 18860 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _68_
timestamp 1701704242
transform 1 0 13708 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _69_
timestamp 1701704242
transform 1 0 11592 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _70_
timestamp 1701704242
transform -1 0 10304 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _71_
timestamp 1701704242
transform -1 0 11316 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _72_
timestamp 1701704242
transform 1 0 14536 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _73_
timestamp 1701704242
transform 1 0 19412 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _74_
timestamp 1701704242
transform -1 0 18492 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _75_
timestamp 1701704242
transform 1 0 16836 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _76_
timestamp 1701704242
transform 1 0 15088 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _77_
timestamp 1701704242
transform -1 0 10212 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _78_
timestamp 1701704242
transform 1 0 9936 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _79_
timestamp 1701704242
transform -1 0 13340 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _80_
timestamp 1701704242
transform 1 0 20148 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _81_
timestamp 1701704242
transform 1 0 20884 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _82_
timestamp 1701704242
transform 1 0 20148 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _83_
timestamp 1701704242
transform 1 0 14720 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _84_
timestamp 1701704242
transform 1 0 18124 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _85_
timestamp 1701704242
transform 1 0 19964 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _86_
timestamp 1701704242
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _87_
timestamp 1701704242
transform 1 0 14812 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _88_
timestamp 1701704242
transform 1 0 12696 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _89_
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _90_
timestamp 1701704242
transform -1 0 12328 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _91_
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _92_
timestamp 1701704242
transform 1 0 21252 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _93_
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _94_
timestamp 1701704242
transform 1 0 18216 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _95_
timestamp 1701704242
transform 1 0 16468 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _96_
timestamp 1701704242
transform 1 0 10672 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _97_
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _98_
timestamp 1701704242
transform 1 0 14076 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _99_
timestamp 1701704242
transform -1 0 12788 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout3
timestamp 1701704242
transform -1 0 12512 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout4
timestamp 1701704242
transform -1 0 12788 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout5 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout6
timestamp 1701704242
transform 1 0 15640 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout7
timestamp 1701704242
transform -1 0 9844 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1701704242
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10672 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_125
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_132 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12696 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1701704242
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1701704242
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1701704242
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1701704242
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1701704242
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1701704242
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1701704242
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_329
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1701704242
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1701704242
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1701704242
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1701704242
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1701704242
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1701704242
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1701704242
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1701704242
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1701704242
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1701704242
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1701704242
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1701704242
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1701704242
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1701704242
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1701704242
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1701704242
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1701704242
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1701704242
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1701704242
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1701704242
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1701704242
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1701704242
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1701704242
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1701704242
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1701704242
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1701704242
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1701704242
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1701704242
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1701704242
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1701704242
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1701704242
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1701704242
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1701704242
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1701704242
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1701704242
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1701704242
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1701704242
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1701704242
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1701704242
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1701704242
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1701704242
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_329
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1701704242
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1701704242
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1701704242
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1701704242
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1701704242
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1701704242
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1701704242
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1701704242
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1701704242
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1701704242
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1701704242
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1701704242
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1701704242
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1701704242
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1701704242
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1701704242
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1701704242
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1701704242
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1701704242
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1701704242
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1701704242
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1701704242
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1701704242
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1701704242
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1701704242
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1701704242
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1701704242
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1701704242
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1701704242
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1701704242
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1701704242
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1701704242
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1701704242
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1701704242
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1701704242
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1701704242
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1701704242
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1701704242
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1701704242
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1701704242
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1701704242
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1701704242
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1701704242
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_329
timestamp 1701704242
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1701704242
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1701704242
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1701704242
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1701704242
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1701704242
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1701704242
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1701704242
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1701704242
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1701704242
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1701704242
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1701704242
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1701704242
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1701704242
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1701704242
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1701704242
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1701704242
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1701704242
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1701704242
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1701704242
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1701704242
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1701704242
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_329
timestamp 1701704242
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1701704242
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1701704242
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1701704242
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1701704242
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1701704242
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1701704242
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1701704242
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1701704242
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1701704242
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1701704242
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1701704242
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1701704242
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1701704242
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1701704242
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1701704242
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1701704242
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1701704242
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1701704242
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1701704242
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1701704242
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1701704242
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1701704242
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1701704242
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1701704242
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 1701704242
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_329
timestamp 1701704242
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1701704242
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1701704242
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1701704242
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1701704242
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1701704242
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1701704242
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1701704242
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1701704242
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1701704242
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1701704242
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1701704242
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1701704242
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1701704242
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1701704242
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1701704242
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1701704242
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1701704242
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1701704242
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1701704242
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1701704242
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1701704242
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1701704242
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1701704242
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1701704242
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1701704242
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1701704242
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_329
timestamp 1701704242
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1701704242
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1701704242
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1701704242
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1701704242
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1701704242
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1701704242
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1701704242
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1701704242
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1701704242
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1701704242
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1701704242
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1701704242
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1701704242
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1701704242
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1701704242
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1701704242
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1701704242
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1701704242
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1701704242
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1701704242
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1701704242
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1701704242
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1701704242
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1701704242
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1701704242
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1701704242
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_321
timestamp 1701704242
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 1701704242
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1701704242
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1701704242
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1701704242
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1701704242
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1701704242
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1701704242
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1701704242
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_137
timestamp 1701704242
transform 1 0 13156 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_149
timestamp 1701704242
transform 1 0 14260 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1701704242
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1701704242
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_179
timestamp 1701704242
transform 1 0 17020 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_191
timestamp 1701704242
transform 1 0 18124 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_203
timestamp 1701704242
transform 1 0 19228 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_215
timestamp 1701704242
transform 1 0 20332 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1701704242
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1701704242
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1701704242
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1701704242
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1701704242
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1701704242
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1701704242
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1701704242
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1701704242
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_329
timestamp 1701704242
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1701704242
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1701704242
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1701704242
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1701704242
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1701704242
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1701704242
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1701704242
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_97
timestamp 1701704242
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_105
timestamp 1701704242
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_109
timestamp 1701704242
transform 1 0 10580 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_116
timestamp 1701704242
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_126
timestamp 1701704242
transform 1 0 12144 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1701704242
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_173
timestamp 1701704242
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_183
timestamp 1701704242
transform 1 0 17388 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1701704242
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_205
timestamp 1701704242
transform 1 0 19412 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_217
timestamp 1701704242
transform 1 0 20516 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_229
timestamp 1701704242
transform 1 0 21620 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_241
timestamp 1701704242
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1701704242
transform 1 0 23460 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1701704242
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1701704242
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1701704242
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1701704242
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1701704242
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1701704242
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_321
timestamp 1701704242
transform 1 0 30084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_329
timestamp 1701704242
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1701704242
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1701704242
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1701704242
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1701704242
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1701704242
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1701704242
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_93
timestamp 1701704242
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_138
timestamp 1701704242
transform 1 0 13248 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_145
timestamp 1701704242
transform 1 0 13892 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_153
timestamp 1701704242
transform 1 0 14628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_157
timestamp 1701704242
transform 1 0 14996 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_169
timestamp 1701704242
transform 1 0 16100 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_175
timestamp 1701704242
transform 1 0 16652 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1701704242
transform 1 0 20792 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1701704242
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1701704242
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1701704242
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1701704242
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1701704242
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1701704242
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1701704242
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1701704242
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1701704242
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_329
timestamp 1701704242
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1701704242
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1701704242
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1701704242
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_101
timestamp 1701704242
transform 1 0 9844 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_111
timestamp 1701704242
transform 1 0 10764 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_119
timestamp 1701704242
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_124
timestamp 1701704242
transform 1 0 11960 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_148
timestamp 1701704242
transform 1 0 14168 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_163
timestamp 1701704242
transform 1 0 15548 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_171
timestamp 1701704242
transform 1 0 16284 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_175
timestamp 1701704242
transform 1 0 16652 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_187
timestamp 1701704242
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1701704242
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_200
timestamp 1701704242
transform 1 0 18952 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_204
timestamp 1701704242
transform 1 0 19320 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1701704242
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1701704242
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1701704242
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1701704242
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1701704242
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1701704242
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1701704242
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1701704242
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1701704242
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1701704242
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_321
timestamp 1701704242
transform 1 0 30084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_329
timestamp 1701704242
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1701704242
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1701704242
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1701704242
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1701704242
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_119
timestamp 1701704242
transform 1 0 11500 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_139
timestamp 1701704242
transform 1 0 13340 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_143
timestamp 1701704242
transform 1 0 13708 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_152
timestamp 1701704242
transform 1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_158
timestamp 1701704242
transform 1 0 15088 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_164
timestamp 1701704242
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_186
timestamp 1701704242
transform 1 0 17664 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_209
timestamp 1701704242
transform 1 0 19780 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1701704242
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_231
timestamp 1701704242
transform 1 0 21804 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_243
timestamp 1701704242
transform 1 0 22908 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_255
timestamp 1701704242
transform 1 0 24012 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_267
timestamp 1701704242
transform 1 0 25116 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1701704242
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1701704242
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1701704242
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1701704242
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1701704242
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_329
timestamp 1701704242
transform 1 0 30820 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1701704242
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1701704242
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1701704242
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1701704242
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1701704242
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_97
timestamp 1701704242
transform 1 0 9476 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_109
timestamp 1701704242
transform 1 0 10580 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_117
timestamp 1701704242
transform 1 0 11316 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1701704242
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_158
timestamp 1701704242
transform 1 0 15088 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_185
timestamp 1701704242
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_190
timestamp 1701704242
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_197
timestamp 1701704242
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_202
timestamp 1701704242
transform 1 0 19136 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_217
timestamp 1701704242
transform 1 0 20516 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_229
timestamp 1701704242
transform 1 0 21620 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_241
timestamp 1701704242
transform 1 0 22724 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_249
timestamp 1701704242
transform 1 0 23460 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1701704242
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1701704242
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1701704242
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1701704242
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1701704242
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1701704242
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1701704242
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1701704242
transform 1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_329
timestamp 1701704242
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1701704242
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1701704242
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1701704242
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1701704242
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_93
timestamp 1701704242
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_119
timestamp 1701704242
transform 1 0 11500 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_141
timestamp 1701704242
transform 1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1701704242
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_197
timestamp 1701704242
transform 1 0 18676 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_203
timestamp 1701704242
transform 1 0 19228 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_220
timestamp 1701704242
transform 1 0 20792 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_231
timestamp 1701704242
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_243
timestamp 1701704242
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_255
timestamp 1701704242
transform 1 0 24012 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_267
timestamp 1701704242
transform 1 0 25116 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1701704242
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1701704242
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1701704242
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1701704242
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_329
timestamp 1701704242
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1701704242
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1701704242
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1701704242
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1701704242
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1701704242
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1701704242
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1701704242
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_109
timestamp 1701704242
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_120
timestamp 1701704242
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_128
timestamp 1701704242
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1701704242
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_149
timestamp 1701704242
transform 1 0 14260 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_161
timestamp 1701704242
transform 1 0 15364 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_187
timestamp 1701704242
transform 1 0 17756 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1701704242
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_219
timestamp 1701704242
transform 1 0 20700 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_231
timestamp 1701704242
transform 1 0 21804 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_243
timestamp 1701704242
transform 1 0 22908 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1701704242
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1701704242
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1701704242
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1701704242
transform 1 0 27140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1701704242
transform 1 0 28244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1701704242
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_321
timestamp 1701704242
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_329
timestamp 1701704242
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1701704242
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1701704242
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1701704242
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1701704242
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1701704242
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1701704242
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1701704242
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1701704242
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1701704242
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_129
timestamp 1701704242
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_153
timestamp 1701704242
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_160
timestamp 1701704242
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1701704242
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_169
timestamp 1701704242
transform 1 0 16100 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_181
timestamp 1701704242
transform 1 0 17204 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_189
timestamp 1701704242
transform 1 0 17940 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_198
timestamp 1701704242
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_216
timestamp 1701704242
transform 1 0 20424 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1701704242
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1701704242
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1701704242
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1701704242
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1701704242
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1701704242
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1701704242
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1701704242
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1701704242
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1701704242
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_329
timestamp 1701704242
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1701704242
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1701704242
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1701704242
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1701704242
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1701704242
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1701704242
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1701704242
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_109
timestamp 1701704242
transform 1 0 10580 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1701704242
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_149
timestamp 1701704242
transform 1 0 14260 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_173
timestamp 1701704242
transform 1 0 16468 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_177
timestamp 1701704242
transform 1 0 16836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1701704242
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_203
timestamp 1701704242
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_227
timestamp 1701704242
transform 1 0 21436 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_239
timestamp 1701704242
transform 1 0 22540 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1701704242
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1701704242
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1701704242
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1701704242
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1701704242
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1701704242
transform 1 0 28244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1701704242
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1701704242
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_329
timestamp 1701704242
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1701704242
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1701704242
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1701704242
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1701704242
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1701704242
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1701704242
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_125
timestamp 1701704242
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_132
timestamp 1701704242
transform 1 0 12696 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_160
timestamp 1701704242
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_196
timestamp 1701704242
transform 1 0 18584 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_219
timestamp 1701704242
transform 1 0 20700 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1701704242
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1701704242
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1701704242
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1701704242
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1701704242
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1701704242
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1701704242
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1701704242
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1701704242
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1701704242
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_329
timestamp 1701704242
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1701704242
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1701704242
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1701704242
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1701704242
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1701704242
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1701704242
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1701704242
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1701704242
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1701704242
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1701704242
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1701704242
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1701704242
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1701704242
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1701704242
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1701704242
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1701704242
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1701704242
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1701704242
transform 1 0 20884 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1701704242
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1701704242
transform 1 0 23092 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1701704242
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1701704242
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1701704242
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1701704242
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1701704242
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1701704242
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 1701704242
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1701704242
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1701704242
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1701704242
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1701704242
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1701704242
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1701704242
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1701704242
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1701704242
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1701704242
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1701704242
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1701704242
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1701704242
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1701704242
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1701704242
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1701704242
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1701704242
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1701704242
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1701704242
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1701704242
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1701704242
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1701704242
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1701704242
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1701704242
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1701704242
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1701704242
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1701704242
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1701704242
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1701704242
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1701704242
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_329
timestamp 1701704242
transform 1 0 30820 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1701704242
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1701704242
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1701704242
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1701704242
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1701704242
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1701704242
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1701704242
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1701704242
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1701704242
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1701704242
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1701704242
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1701704242
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1701704242
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1701704242
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1701704242
transform 1 0 17940 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1701704242
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1701704242
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1701704242
transform 1 0 20884 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1701704242
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1701704242
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1701704242
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1701704242
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1701704242
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1701704242
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1701704242
transform 1 0 27140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1701704242
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1701704242
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 1701704242
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_329
timestamp 1701704242
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1701704242
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1701704242
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1701704242
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1701704242
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1701704242
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1701704242
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1701704242
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1701704242
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1701704242
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1701704242
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1701704242
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1701704242
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1701704242
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1701704242
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1701704242
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1701704242
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1701704242
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1701704242
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1701704242
transform 1 0 20516 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1701704242
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1701704242
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1701704242
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1701704242
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1701704242
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1701704242
transform 1 0 25668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1701704242
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1701704242
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1701704242
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1701704242
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_329
timestamp 1701704242
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1701704242
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1701704242
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1701704242
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1701704242
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1701704242
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1701704242
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1701704242
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1701704242
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1701704242
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1701704242
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1701704242
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1701704242
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1701704242
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1701704242
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1701704242
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1701704242
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1701704242
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1701704242
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1701704242
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1701704242
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1701704242
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1701704242
transform 1 0 23092 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1701704242
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1701704242
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1701704242
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1701704242
transform 1 0 27140 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1701704242
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1701704242
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1701704242
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1701704242
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1701704242
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1701704242
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1701704242
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1701704242
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1701704242
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1701704242
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1701704242
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1701704242
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1701704242
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1701704242
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1701704242
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1701704242
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1701704242
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1701704242
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1701704242
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1701704242
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1701704242
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1701704242
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1701704242
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1701704242
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1701704242
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1701704242
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1701704242
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_329
timestamp 1701704242
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1701704242
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1701704242
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1701704242
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1701704242
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1701704242
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1701704242
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1701704242
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1701704242
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1701704242
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1701704242
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1701704242
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1701704242
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1701704242
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1701704242
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1701704242
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1701704242
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1701704242
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1701704242
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1701704242
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1701704242
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1701704242
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1701704242
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1701704242
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1701704242
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1701704242
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1701704242
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1701704242
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1701704242
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1701704242
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1701704242
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1701704242
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1701704242
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1701704242
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1701704242
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1701704242
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1701704242
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1701704242
transform 1 0 20516 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1701704242
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1701704242
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1701704242
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1701704242
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1701704242
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1701704242
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1701704242
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1701704242
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1701704242
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1701704242
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1701704242
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1701704242
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1701704242
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1701704242
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1701704242
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1701704242
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1701704242
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1701704242
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1701704242
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1701704242
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1701704242
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1701704242
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1701704242
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1701704242
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1701704242
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1701704242
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1701704242
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1701704242
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1701704242
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1701704242
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1701704242
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1701704242
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1701704242
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1701704242
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1701704242
transform 1 0 20516 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1701704242
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1701704242
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1701704242
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1701704242
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1701704242
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1701704242
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1701704242
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1701704242
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1701704242
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1701704242
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1701704242
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1701704242
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1701704242
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1701704242
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1701704242
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1701704242
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1701704242
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1701704242
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1701704242
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_137
timestamp 1701704242
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_153
timestamp 1701704242
transform 1 0 14628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1701704242
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 1701704242
transform 1 0 19780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1701704242
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22356 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_249
timestamp 1701704242
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1701704242
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1701704242
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_305
timestamp 1701704242
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_329
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  g_buf2.ctr_buf pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13984 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  g_dly_stp\[0\].dly_stp
timestamp 1701704242
transform -1 0 11592 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  g_dly_stp\[1\].dly_stp
timestamp 1701704242
transform -1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  g_dly_stp\[2\].dly_stp
timestamp 1701704242
transform 1 0 11868 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  g_ring1\[1\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 16744 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring1\[1\].stg01 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13800 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring1\[1\].stg02 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14168 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring1\[2\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring1\[2\].stg01
timestamp 1701704242
transform -1 0 15456 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring1\[2\].stg02
timestamp 1701704242
transform -1 0 16100 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring1\[3\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 18952 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring1\[3\].stg01
timestamp 1701704242
transform 1 0 15732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring1\[3\].stg02
timestamp 1701704242
transform -1 0 16836 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring1\[4\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 13892 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring1\[4\].stg01
timestamp 1701704242
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring1\[4\].stg02
timestamp 1701704242
transform -1 0 15272 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring1\[5\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring1\[5\].stg01
timestamp 1701704242
transform 1 0 13892 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring1\[5\].stg02
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring1\[6\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring1\[6\].stg01
timestamp 1701704242
transform 1 0 12788 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring1\[6\].stg02
timestamp 1701704242
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring1\[7\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring1\[7\].stg01
timestamp 1701704242
transform -1 0 11960 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring1\[7\].stg02
timestamp 1701704242
transform -1 0 12972 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring2\[8\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring2\[8\].stg01_8 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11868 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring2\[8\].stg01
timestamp 1701704242
transform 1 0 12972 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring2\[8\].stg02
timestamp 1701704242
transform -1 0 13248 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring3\[9\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 19136 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring3\[9\].stg01_15
timestamp 1701704242
transform 1 0 13800 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring3\[9\].stg01
timestamp 1701704242
transform -1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring3\[9\].stg02
timestamp 1701704242
transform 1 0 14168 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring3\[10\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 17664 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring3\[10\].stg01
timestamp 1701704242
transform 1 0 17296 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring3\[10\].stg01_9
timestamp 1701704242
transform 1 0 15456 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring3\[10\].stg02
timestamp 1701704242
transform 1 0 16100 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring3\[11\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 16652 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring3\[11\].stg01_10
timestamp 1701704242
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring3\[11\].stg01
timestamp 1701704242
transform 1 0 17112 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring3\[11\].stg02
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring3\[12\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 14996 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring3\[12\].stg01_11
timestamp 1701704242
transform 1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring3\[12\].stg01
timestamp 1701704242
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring3\[12\].stg02
timestamp 1701704242
transform 1 0 14536 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring3\[13\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 10488 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring3\[13\].stg01_12
timestamp 1701704242
transform -1 0 13708 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring3\[13\].stg01
timestamp 1701704242
transform 1 0 13340 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring3\[13\].stg02
timestamp 1701704242
transform 1 0 13064 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring3\[14\].g_buf2.ctr_buf
timestamp 1701704242
transform -1 0 9384 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring3\[14\].stg01_13
timestamp 1701704242
transform -1 0 13340 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring3\[14\].stg01
timestamp 1701704242
transform -1 0 12052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring3\[14\].stg02
timestamp 1701704242
transform -1 0 12420 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  g_ring3\[15\].g_buf2.ctr_buf
timestamp 1701704242
transform 1 0 13248 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  g_ring3\[15\].stg01_14
timestamp 1701704242
transform -1 0 12236 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_ring3\[15\].stg01
timestamp 1701704242
transform -1 0 11684 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  g_ring3\[15\].stg02
timestamp 1701704242
transform -1 0 12604 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1701704242
transform 1 0 12328 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9752 0 1 544
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stg01_16
timestamp 1701704242
transform -1 0 14260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  stg01
timestamp 1701704242
transform -1 0 11868 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  stg02
timestamp 1701704242
transform -1 0 12880 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 15474 19600 15530 20000 0 FreeSans 224 90 0 0 dbg_reset
port 2 nsew signal tristate
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[0]
port 3 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[1]
port 4 nsew signal tristate
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[2]
port 5 nsew signal tristate
flabel metal2 s 13542 19600 13598 20000 0 FreeSans 224 90 0 0 dbg_ring_sig[0]
port 6 nsew signal tristate
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 dbg_ring_sig[10]
port 7 nsew signal tristate
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 dbg_ring_sig[11]
port 8 nsew signal tristate
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 dbg_ring_sig[12]
port 9 nsew signal tristate
flabel metal3 s 0 7488 400 7608 0 FreeSans 480 0 0 0 dbg_ring_sig[13]
port 10 nsew signal tristate
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 dbg_ring_sig[14]
port 11 nsew signal tristate
flabel metal2 s 12898 19600 12954 20000 0 FreeSans 224 90 0 0 dbg_ring_sig[15]
port 12 nsew signal tristate
flabel metal2 s 16762 19600 16818 20000 0 FreeSans 224 90 0 0 dbg_ring_sig[1]
port 13 nsew signal tristate
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 dbg_ring_sig[2]
port 14 nsew signal tristate
flabel metal2 s 19338 0 19394 400 0 FreeSans 224 90 0 0 dbg_ring_sig[3]
port 15 nsew signal tristate
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 dbg_ring_sig[4]
port 16 nsew signal tristate
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 dbg_ring_sig[5]
port 17 nsew signal tristate
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 dbg_ring_sig[6]
port 18 nsew signal tristate
flabel metal3 s 0 10888 400 11008 0 FreeSans 480 0 0 0 dbg_ring_sig[7]
port 19 nsew signal tristate
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 dbg_ring_sig[8]
port 20 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 dbg_ring_sig[9]
port 21 nsew signal tristate
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 i_start
port 22 nsew signal input
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 i_stop
port 23 nsew signal input
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 o_result_ctr[0]
port 24 nsew signal tristate
flabel metal3 s 31600 11568 32000 11688 0 FreeSans 480 0 0 0 o_result_ctr[1]
port 25 nsew signal tristate
flabel metal2 s 20626 19600 20682 20000 0 FreeSans 224 90 0 0 o_result_ctr[2]
port 26 nsew signal tristate
flabel metal2 s 14830 19600 14886 20000 0 FreeSans 224 90 0 0 o_result_ring[0]
port 27 nsew signal tristate
flabel metal3 s 31600 8168 32000 8288 0 FreeSans 480 0 0 0 o_result_ring[10]
port 28 nsew signal tristate
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 o_result_ring[11]
port 29 nsew signal tristate
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 o_result_ring[12]
port 30 nsew signal tristate
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 o_result_ring[13]
port 31 nsew signal tristate
flabel metal3 s 0 8848 400 8968 0 FreeSans 480 0 0 0 o_result_ring[14]
port 32 nsew signal tristate
flabel metal2 s 14186 19600 14242 20000 0 FreeSans 224 90 0 0 o_result_ring[15]
port 33 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 o_result_ring[1]
port 34 nsew signal tristate
flabel metal3 s 31600 8848 32000 8968 0 FreeSans 480 0 0 0 o_result_ring[2]
port 35 nsew signal tristate
flabel metal2 s 20626 0 20682 400 0 FreeSans 224 90 0 0 o_result_ring[3]
port 36 nsew signal tristate
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 o_result_ring[4]
port 37 nsew signal tristate
flabel metal2 s 12898 0 12954 400 0 FreeSans 224 90 0 0 o_result_ring[5]
port 38 nsew signal tristate
flabel metal3 s 0 10208 400 10328 0 FreeSans 480 0 0 0 o_result_ring[6]
port 39 nsew signal tristate
flabel metal3 s 0 11568 400 11688 0 FreeSans 480 0 0 0 o_result_ring[7]
port 40 nsew signal tristate
flabel metal2 s 16118 19600 16174 20000 0 FreeSans 224 90 0 0 o_result_ring[8]
port 41 nsew signal tristate
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 o_result_ring[9]
port 42 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal1 16560 10642 16560 10642 0 _00_
rlabel metal1 14996 11322 14996 11322 0 _01_
rlabel metal1 17986 12172 17986 12172 0 _02_
rlabel metal2 16790 10744 16790 10744 0 _03_
rlabel metal2 15686 11458 15686 11458 0 _04_
rlabel metal1 16790 11866 16790 11866 0 _05_
rlabel metal1 17756 11730 17756 11730 0 _06_
rlabel metal1 18216 11866 18216 11866 0 _07_
rlabel metal1 15226 11220 15226 11220 0 _08_
rlabel metal1 13064 12342 13064 12342 0 dbg_reset
rlabel metal2 17434 16029 17434 16029 0 dbg_ring_ctr[0]
rlabel metal1 19550 11322 19550 11322 0 dbg_ring_ctr[1]
rlabel metal2 18722 18099 18722 18099 0 dbg_ring_ctr[2]
rlabel metal1 13708 11866 13708 11866 0 dbg_ring_sig[0]
rlabel metal1 17710 8330 17710 8330 0 dbg_ring_sig[10]
rlabel metal1 16928 7174 16928 7174 0 dbg_ring_sig[11]
rlabel metal2 15502 4036 15502 4036 0 dbg_ring_sig[12]
rlabel metal3 1533 7548 1533 7548 0 dbg_ring_sig[13]
rlabel metal3 1533 8228 1533 8228 0 dbg_ring_sig[14]
rlabel metal2 12926 15208 12926 15208 0 dbg_ring_sig[15]
rlabel metal2 16974 19652 16974 19652 0 dbg_ring_sig[1]
rlabel metal1 18446 8806 18446 8806 0 dbg_ring_sig[2]
rlabel metal2 19366 3798 19366 3798 0 dbg_ring_sig[3]
rlabel metal1 13754 6630 13754 6630 0 dbg_ring_sig[4]
rlabel metal2 11638 1557 11638 1557 0 dbg_ring_sig[5]
rlabel metal2 9798 9537 9798 9537 0 dbg_ring_sig[6]
rlabel metal3 1533 10948 1533 10948 0 dbg_ring_sig[7]
rlabel metal2 14214 1557 14214 1557 0 dbg_ring_sig[8]
rlabel metal2 28290 9537 28290 9537 0 dbg_ring_sig[9]
rlabel metal2 12282 534 12282 534 0 i_start
rlabel metal2 9706 415 9706 415 0 i_stop
rlabel metal1 12742 9010 12742 9010 0 net1
rlabel metal1 17112 9010 17112 9010 0 net10
rlabel metal2 15318 8602 15318 8602 0 net11
rlabel metal1 13432 7922 13432 7922 0 net12
rlabel via2 13110 9027 13110 9027 0 net13
rlabel metal1 11638 9520 11638 9520 0 net14
rlabel metal1 14444 9010 14444 9010 0 net15
rlabel metal2 13018 10302 13018 10302 0 net16
rlabel metal2 19366 9894 19366 9894 0 net2
rlabel via2 13570 8381 13570 8381 0 net3
rlabel metal2 12466 10268 12466 10268 0 net4
rlabel metal1 16100 11186 16100 11186 0 net5
rlabel metal1 15456 7786 15456 7786 0 net6
rlabel metal1 12696 11186 12696 11186 0 net7
rlabel metal1 12650 9996 12650 9996 0 net8
rlabel metal1 17342 9520 17342 9520 0 net9
rlabel metal1 20194 10778 20194 10778 0 o_result_ctr[0]
rlabel via2 28290 11611 28290 11611 0 o_result_ctr[1]
rlabel metal1 20608 12410 20608 12410 0 o_result_ctr[2]
rlabel metal2 14858 18099 14858 18099 0 o_result_ring[0]
rlabel metal2 31694 8517 31694 8517 0 o_result_ring[10]
rlabel metal1 18262 7718 18262 7718 0 o_result_ring[11]
rlabel metal1 16514 6630 16514 6630 0 o_result_ring[12]
rlabel metal2 10994 1557 10994 1557 0 o_result_ring[13]
rlabel metal2 11178 8857 11178 8857 0 o_result_ring[14]
rlabel metal2 14214 18099 14214 18099 0 o_result_ring[15]
rlabel metal2 18078 18099 18078 18099 0 o_result_ring[1]
rlabel metal1 21275 9418 21275 9418 0 o_result_ring[2]
rlabel metal2 20654 4036 20654 4036 0 o_result_ring[3]
rlabel metal2 14858 1557 14858 1557 0 o_result_ring[4]
rlabel metal2 12926 4036 12926 4036 0 o_result_ring[5]
rlabel metal3 1533 10268 1533 10268 0 o_result_ring[6]
rlabel metal2 11454 11203 11454 11203 0 o_result_ring[7]
rlabel metal2 16238 19244 16238 19244 0 o_result_ring[8]
rlabel metal2 31694 10183 31694 10183 0 o_result_ring[9]
rlabel metal1 20194 10506 20194 10506 0 r_dly_store_ctr\[0\]
rlabel metal1 20930 11594 20930 11594 0 r_dly_store_ctr\[1\]
rlabel metal1 20286 12376 20286 12376 0 r_dly_store_ctr\[2\]
rlabel metal1 14766 12342 14766 12342 0 r_dly_store_ring\[0\]
rlabel metal1 21114 8602 21114 8602 0 r_dly_store_ring\[10\]
rlabel metal1 18262 7990 18262 7990 0 r_dly_store_ring\[11\]
rlabel metal2 16606 7038 16606 7038 0 r_dly_store_ring\[12\]
rlabel metal1 10810 7412 10810 7412 0 r_dly_store_ring\[13\]
rlabel metal1 10948 9078 10948 9078 0 r_dly_store_ring\[14\]
rlabel metal1 14122 11254 14122 11254 0 r_dly_store_ring\[15\]
rlabel metal1 18170 10166 18170 10166 0 r_dly_store_ring\[1\]
rlabel metal1 19918 9146 19918 9146 0 r_dly_store_ring\[2\]
rlabel metal1 20378 8024 20378 8024 0 r_dly_store_ring\[3\]
rlabel metal2 14950 7038 14950 7038 0 r_dly_store_ring\[4\]
rlabel metal1 12742 7990 12742 7990 0 r_dly_store_ring\[5\]
rlabel metal1 10948 10166 10948 10166 0 r_dly_store_ring\[6\]
rlabel metal1 12282 10574 12282 10574 0 r_dly_store_ring\[7\]
rlabel metal1 16008 10166 16008 10166 0 r_dly_store_ring\[8\]
rlabel metal1 21390 10200 21390 10200 0 r_dly_store_ring\[9\]
rlabel metal1 18722 11186 18722 11186 0 r_ring_ctr\[0\]
rlabel metal2 19642 11424 19642 11424 0 r_ring_ctr\[1\]
rlabel metal1 18124 12274 18124 12274 0 r_ring_ctr\[2\]
rlabel metal1 11592 11662 11592 11662 0 w_dly_stop\[1\]
rlabel metal1 12006 11560 12006 11560 0 w_dly_stop\[2\]
rlabel metal1 15962 10710 15962 10710 0 w_ring_buf\[0\]
rlabel metal1 17986 8398 17986 8398 0 w_ring_buf\[10\]
rlabel metal1 16820 7990 16820 7990 0 w_ring_buf\[11\]
rlabel metal1 15088 7990 15088 7990 0 w_ring_buf\[12\]
rlabel metal1 10115 7990 10115 7990 0 w_ring_buf\[13\]
rlabel metal1 9506 9078 9506 9078 0 w_ring_buf\[14\]
rlabel metal2 13202 10880 13202 10880 0 w_ring_buf\[15\]
rlabel metal1 16744 9690 16744 9690 0 w_ring_buf\[1\]
rlabel metal1 17940 9078 17940 9078 0 w_ring_buf\[2\]
rlabel metal1 18982 7990 18982 7990 0 w_ring_buf\[3\]
rlabel via1 13841 7310 13841 7310 0 w_ring_buf\[4\]
rlabel metal1 11633 7990 11633 7990 0 w_ring_buf\[5\]
rlabel metal1 10212 9690 10212 9690 0 w_ring_buf\[6\]
rlabel metal1 11316 10778 11316 10778 0 w_ring_buf\[7\]
rlabel metal1 14474 10166 14474 10166 0 w_ring_buf\[8\]
rlabel metal1 19504 9486 19504 9486 0 w_ring_buf\[9\]
rlabel metal1 11822 9996 11822 9996 0 w_ring_int_norsz\[0\]
rlabel metal1 17204 9418 17204 9418 0 w_ring_int_norsz\[10\]
rlabel metal1 16836 8942 16836 8942 0 w_ring_int_norsz\[11\]
rlabel metal2 14858 8330 14858 8330 0 w_ring_int_norsz\[12\]
rlabel metal1 13432 8058 13432 8058 0 w_ring_int_norsz\[13\]
rlabel metal1 12006 8942 12006 8942 0 w_ring_int_norsz\[14\]
rlabel metal1 12052 9418 12052 9418 0 w_ring_int_norsz\[15\]
rlabel metal1 13754 9418 13754 9418 0 w_ring_int_norsz\[1\]
rlabel metal1 15548 9418 15548 9418 0 w_ring_int_norsz\[2\]
rlabel metal1 16192 9078 16192 9078 0 w_ring_int_norsz\[3\]
rlabel metal1 14674 8330 14674 8330 0 w_ring_int_norsz\[4\]
rlabel metal2 13846 8534 13846 8534 0 w_ring_int_norsz\[5\]
rlabel metal1 12834 8942 12834 8942 0 w_ring_int_norsz\[6\]
rlabel metal1 12650 9588 12650 9588 0 w_ring_int_norsz\[7\]
rlabel metal1 12972 9690 12972 9690 0 w_ring_int_norsz\[8\]
rlabel metal1 14444 9146 14444 9146 0 w_ring_int_norsz\[9\]
rlabel metal1 13524 9486 13524 9486 0 w_ring_norsz\[0\]
rlabel metal1 16698 9078 16698 9078 0 w_ring_norsz\[10\]
rlabel metal1 16376 8398 16376 8398 0 w_ring_norsz\[11\]
rlabel metal1 14674 7922 14674 7922 0 w_ring_norsz\[12\]
rlabel metal2 12558 8738 12558 8738 0 w_ring_norsz\[13\]
rlabel metal1 9154 9384 9154 9384 0 w_ring_norsz\[14\]
rlabel metal1 12926 9962 12926 9962 0 w_ring_norsz\[15\]
rlabel metal1 15226 9520 15226 9520 0 w_ring_norsz\[1\]
rlabel metal1 16284 9690 16284 9690 0 w_ring_norsz\[2\]
rlabel metal1 17250 8874 17250 8874 0 w_ring_norsz\[3\]
rlabel metal1 14122 8466 14122 8466 0 w_ring_norsz\[4\]
rlabel metal1 13018 8976 13018 8976 0 w_ring_norsz\[5\]
rlabel viali 11733 9486 11733 9486 0 w_ring_norsz\[6\]
rlabel metal1 12650 9690 12650 9690 0 w_ring_norsz\[7\]
rlabel metal1 13846 10098 13846 10098 0 w_ring_norsz\[8\]
rlabel metal1 15916 9486 15916 9486 0 w_ring_norsz\[9\]
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
