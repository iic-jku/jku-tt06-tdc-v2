magic
tech sky130A
magscale 1 2
timestamp 1710764608
<< viali >>
rect 12357 18785 12391 18819
rect 12541 18581 12575 18615
rect 13829 12733 13863 12767
rect 15485 12733 15519 12767
rect 17325 12733 17359 12767
rect 18889 12733 18923 12767
rect 13921 12597 13955 12631
rect 15577 12597 15611 12631
rect 17509 12597 17543 12631
rect 18797 12597 18831 12631
rect 12633 12393 12667 12427
rect 13185 12393 13219 12427
rect 19717 12393 19751 12427
rect 13522 12325 13556 12359
rect 17570 12325 17604 12359
rect 18981 12325 19015 12359
rect 11494 12257 11528 12291
rect 11667 12257 11701 12291
rect 11770 12256 11804 12290
rect 11897 12257 11931 12291
rect 12173 12257 12207 12291
rect 12449 12257 12483 12291
rect 12909 12257 12943 12291
rect 13001 12257 13035 12291
rect 13277 12257 13311 12291
rect 15033 12247 15067 12281
rect 15945 12257 15979 12291
rect 16773 12257 16807 12291
rect 16865 12257 16899 12291
rect 17049 12257 17083 12291
rect 19349 12257 19383 12291
rect 19625 12257 19659 12291
rect 15669 12189 15703 12223
rect 15853 12189 15887 12223
rect 17325 12189 17359 12223
rect 12265 12121 12299 12155
rect 11391 12053 11425 12087
rect 11989 12053 12023 12087
rect 12817 12053 12851 12087
rect 14657 12053 14691 12087
rect 14933 12053 14967 12087
rect 15761 12053 15795 12087
rect 17233 12053 17267 12087
rect 18705 12053 18739 12087
rect 11989 11849 12023 11883
rect 12541 11849 12575 11883
rect 13645 11849 13679 11883
rect 16313 11849 16347 11883
rect 17141 11849 17175 11883
rect 17325 11849 17359 11883
rect 17877 11849 17911 11883
rect 20821 11849 20855 11883
rect 10655 11781 10689 11815
rect 13829 11781 13863 11815
rect 14565 11781 14599 11815
rect 17601 11781 17635 11815
rect 11161 11713 11195 11747
rect 10584 11645 10618 11679
rect 10977 11645 11011 11679
rect 11069 11645 11103 11679
rect 11253 11645 11287 11679
rect 11529 11645 11563 11679
rect 11805 11645 11839 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 12633 11645 12667 11679
rect 13369 11645 13403 11679
rect 14289 11645 14323 11679
rect 14933 11645 14967 11679
rect 15189 11645 15223 11679
rect 16405 11645 16439 11679
rect 17417 11645 17451 11679
rect 17509 11645 17543 11679
rect 17693 11645 17727 11679
rect 17785 11645 17819 11679
rect 18245 11645 18279 11679
rect 18521 11645 18555 11679
rect 18705 11645 18739 11679
rect 19165 11645 19199 11679
rect 19432 11645 19466 11679
rect 12357 11577 12391 11611
rect 14105 11577 14139 11611
rect 14381 11577 14415 11611
rect 14565 11577 14599 11611
rect 16957 11577 16991 11611
rect 17173 11577 17207 11611
rect 18153 11577 18187 11611
rect 20729 11577 20763 11611
rect 10885 11509 10919 11543
rect 11437 11509 11471 11543
rect 11713 11509 11747 11543
rect 13277 11509 13311 11543
rect 16497 11509 16531 11543
rect 18429 11509 18463 11543
rect 18797 11509 18831 11543
rect 20545 11509 20579 11543
rect 10655 11305 10689 11339
rect 11253 11305 11287 11339
rect 12449 11305 12483 11339
rect 13829 11305 13863 11339
rect 15393 11305 15427 11339
rect 15669 11305 15703 11339
rect 16221 11305 16255 11339
rect 17049 11305 17083 11339
rect 20361 11305 20395 11339
rect 11897 11237 11931 11271
rect 12265 11237 12299 11271
rect 13553 11237 13587 11271
rect 14280 11237 14314 11271
rect 15577 11237 15611 11271
rect 19248 11237 19282 11271
rect 20545 11237 20579 11271
rect 9505 11169 9539 11203
rect 9597 11169 9631 11203
rect 9965 11169 9999 11203
rect 10241 11169 10275 11203
rect 10517 11169 10551 11203
rect 10758 11169 10792 11203
rect 11069 11169 11103 11203
rect 11253 11167 11287 11201
rect 11437 11169 11471 11203
rect 11529 11169 11563 11203
rect 11621 11169 11655 11203
rect 12633 11169 12667 11203
rect 12909 11169 12943 11203
rect 16497 11169 16531 11203
rect 16681 11169 16715 11203
rect 16957 11169 16991 11203
rect 17489 11169 17523 11203
rect 18889 11169 18923 11203
rect 12817 11101 12851 11135
rect 14013 11101 14047 11135
rect 17233 11101 17267 11135
rect 18981 11101 19015 11135
rect 10149 11033 10183 11067
rect 10425 11033 10459 11067
rect 16773 11033 16807 11067
rect 18797 11033 18831 11067
rect 20821 11033 20855 11067
rect 9873 10965 9907 10999
rect 11713 10965 11747 10999
rect 18613 10965 18647 10999
rect 11161 10761 11195 10795
rect 11713 10761 11747 10795
rect 17509 10761 17543 10795
rect 18245 10761 18279 10795
rect 18889 10761 18923 10795
rect 19625 10761 19659 10795
rect 13829 10693 13863 10727
rect 20177 10693 20211 10727
rect 10517 10625 10551 10659
rect 15393 10625 15427 10659
rect 8861 10557 8895 10591
rect 8953 10557 8987 10591
rect 9229 10557 9263 10591
rect 9321 10557 9355 10591
rect 9413 10557 9447 10591
rect 9781 10557 9815 10591
rect 9873 10557 9907 10591
rect 10333 10557 10367 10591
rect 10609 10557 10643 10591
rect 10885 10557 10919 10591
rect 11805 10557 11839 10591
rect 11897 10557 11931 10591
rect 14197 10557 14231 10591
rect 14473 10557 14507 10591
rect 14933 10557 14967 10591
rect 15209 10557 15243 10591
rect 15485 10557 15519 10591
rect 15761 10557 15795 10591
rect 15853 10557 15887 10591
rect 17877 10557 17911 10591
rect 17969 10557 18003 10591
rect 18153 10557 18187 10591
rect 18797 10557 18831 10591
rect 19257 10557 19291 10591
rect 19533 10557 19567 10591
rect 19809 10557 19843 10591
rect 20085 10557 20119 10591
rect 20545 10557 20579 10591
rect 20637 10557 20671 10591
rect 20913 10557 20947 10591
rect 21005 10557 21039 10591
rect 21189 10557 21223 10591
rect 21465 10557 21499 10591
rect 9965 10489 9999 10523
rect 11069 10489 11103 10523
rect 12142 10489 12176 10523
rect 13645 10489 13679 10523
rect 15669 10489 15703 10523
rect 16120 10489 16154 10523
rect 17417 10489 17451 10523
rect 20453 10489 20487 10523
rect 9137 10421 9171 10455
rect 9689 10421 9723 10455
rect 10241 10421 10275 10455
rect 10793 10421 10827 10455
rect 13277 10421 13311 10455
rect 14289 10421 14323 10455
rect 14565 10421 14599 10455
rect 14841 10421 14875 10455
rect 15117 10421 15151 10455
rect 17233 10421 17267 10455
rect 19349 10421 19383 10455
rect 19901 10421 19935 10455
rect 20729 10421 20763 10455
rect 21281 10421 21315 10455
rect 21557 10421 21591 10455
rect 10793 10217 10827 10251
rect 11345 10217 11379 10251
rect 13737 10217 13771 10251
rect 20637 10217 20671 10251
rect 21649 10217 21683 10251
rect 9658 10149 9692 10183
rect 14013 10149 14047 10183
rect 14749 10149 14783 10183
rect 15301 10149 15335 10183
rect 15853 10149 15887 10183
rect 19524 10149 19558 10183
rect 21373 10149 21407 10183
rect 8769 10081 8803 10115
rect 8861 10081 8895 10115
rect 9321 10081 9355 10115
rect 11069 10081 11103 10115
rect 11713 10081 11747 10115
rect 12173 10081 12207 10115
rect 12265 10081 12299 10115
rect 12357 10081 12391 10115
rect 12541 10081 12575 10115
rect 12817 10081 12851 10115
rect 13093 10081 13127 10115
rect 13436 10081 13470 10115
rect 13645 10081 13679 10115
rect 15761 10081 15795 10115
rect 16773 10081 16807 10115
rect 16957 10081 16991 10115
rect 17141 10081 17175 10115
rect 17417 10081 17451 10115
rect 17693 10081 17727 10115
rect 17960 10081 17994 10115
rect 19257 10081 19291 10115
rect 20729 10081 20763 10115
rect 21833 10081 21867 10115
rect 22109 10081 22143 10115
rect 9413 10013 9447 10047
rect 16313 10013 16347 10047
rect 21925 10013 21959 10047
rect 8953 9945 8987 9979
rect 9229 9945 9263 9979
rect 12081 9945 12115 9979
rect 12633 9945 12667 9979
rect 13185 9945 13219 9979
rect 13507 9945 13541 9979
rect 8677 9877 8711 9911
rect 11805 9877 11839 9911
rect 12909 9877 12943 9911
rect 14105 9877 14139 9911
rect 14841 9877 14875 9911
rect 15577 9877 15611 9911
rect 17049 9877 17083 9911
rect 17325 9877 17359 9911
rect 19073 9877 19107 9911
rect 20821 9877 20855 9911
rect 22201 9877 22235 9911
rect 9505 9673 9539 9707
rect 9965 9673 9999 9707
rect 10885 9673 10919 9707
rect 14473 9673 14507 9707
rect 20545 9673 20579 9707
rect 22017 9673 22051 9707
rect 22293 9673 22327 9707
rect 23397 9673 23431 9707
rect 7849 9605 7883 9639
rect 8677 9605 8711 9639
rect 8953 9605 8987 9639
rect 9229 9605 9263 9639
rect 12081 9605 12115 9639
rect 18797 9605 18831 9639
rect 19533 9605 19567 9639
rect 8125 9537 8159 9571
rect 10333 9537 10367 9571
rect 11437 9537 11471 9571
rect 7757 9469 7791 9503
rect 8217 9469 8251 9503
rect 8585 9469 8619 9503
rect 9021 9479 9055 9513
rect 9137 9479 9171 9513
rect 9597 9469 9631 9503
rect 9873 9469 9907 9503
rect 9971 9469 10005 9503
rect 10149 9469 10183 9503
rect 10425 9469 10459 9503
rect 10517 9469 10551 9503
rect 10977 9469 11011 9503
rect 11253 9469 11287 9503
rect 11345 9469 11379 9503
rect 14156 9469 14190 9503
rect 14381 9469 14415 9503
rect 18889 9469 18923 9503
rect 19257 9469 19291 9503
rect 20821 9469 20855 9503
rect 21097 9469 21131 9503
rect 21465 9469 21499 9503
rect 21557 9469 21591 9503
rect 21649 9469 21683 9503
rect 21925 9469 21959 9503
rect 22385 9469 22419 9503
rect 22477 9469 22511 9503
rect 22937 9469 22971 9503
rect 23029 9469 23063 9503
rect 23121 9469 23155 9503
rect 23305 9469 23339 9503
rect 11161 9401 11195 9435
rect 13369 9401 13403 9435
rect 13645 9401 13679 9435
rect 14013 9401 14047 9435
rect 14243 9401 14277 9435
rect 14841 9401 14875 9435
rect 16773 9401 16807 9435
rect 19717 9401 19751 9435
rect 20085 9401 20119 9435
rect 20637 9401 20671 9435
rect 9781 9333 9815 9367
rect 10609 9333 10643 9367
rect 16129 9333 16163 9367
rect 18061 9333 18095 9367
rect 20913 9333 20947 9367
rect 21189 9333 21223 9367
rect 21741 9333 21775 9367
rect 22569 9333 22603 9367
rect 22845 9333 22879 9367
rect 7941 9129 7975 9163
rect 8125 9129 8159 9163
rect 8953 9129 8987 9163
rect 10609 9129 10643 9163
rect 11805 9129 11839 9163
rect 12081 9129 12115 9163
rect 15485 9129 15519 9163
rect 16681 9129 16715 9163
rect 16957 9129 16991 9163
rect 17233 9129 17267 9163
rect 21925 9129 21959 9163
rect 11069 9061 11103 9095
rect 14013 9061 14047 9095
rect 17417 9061 17451 9095
rect 19165 9061 19199 9095
rect 7389 8993 7423 9027
rect 7665 8993 7699 9027
rect 7757 8993 7791 9027
rect 7941 8993 7975 9027
rect 8217 8993 8251 9027
rect 8493 8993 8527 9027
rect 8585 8993 8619 9027
rect 8861 8993 8895 9027
rect 9229 8993 9263 9027
rect 9496 8993 9530 9027
rect 11897 8993 11931 9027
rect 12173 8993 12207 9027
rect 14197 8993 14231 9027
rect 16405 8993 16439 9027
rect 16589 8993 16623 9027
rect 16865 8993 16899 9027
rect 17325 8993 17359 9027
rect 19524 8993 19558 9027
rect 20729 8993 20763 9027
rect 20913 8993 20947 9027
rect 21373 8993 21407 9027
rect 21833 8993 21867 9027
rect 22109 8993 22143 9027
rect 22385 8983 22419 9017
rect 7573 8925 7607 8959
rect 19257 8925 19291 8959
rect 7297 8857 7331 8891
rect 20637 8857 20671 8891
rect 21649 8857 21683 8891
rect 8401 8789 8435 8823
rect 8677 8789 8711 8823
rect 11161 8789 11195 8823
rect 12541 8789 12575 8823
rect 20821 8789 20855 8823
rect 22201 8789 22235 8823
rect 22477 8789 22511 8823
rect 11253 8585 11287 8619
rect 12725 8585 12759 8619
rect 16727 8585 16761 8619
rect 22109 8585 22143 8619
rect 8125 8517 8159 8551
rect 8769 8517 8803 8551
rect 13277 8517 13311 8551
rect 14933 8517 14967 8551
rect 18797 8517 18831 8551
rect 20545 8517 20579 8551
rect 13553 8449 13587 8483
rect 17601 8449 17635 8483
rect 8217 8381 8251 8415
rect 8585 8381 8619 8415
rect 8677 8381 8711 8415
rect 9137 8381 9171 8415
rect 9321 8381 9355 8415
rect 9689 8381 9723 8415
rect 11345 8381 11379 8415
rect 11621 8381 11655 8415
rect 11713 8381 11747 8415
rect 12265 8381 12299 8415
rect 12541 8381 12575 8415
rect 12633 8381 12667 8415
rect 13093 8375 13127 8409
rect 13185 8381 13219 8415
rect 13809 8381 13843 8415
rect 15117 8381 15151 8415
rect 15853 8381 15887 8415
rect 16037 8381 16071 8415
rect 16129 8381 16163 8415
rect 16565 8381 16599 8415
rect 16798 8389 16832 8423
rect 17141 8381 17175 8415
rect 17325 8381 17359 8415
rect 17417 8381 17451 8415
rect 17693 8375 17727 8409
rect 17785 8381 17819 8415
rect 18705 8381 18739 8415
rect 19165 8381 19199 8415
rect 19432 8381 19466 8415
rect 20729 8381 20763 8415
rect 21373 8381 21407 8415
rect 21465 8381 21499 8415
rect 21741 8381 21775 8415
rect 22017 8381 22051 8415
rect 9045 8313 9079 8347
rect 9873 8313 9907 8347
rect 10241 8313 10275 8347
rect 10609 8313 10643 8347
rect 11529 8313 11563 8347
rect 11805 8313 11839 8347
rect 12173 8313 12207 8347
rect 12449 8313 12483 8347
rect 13001 8313 13035 8347
rect 15485 8313 15519 8347
rect 17877 8313 17911 8347
rect 18061 8313 18095 8347
rect 18429 8313 18463 8347
rect 21281 8313 21315 8347
rect 21557 8313 21591 8347
rect 8493 8245 8527 8279
rect 10701 8245 10735 8279
rect 16497 8245 16531 8279
rect 17049 8245 17083 8279
rect 21005 8245 21039 8279
rect 21833 8245 21867 8279
rect 8401 8041 8435 8075
rect 10609 8041 10643 8075
rect 13001 8041 13035 8075
rect 13645 8041 13679 8075
rect 13829 8041 13863 8075
rect 14979 8041 15013 8075
rect 15669 8041 15703 8075
rect 17417 8041 17451 8075
rect 17693 8041 17727 8075
rect 9474 7973 9508 8007
rect 12265 7973 12299 8007
rect 13277 7973 13311 8007
rect 18521 7973 18555 8007
rect 8493 7905 8527 7939
rect 8769 7905 8803 7939
rect 9045 7905 9079 7939
rect 9229 7905 9263 7939
rect 11161 7905 11195 7939
rect 11621 7905 11655 7939
rect 11989 7905 12023 7939
rect 12081 7905 12115 7939
rect 13093 7905 13127 7939
rect 13369 7905 13403 7939
rect 13461 7905 13495 7939
rect 13645 7905 13679 7939
rect 13921 7905 13955 7939
rect 14197 7905 14231 7939
rect 14381 7905 14415 7939
rect 14841 7905 14875 7939
rect 15050 7911 15084 7945
rect 15209 7905 15243 7939
rect 15485 7905 15519 7939
rect 15669 7905 15703 7939
rect 15761 7905 15795 7939
rect 16497 7905 16531 7939
rect 17141 7905 17175 7939
rect 17509 7905 17543 7939
rect 17785 7905 17819 7939
rect 18061 7905 18095 7939
rect 18972 7905 19006 7939
rect 20269 7905 20303 7939
rect 20729 7905 20763 7939
rect 18705 7837 18739 7871
rect 20821 7837 20855 7871
rect 8677 7769 8711 7803
rect 14473 7769 14507 7803
rect 15853 7769 15887 7803
rect 20085 7769 20119 7803
rect 8953 7701 8987 7735
rect 11253 7701 11287 7735
rect 11713 7701 11747 7735
rect 12357 7701 12391 7735
rect 14105 7701 14139 7735
rect 14749 7701 14783 7735
rect 15301 7701 15335 7735
rect 16405 7701 16439 7735
rect 17049 7701 17083 7735
rect 17969 7701 18003 7735
rect 18429 7701 18463 7735
rect 20545 7701 20579 7735
rect 9689 7497 9723 7531
rect 13277 7497 13311 7531
rect 19901 7497 19935 7531
rect 20177 7497 20211 7531
rect 20453 7497 20487 7531
rect 10241 7429 10275 7463
rect 12081 7429 12115 7463
rect 13829 7429 13863 7463
rect 20729 7429 20763 7463
rect 9413 7361 9447 7395
rect 10701 7361 10735 7395
rect 16957 7361 16991 7395
rect 8953 7293 8987 7327
rect 9321 7293 9355 7327
rect 9781 7293 9815 7327
rect 9965 7293 9999 7327
rect 10057 7293 10091 7327
rect 10333 7293 10367 7327
rect 10425 7293 10459 7327
rect 10517 7293 10551 7327
rect 12541 7293 12575 7327
rect 13185 7293 13219 7327
rect 13921 7293 13955 7327
rect 15209 7293 15243 7327
rect 16681 7293 16715 7327
rect 19257 7293 19291 7327
rect 19717 7293 19751 7327
rect 19993 7293 20027 7327
rect 20269 7303 20303 7337
rect 20361 7293 20395 7327
rect 20637 7293 20671 7327
rect 9045 7225 9079 7259
rect 10946 7225 10980 7259
rect 13001 7225 13035 7259
rect 14105 7225 14139 7259
rect 15025 7225 15059 7259
rect 15476 7225 15510 7259
rect 17202 7225 17236 7259
rect 18797 7225 18831 7259
rect 12449 7157 12483 7191
rect 12909 7157 12943 7191
rect 14197 7157 14231 7191
rect 14933 7157 14967 7191
rect 16589 7157 16623 7191
rect 16773 7157 16807 7191
rect 18337 7157 18371 7191
rect 18889 7157 18923 7191
rect 19349 7157 19383 7191
rect 19625 7157 19659 7191
rect 11897 6953 11931 6987
rect 14657 6953 14691 6987
rect 15485 6953 15519 6987
rect 17233 6953 17267 6987
rect 18705 6953 18739 6987
rect 18981 6953 19015 6987
rect 19257 6953 19291 6987
rect 20361 6953 20395 6987
rect 12265 6885 12299 6919
rect 16681 6885 16715 6919
rect 20085 6885 20119 6919
rect 9781 6817 9815 6851
rect 9873 6817 9907 6851
rect 10057 6817 10091 6851
rect 10149 6817 10183 6851
rect 10517 6817 10551 6851
rect 10793 6817 10827 6851
rect 11161 6817 11195 6851
rect 11437 6817 11471 6851
rect 11621 6817 11655 6851
rect 11897 6817 11931 6851
rect 12081 6817 12115 6851
rect 12173 6817 12207 6851
rect 12633 6817 12667 6851
rect 12900 6817 12934 6851
rect 14473 6817 14507 6851
rect 14565 6817 14599 6851
rect 14841 6817 14875 6851
rect 15025 6817 15059 6851
rect 15301 6817 15335 6851
rect 15393 6817 15427 6851
rect 15669 6817 15703 6851
rect 16313 6817 16347 6851
rect 17325 6817 17359 6851
rect 17417 6817 17451 6851
rect 17877 6817 17911 6851
rect 18061 6817 18095 6851
rect 18521 6817 18555 6851
rect 18613 6817 18647 6851
rect 18889 6817 18923 6851
rect 19349 6817 19383 6851
rect 19441 6817 19475 6851
rect 19717 6817 19751 6851
rect 20177 6817 20211 6851
rect 20269 6817 20303 6851
rect 10425 6749 10459 6783
rect 11345 6749 11379 6783
rect 11713 6681 11747 6715
rect 14013 6681 14047 6715
rect 14381 6681 14415 6715
rect 15761 6681 15795 6715
rect 16865 6681 16899 6715
rect 17509 6681 17543 6715
rect 19809 6681 19843 6715
rect 10701 6613 10735 6647
rect 11069 6613 11103 6647
rect 14933 6613 14967 6647
rect 15209 6613 15243 6647
rect 16405 6613 16439 6647
rect 17969 6613 18003 6647
rect 18429 6613 18463 6647
rect 19533 6613 19567 6647
rect 10793 6409 10827 6443
rect 11345 6409 11379 6443
rect 11621 6409 11655 6443
rect 11897 6409 11931 6443
rect 12173 6409 12207 6443
rect 14657 6409 14691 6443
rect 15577 6409 15611 6443
rect 16865 6409 16899 6443
rect 17417 6409 17451 6443
rect 17785 6409 17819 6443
rect 11069 6341 11103 6375
rect 12725 6341 12759 6375
rect 13001 6341 13035 6375
rect 14289 6341 14323 6375
rect 15301 6341 15335 6375
rect 12449 6273 12483 6307
rect 10701 6205 10735 6239
rect 10977 6205 11011 6239
rect 11161 6205 11195 6239
rect 11437 6205 11471 6239
rect 11713 6205 11747 6239
rect 11989 6205 12023 6239
rect 12265 6205 12299 6239
rect 12357 6205 12391 6239
rect 12633 6205 12667 6239
rect 13093 6205 13127 6239
rect 13185 6205 13219 6239
rect 13645 6205 13679 6239
rect 13921 6205 13955 6239
rect 14381 6205 14415 6239
rect 14565 6205 14599 6239
rect 14933 6205 14967 6239
rect 15025 6205 15059 6239
rect 15209 6205 15243 6239
rect 15669 6205 15703 6239
rect 15761 6205 15795 6239
rect 16497 6205 16531 6239
rect 16957 6205 16991 6239
rect 17049 6205 17083 6239
rect 17141 6205 17175 6239
rect 17325 6205 17359 6239
rect 17693 6205 17727 6239
rect 17877 6205 17911 6239
rect 17969 6205 18003 6239
rect 18245 6205 18279 6239
rect 18429 6205 18463 6239
rect 13277 6137 13311 6171
rect 13737 6137 13771 6171
rect 16405 6137 16439 6171
rect 14013 6069 14047 6103
rect 15853 6069 15887 6103
rect 18061 6069 18095 6103
rect 18245 6069 18279 6103
rect 11897 5865 11931 5899
rect 12541 5865 12575 5899
rect 13553 5865 13587 5899
rect 14105 5865 14139 5899
rect 11897 5729 11931 5763
rect 12081 5729 12115 5763
rect 12173 5729 12207 5763
rect 12265 5729 12299 5763
rect 12449 5729 12483 5763
rect 13093 5729 13127 5763
rect 13185 5729 13219 5763
rect 13277 5729 13311 5763
rect 13461 5729 13495 5763
rect 13921 5729 13955 5763
rect 14105 5729 14139 5763
rect 13001 5525 13035 5559
rect 12357 5321 12391 5355
rect 12633 5321 12667 5355
rect 13001 5321 13035 5355
rect 12449 5117 12483 5151
rect 12541 5117 12575 5151
rect 12909 5117 12943 5151
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 12250 18912 12256 18964
rect 12308 18912 12314 18964
rect 12268 18816 12296 18912
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 12268 18788 12357 18816
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 12526 18572 12532 18624
rect 12584 18572 12590 18624
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 15010 12764 15016 12776
rect 13863 12736 15016 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 15010 12724 15016 12736
rect 15068 12764 15074 12776
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 15068 12736 15485 12764
rect 15068 12724 15074 12736
rect 15473 12733 15485 12736
rect 15519 12764 15531 12767
rect 15519 12736 16344 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 16316 12640 16344 12736
rect 17310 12724 17316 12776
rect 17368 12724 17374 12776
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12764 18935 12767
rect 21266 12764 21272 12776
rect 18923 12736 21272 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 13906 12588 13912 12640
rect 13964 12588 13970 12640
rect 15562 12588 15568 12640
rect 15620 12588 15626 12640
rect 16298 12588 16304 12640
rect 16356 12588 16362 12640
rect 17494 12588 17500 12640
rect 17552 12588 17558 12640
rect 18785 12631 18843 12637
rect 18785 12597 18797 12631
rect 18831 12628 18843 12631
rect 22002 12628 22008 12640
rect 18831 12600 22008 12628
rect 18831 12597 18843 12600
rect 18785 12591 18843 12597
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 12621 12427 12679 12433
rect 12621 12393 12633 12427
rect 12667 12424 12679 12427
rect 13173 12427 13231 12433
rect 12667 12396 13124 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 11482 12291 11540 12297
rect 11482 12257 11494 12291
rect 11528 12288 11540 12291
rect 11655 12291 11713 12297
rect 11655 12288 11667 12291
rect 11528 12260 11667 12288
rect 11528 12257 11540 12260
rect 11482 12251 11540 12257
rect 11655 12257 11667 12260
rect 11701 12257 11713 12291
rect 11655 12251 11713 12257
rect 11758 12290 11816 12296
rect 11758 12256 11770 12290
rect 11804 12256 11816 12290
rect 11758 12250 11816 12256
rect 11773 12220 11801 12250
rect 11882 12248 11888 12300
rect 11940 12248 11946 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12342 12288 12348 12300
rect 12207 12260 12348 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 12434 12248 12440 12300
rect 12492 12248 12498 12300
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 12897 12291 12955 12297
rect 12897 12288 12909 12291
rect 12768 12260 12909 12288
rect 12768 12248 12774 12260
rect 12897 12257 12909 12260
rect 12943 12257 12955 12291
rect 12897 12251 12955 12257
rect 12986 12248 12992 12300
rect 13044 12248 13050 12300
rect 13096 12288 13124 12396
rect 13173 12393 13185 12427
rect 13219 12393 13231 12427
rect 13173 12387 13231 12393
rect 13188 12356 13216 12387
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 16816 12396 17816 12424
rect 16816 12384 16822 12396
rect 17788 12368 17816 12396
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19392 12396 19717 12424
rect 19392 12384 19398 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 19705 12387 19763 12393
rect 13510 12359 13568 12365
rect 13510 12356 13522 12359
rect 13188 12328 13522 12356
rect 13510 12325 13522 12328
rect 13556 12325 13568 12359
rect 13510 12319 13568 12325
rect 15010 12316 15016 12368
rect 15068 12356 15074 12368
rect 17586 12365 17592 12368
rect 17558 12359 17592 12365
rect 15068 12316 15081 12356
rect 17558 12325 17570 12359
rect 17558 12319 17592 12325
rect 17586 12316 17592 12319
rect 17644 12316 17650 12368
rect 17770 12316 17776 12368
rect 17828 12316 17834 12368
rect 18046 12316 18052 12368
rect 18104 12356 18110 12368
rect 18969 12359 19027 12365
rect 18969 12356 18981 12359
rect 18104 12328 18981 12356
rect 18104 12316 18110 12328
rect 18969 12325 18981 12328
rect 19015 12325 19027 12359
rect 18969 12319 19027 12325
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 13096 12260 13277 12288
rect 13265 12257 13277 12260
rect 13311 12288 13323 12291
rect 14826 12288 14832 12300
rect 13311 12260 14832 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 15053 12287 15081 12316
rect 15933 12291 15991 12297
rect 15933 12288 15945 12291
rect 15021 12281 15081 12287
rect 15021 12247 15033 12281
rect 15067 12250 15081 12281
rect 15488 12260 15945 12288
rect 15067 12247 15079 12250
rect 15021 12241 15079 12247
rect 12526 12220 12532 12232
rect 11773 12192 12532 12220
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 8846 12112 8852 12164
rect 8904 12152 8910 12164
rect 12253 12155 12311 12161
rect 12253 12152 12265 12155
rect 8904 12124 12265 12152
rect 8904 12112 8910 12124
rect 12253 12121 12265 12124
rect 12299 12121 12311 12155
rect 15488 12152 15516 12260
rect 15933 12257 15945 12260
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 16758 12248 16764 12300
rect 16816 12248 16822 12300
rect 16853 12291 16911 12297
rect 16853 12257 16865 12291
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 17037 12291 17095 12297
rect 17037 12257 17049 12291
rect 17083 12257 17095 12291
rect 17037 12251 17095 12257
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15620 12192 15669 12220
rect 15620 12180 15626 12192
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12220 15899 12223
rect 16776 12220 16804 12248
rect 15887 12192 16804 12220
rect 15887 12189 15899 12192
rect 15841 12183 15899 12189
rect 16868 12152 16896 12251
rect 12253 12115 12311 12121
rect 14660 12124 16896 12152
rect 17052 12152 17080 12251
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19337 12291 19395 12297
rect 19337 12288 19349 12291
rect 19300 12260 19349 12288
rect 19300 12248 19306 12260
rect 19337 12257 19349 12260
rect 19383 12257 19395 12291
rect 19337 12251 19395 12257
rect 19613 12291 19671 12297
rect 19613 12257 19625 12291
rect 19659 12257 19671 12291
rect 19613 12251 19671 12257
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17313 12223 17371 12229
rect 17313 12220 17325 12223
rect 17184 12192 17325 12220
rect 17184 12180 17190 12192
rect 17313 12189 17325 12192
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 17052 12124 17356 12152
rect 10870 12044 10876 12096
rect 10928 12084 10934 12096
rect 11379 12087 11437 12093
rect 11379 12084 11391 12087
rect 10928 12056 11391 12084
rect 10928 12044 10934 12056
rect 11379 12053 11391 12056
rect 11425 12053 11437 12087
rect 11379 12047 11437 12053
rect 11606 12044 11612 12096
rect 11664 12084 11670 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11664 12056 11989 12084
rect 11664 12044 11670 12056
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 11977 12047 12035 12053
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 12894 12084 12900 12096
rect 12851 12056 12900 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14660 12093 14688 12124
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14424 12056 14657 12084
rect 14424 12044 14430 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 14918 12044 14924 12096
rect 14976 12044 14982 12096
rect 15746 12044 15752 12096
rect 15804 12044 15810 12096
rect 16868 12084 16896 12124
rect 17034 12084 17040 12096
rect 16868 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17218 12044 17224 12096
rect 17276 12044 17282 12096
rect 17328 12084 17356 12124
rect 17678 12084 17684 12096
rect 17328 12056 17684 12084
rect 17678 12044 17684 12056
rect 17736 12084 17742 12096
rect 18693 12087 18751 12093
rect 18693 12084 18705 12087
rect 17736 12056 18705 12084
rect 17736 12044 17742 12056
rect 18693 12053 18705 12056
rect 18739 12084 18751 12087
rect 19426 12084 19432 12096
rect 18739 12056 19432 12084
rect 18739 12053 18751 12056
rect 18693 12047 18751 12053
rect 19426 12044 19432 12056
rect 19484 12084 19490 12096
rect 19628 12084 19656 12251
rect 19484 12056 19656 12084
rect 19484 12044 19490 12056
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9180 11852 11376 11880
rect 9180 11840 9186 11852
rect 10643 11815 10701 11821
rect 10643 11781 10655 11815
rect 10689 11812 10701 11815
rect 11238 11812 11244 11824
rect 10689 11784 11244 11812
rect 10689 11781 10701 11784
rect 10643 11775 10701 11781
rect 11238 11772 11244 11784
rect 11296 11772 11302 11824
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 8720 11716 11161 11744
rect 8720 11704 8726 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11348 11744 11376 11852
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11572 11852 11989 11880
rect 11572 11840 11578 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 11977 11843 12035 11849
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12529 11883 12587 11889
rect 12529 11880 12541 11883
rect 12492 11852 12541 11880
rect 12492 11840 12498 11852
rect 12529 11849 12541 11852
rect 12575 11849 12587 11883
rect 12529 11843 12587 11849
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13044 11852 13645 11880
rect 13044 11840 13050 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 13633 11843 13691 11849
rect 14476 11852 16313 11880
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 12802 11812 12808 11824
rect 11480 11784 12808 11812
rect 11480 11772 11486 11784
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 13817 11815 13875 11821
rect 13817 11781 13829 11815
rect 13863 11812 13875 11815
rect 13906 11812 13912 11824
rect 13863 11784 13912 11812
rect 13863 11781 13875 11784
rect 13817 11775 13875 11781
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 11149 11707 11207 11713
rect 11256 11716 11376 11744
rect 10594 11685 10600 11688
rect 10572 11679 10600 11685
rect 10572 11645 10584 11679
rect 10572 11639 10600 11645
rect 10594 11636 10600 11639
rect 10652 11636 10658 11688
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 11256 11685 11284 11716
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11664 11716 12204 11744
rect 11664 11704 11670 11716
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10744 11648 10977 11676
rect 10744 11636 10750 11648
rect 10965 11645 10977 11648
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11645 11299 11679
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11241 11639 11299 11645
rect 11348 11648 11529 11676
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 11072 11608 11100 11639
rect 11348 11620 11376 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 11974 11676 11980 11688
rect 11839 11648 11980 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12176 11685 12204 11716
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11645 12219 11679
rect 12161 11639 12219 11645
rect 8996 11580 11100 11608
rect 8996 11568 9002 11580
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 12084 11608 12112 11639
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12584 11648 12633 11676
rect 12584 11636 12590 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 13998 11676 14004 11688
rect 13403 11648 14004 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 13998 11636 14004 11648
rect 14056 11636 14062 11688
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11676 14335 11679
rect 14476 11676 14504 11852
rect 16301 11849 16313 11852
rect 16347 11880 16359 11883
rect 16758 11880 16764 11892
rect 16347 11852 16764 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 17129 11883 17187 11889
rect 17129 11849 17141 11883
rect 17175 11880 17187 11883
rect 17218 11880 17224 11892
rect 17175 11852 17224 11880
rect 17175 11849 17187 11852
rect 17129 11843 17187 11849
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 17310 11840 17316 11892
rect 17368 11840 17374 11892
rect 17865 11883 17923 11889
rect 17865 11880 17877 11883
rect 17420 11852 17877 11880
rect 14553 11815 14611 11821
rect 14553 11781 14565 11815
rect 14599 11781 14611 11815
rect 17420 11812 17448 11852
rect 17865 11849 17877 11852
rect 17911 11849 17923 11883
rect 17865 11843 17923 11849
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20680 11852 20821 11880
rect 20680 11840 20686 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 14553 11775 14611 11781
rect 16960 11784 17448 11812
rect 17589 11815 17647 11821
rect 14568 11744 14596 11775
rect 14568 11716 15056 11744
rect 14323 11648 14504 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14884 11648 14933 11676
rect 14884 11636 14890 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 15028 11676 15056 11716
rect 15177 11679 15235 11685
rect 15177 11676 15189 11679
rect 15028 11648 15189 11676
rect 14921 11639 14979 11645
rect 15177 11645 15189 11648
rect 15223 11645 15235 11679
rect 15177 11639 15235 11645
rect 15746 11636 15752 11688
rect 15804 11636 15810 11688
rect 16393 11679 16451 11685
rect 16393 11676 16405 11679
rect 16316 11648 16405 11676
rect 12250 11608 12256 11620
rect 11388 11580 12256 11608
rect 11388 11568 11394 11580
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 12345 11611 12403 11617
rect 12345 11577 12357 11611
rect 12391 11608 12403 11611
rect 12544 11608 12572 11636
rect 12391 11580 12572 11608
rect 12391 11577 12403 11580
rect 12345 11571 12403 11577
rect 13538 11568 13544 11620
rect 13596 11608 13602 11620
rect 14093 11611 14151 11617
rect 14093 11608 14105 11611
rect 13596 11580 14105 11608
rect 13596 11568 13602 11580
rect 14093 11577 14105 11580
rect 14139 11608 14151 11611
rect 14366 11608 14372 11620
rect 14139 11580 14372 11608
rect 14139 11577 14151 11580
rect 14093 11571 14151 11577
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 14553 11611 14611 11617
rect 14553 11577 14565 11611
rect 14599 11608 14611 11611
rect 15764 11608 15792 11636
rect 14599 11580 15792 11608
rect 16316 11608 16344 11648
rect 16393 11645 16405 11648
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 16960 11617 16988 11784
rect 17589 11781 17601 11815
rect 17635 11781 17647 11815
rect 17589 11775 17647 11781
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 17310 11676 17316 11688
rect 17092 11648 17316 11676
rect 17092 11636 17098 11648
rect 17310 11636 17316 11648
rect 17368 11676 17374 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 17368 11648 17417 11676
rect 17368 11636 17374 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 17494 11636 17500 11688
rect 17552 11636 17558 11688
rect 16945 11611 17003 11617
rect 16316 11580 16896 11608
rect 14599 11577 14611 11580
rect 14553 11571 14611 11577
rect 16316 11552 16344 11580
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10192 11512 10885 11540
rect 10192 11500 10198 11512
rect 10873 11509 10885 11512
rect 10919 11509 10931 11543
rect 10873 11503 10931 11509
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 11425 11543 11483 11549
rect 11425 11540 11437 11543
rect 11020 11512 11437 11540
rect 11020 11500 11026 11512
rect 11425 11509 11437 11512
rect 11471 11509 11483 11543
rect 11425 11503 11483 11509
rect 11698 11500 11704 11552
rect 11756 11500 11762 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12710 11540 12716 11552
rect 12492 11512 12716 11540
rect 12492 11500 12498 11512
rect 12710 11500 12716 11512
rect 12768 11540 12774 11552
rect 13265 11543 13323 11549
rect 13265 11540 13277 11543
rect 12768 11512 13277 11540
rect 12768 11500 12774 11512
rect 13265 11509 13277 11512
rect 13311 11509 13323 11543
rect 13265 11503 13323 11509
rect 16298 11500 16304 11552
rect 16356 11500 16362 11552
rect 16482 11500 16488 11552
rect 16540 11500 16546 11552
rect 16868 11540 16896 11580
rect 16945 11577 16957 11611
rect 16991 11577 17003 11611
rect 16945 11571 17003 11577
rect 17161 11611 17219 11617
rect 17161 11577 17173 11611
rect 17207 11608 17219 11611
rect 17604 11608 17632 11775
rect 17678 11772 17684 11824
rect 17736 11772 17742 11824
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 19150 11812 19156 11824
rect 17828 11784 19156 11812
rect 17828 11772 17834 11784
rect 19150 11772 19156 11784
rect 19208 11772 19214 11824
rect 17696 11685 17724 11772
rect 18524 11716 19288 11744
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11645 17739 11679
rect 17681 11639 17739 11645
rect 17773 11679 17831 11685
rect 17773 11645 17785 11679
rect 17819 11645 17831 11679
rect 17773 11639 17831 11645
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18414 11676 18420 11688
rect 18279 11648 18420 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 17788 11608 17816 11639
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 18524 11685 18552 11716
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 17207 11580 17632 11608
rect 17696 11580 17816 11608
rect 17207 11577 17219 11580
rect 17161 11571 17219 11577
rect 17696 11540 17724 11580
rect 17862 11568 17868 11620
rect 17920 11608 17926 11620
rect 18141 11611 18199 11617
rect 18141 11608 18153 11611
rect 17920 11580 18153 11608
rect 17920 11568 17926 11580
rect 18141 11577 18153 11580
rect 18187 11577 18199 11611
rect 18708 11608 18736 11639
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 19116 11648 19165 11676
rect 19116 11636 19122 11648
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 19153 11639 19211 11645
rect 18141 11571 18199 11577
rect 18524 11580 18736 11608
rect 19260 11608 19288 11716
rect 19426 11685 19432 11688
rect 19420 11676 19432 11685
rect 19387 11648 19432 11676
rect 19420 11639 19432 11648
rect 19426 11636 19432 11639
rect 19484 11636 19490 11688
rect 21450 11676 21456 11688
rect 20456 11648 21456 11676
rect 20456 11608 20484 11648
rect 21450 11636 21456 11648
rect 21508 11636 21514 11688
rect 20717 11611 20775 11617
rect 20717 11608 20729 11611
rect 19260 11580 20484 11608
rect 20548 11580 20729 11608
rect 18524 11552 18552 11580
rect 16868 11512 17724 11540
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18417 11543 18475 11549
rect 18417 11540 18429 11543
rect 18104 11512 18429 11540
rect 18104 11500 18110 11512
rect 18417 11509 18429 11512
rect 18463 11509 18475 11543
rect 18417 11503 18475 11509
rect 18506 11500 18512 11552
rect 18564 11500 18570 11552
rect 18785 11543 18843 11549
rect 18785 11509 18797 11543
rect 18831 11540 18843 11543
rect 18874 11540 18880 11552
rect 18831 11512 18880 11540
rect 18831 11509 18843 11512
rect 18785 11503 18843 11509
rect 18874 11500 18880 11512
rect 18932 11500 18938 11552
rect 20548 11549 20576 11580
rect 20717 11577 20729 11580
rect 20763 11577 20775 11611
rect 20717 11571 20775 11577
rect 20533 11543 20591 11549
rect 20533 11509 20545 11543
rect 20579 11509 20591 11543
rect 20533 11503 20591 11509
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 10594 11296 10600 11348
rect 10652 11345 10658 11348
rect 10652 11339 10701 11345
rect 10652 11305 10655 11339
rect 10689 11305 10701 11339
rect 10652 11299 10701 11305
rect 10652 11296 10658 11299
rect 10962 11296 10968 11348
rect 11020 11296 11026 11348
rect 11146 11336 11152 11348
rect 11072 11308 11152 11336
rect 10980 11268 11008 11296
rect 10520 11240 11008 11268
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 8628 11172 9505 11200
rect 8628 11160 8634 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 9582 11160 9588 11212
rect 9640 11160 9646 11212
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 10042 11200 10048 11212
rect 9999 11172 10048 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10520 11209 10548 11240
rect 10229 11203 10287 11209
rect 10229 11169 10241 11203
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 10746 11203 10804 11209
rect 10746 11169 10758 11203
rect 10792 11200 10804 11203
rect 10870 11200 10876 11212
rect 10792 11172 10876 11200
rect 10792 11169 10804 11172
rect 10746 11163 10804 11169
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 10244 11132 10272 11163
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 11072 11209 11100 11308
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 11514 11336 11520 11348
rect 11287 11308 11520 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 11606 11296 11612 11348
rect 11664 11296 11670 11348
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11305 12495 11339
rect 12437 11299 12495 11305
rect 11624 11268 11652 11296
rect 11885 11271 11943 11277
rect 11885 11268 11897 11271
rect 11624 11240 11897 11268
rect 11885 11237 11897 11240
rect 11931 11237 11943 11271
rect 11885 11231 11943 11237
rect 12253 11271 12311 11277
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 12452 11268 12480 11299
rect 12526 11296 12532 11348
rect 12584 11296 12590 11348
rect 13817 11339 13875 11345
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 14182 11336 14188 11348
rect 13863 11308 14188 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14918 11296 14924 11348
rect 14976 11296 14982 11348
rect 15381 11339 15439 11345
rect 15381 11305 15393 11339
rect 15427 11305 15439 11339
rect 15381 11299 15439 11305
rect 12299 11240 12480 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 11238 11160 11244 11212
rect 11296 11198 11302 11212
rect 11296 11170 11339 11198
rect 11296 11160 11302 11170
rect 11422 11160 11428 11212
rect 11480 11160 11486 11212
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 11606 11160 11612 11212
rect 11664 11160 11670 11212
rect 11900 11132 11928 11231
rect 11974 11160 11980 11212
rect 12032 11200 12038 11212
rect 12434 11200 12440 11212
rect 12032 11172 12440 11200
rect 12032 11160 12038 11172
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 12544 11200 12572 11296
rect 13538 11228 13544 11280
rect 13596 11228 13602 11280
rect 14268 11271 14326 11277
rect 14268 11237 14280 11271
rect 14314 11268 14326 11271
rect 14936 11268 14964 11296
rect 14314 11240 14964 11268
rect 15396 11268 15424 11299
rect 15654 11296 15660 11348
rect 15712 11296 15718 11348
rect 16206 11296 16212 11348
rect 16264 11296 16270 11348
rect 16482 11296 16488 11348
rect 16540 11296 16546 11348
rect 17037 11339 17095 11345
rect 17037 11305 17049 11339
rect 17083 11336 17095 11339
rect 18230 11336 18236 11348
rect 17083 11308 18236 11336
rect 17083 11305 17095 11308
rect 17037 11299 17095 11305
rect 18230 11296 18236 11308
rect 18288 11296 18294 11348
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 20395 11308 20576 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 15565 11271 15623 11277
rect 15565 11268 15577 11271
rect 15396 11240 15577 11268
rect 14314 11237 14326 11240
rect 14268 11231 14326 11237
rect 15565 11237 15577 11240
rect 15611 11237 15623 11271
rect 15565 11231 15623 11237
rect 16500 11209 16528 11296
rect 17126 11268 17132 11280
rect 16960 11240 17132 11268
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12544 11172 12633 11200
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 12897 11203 12955 11209
rect 12897 11200 12909 11203
rect 12621 11163 12679 11169
rect 12728 11172 12909 11200
rect 12728 11132 12756 11172
rect 12897 11169 12909 11172
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 16485 11203 16543 11209
rect 16485 11169 16497 11203
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 16850 11200 16856 11212
rect 16715 11172 16856 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 16960 11209 16988 11240
rect 17126 11228 17132 11240
rect 17184 11228 17190 11280
rect 19058 11268 19064 11280
rect 17236 11240 19064 11268
rect 16945 11203 17003 11209
rect 16945 11169 16957 11203
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 9364 11104 11284 11132
rect 11900 11104 12756 11132
rect 9364 11092 9370 11104
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 10137 11067 10195 11073
rect 10137 11064 10149 11067
rect 9088 11036 10149 11064
rect 9088 11024 9094 11036
rect 10137 11033 10149 11036
rect 10183 11033 10195 11067
rect 10137 11027 10195 11033
rect 10413 11067 10471 11073
rect 10413 11033 10425 11067
rect 10459 11064 10471 11067
rect 11146 11064 11152 11076
rect 10459 11036 11152 11064
rect 10459 11033 10471 11036
rect 10413 11027 10471 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 11256 11064 11284 11104
rect 12802 11092 12808 11144
rect 12860 11092 12866 11144
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 14001 11135 14059 11141
rect 14001 11132 14013 11135
rect 13044 11104 14013 11132
rect 13044 11092 13050 11104
rect 14001 11101 14013 11104
rect 14047 11101 14059 11135
rect 14001 11095 14059 11101
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 17236 11141 17264 11240
rect 19058 11228 19064 11240
rect 19116 11228 19122 11280
rect 19242 11277 19248 11280
rect 19236 11268 19248 11277
rect 19203 11240 19248 11268
rect 19236 11231 19248 11240
rect 19242 11228 19248 11231
rect 19300 11228 19306 11280
rect 20548 11277 20576 11308
rect 20533 11271 20591 11277
rect 20533 11237 20545 11271
rect 20579 11237 20591 11271
rect 20533 11231 20591 11237
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 17477 11203 17535 11209
rect 17477 11200 17489 11203
rect 17368 11172 17489 11200
rect 17368 11160 17374 11172
rect 17477 11169 17489 11172
rect 17523 11169 17535 11203
rect 17477 11163 17535 11169
rect 18414 11160 18420 11212
rect 18472 11200 18478 11212
rect 18877 11203 18935 11209
rect 18877 11200 18889 11203
rect 18472 11172 18889 11200
rect 18472 11160 18478 11172
rect 18877 11169 18889 11172
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 16632 11104 17233 11132
rect 16632 11092 16638 11104
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 11974 11064 11980 11076
rect 11256 11036 11980 11064
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 16758 11024 16764 11076
rect 16816 11024 16822 11076
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 18785 11067 18843 11073
rect 18785 11064 18797 11067
rect 18380 11036 18797 11064
rect 18380 11024 18386 11036
rect 18785 11033 18797 11036
rect 18831 11033 18843 11067
rect 18892 11064 18920 11163
rect 18969 11135 19027 11141
rect 18969 11101 18981 11135
rect 19015 11132 19027 11135
rect 19076 11132 19104 11228
rect 19015 11104 19104 11132
rect 19015 11101 19027 11104
rect 18969 11095 19027 11101
rect 20809 11067 20867 11073
rect 18892 11036 19012 11064
rect 18785 11027 18843 11033
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 9861 10999 9919 11005
rect 9861 10996 9873 10999
rect 9732 10968 9873 10996
rect 9732 10956 9738 10968
rect 9861 10965 9873 10968
rect 9907 10965 9919 10999
rect 9861 10959 9919 10965
rect 11698 10956 11704 11008
rect 11756 10956 11762 11008
rect 18598 10956 18604 11008
rect 18656 10956 18662 11008
rect 18984 10996 19012 11036
rect 20809 11033 20821 11067
rect 20855 11064 20867 11067
rect 28258 11064 28264 11076
rect 20855 11036 28264 11064
rect 20855 11033 20867 11036
rect 20809 11027 20867 11033
rect 28258 11024 28264 11036
rect 28316 11024 28322 11076
rect 19334 10996 19340 11008
rect 18984 10968 19340 10996
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 9674 10792 9680 10804
rect 9140 10764 9680 10792
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 8536 10560 8861 10588
rect 8536 10548 8542 10560
rect 8849 10557 8861 10560
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9140 10588 9168 10764
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 10134 10752 10140 10804
rect 10192 10752 10198 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 11112 10764 11161 10792
rect 11112 10752 11118 10764
rect 11149 10761 11161 10764
rect 11195 10761 11207 10795
rect 11149 10755 11207 10761
rect 11698 10752 11704 10804
rect 11756 10752 11762 10804
rect 12894 10792 12900 10804
rect 11808 10764 12900 10792
rect 10152 10724 10180 10752
rect 11422 10724 11428 10736
rect 9324 10696 10180 10724
rect 10336 10696 11428 10724
rect 9324 10656 9352 10696
rect 9232 10628 9352 10656
rect 9784 10628 10180 10656
rect 9232 10597 9260 10628
rect 8987 10560 9168 10588
rect 9217 10591 9275 10597
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10588 9459 10591
rect 9674 10588 9680 10600
rect 9447 10560 9680 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9784 10597 9812 10628
rect 10152 10600 10180 10628
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 9324 10520 9352 10548
rect 9876 10520 9904 10551
rect 10134 10548 10140 10600
rect 10192 10548 10198 10600
rect 10336 10597 10364 10696
rect 11422 10684 11428 10696
rect 11480 10684 11486 10736
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 10551 10628 11376 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 8812 10492 9352 10520
rect 9416 10492 9904 10520
rect 9953 10523 10011 10529
rect 8812 10480 8818 10492
rect 9416 10464 9444 10492
rect 9953 10489 9965 10523
rect 9999 10520 10011 10523
rect 10612 10520 10640 10551
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 9999 10492 10364 10520
rect 10612 10492 11008 10520
rect 9999 10489 10011 10492
rect 9953 10483 10011 10489
rect 10336 10464 10364 10492
rect 7834 10412 7840 10464
rect 7892 10452 7898 10464
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 7892 10424 9137 10452
rect 7892 10412 7898 10424
rect 9125 10421 9137 10424
rect 9171 10421 9183 10455
rect 9125 10415 9183 10421
rect 9398 10412 9404 10464
rect 9456 10412 9462 10464
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9858 10452 9864 10464
rect 9723 10424 9864 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10226 10412 10232 10464
rect 10284 10412 10290 10464
rect 10318 10412 10324 10464
rect 10376 10412 10382 10464
rect 10778 10412 10784 10464
rect 10836 10412 10842 10464
rect 10980 10452 11008 10492
rect 11054 10480 11060 10532
rect 11112 10480 11118 10532
rect 11348 10520 11376 10628
rect 11808 10597 11836 10764
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 15856 10764 16804 10792
rect 13814 10684 13820 10736
rect 13872 10684 13878 10736
rect 12986 10616 12992 10668
rect 13044 10616 13050 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 14936 10628 15393 10656
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10588 11943 10591
rect 12526 10588 12532 10600
rect 11931 10560 12532 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 12526 10548 12532 10560
rect 12584 10588 12590 10600
rect 13004 10588 13032 10616
rect 12584 10560 13032 10588
rect 12584 10548 12590 10560
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 14056 10560 14197 10588
rect 14056 10548 14062 10560
rect 14185 10557 14197 10560
rect 14231 10588 14243 10591
rect 14366 10588 14372 10600
rect 14231 10560 14372 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14936 10597 14964 10628
rect 15381 10625 15393 10628
rect 15427 10625 15439 10659
rect 15856 10656 15884 10764
rect 16776 10724 16804 10764
rect 17494 10752 17500 10804
rect 17552 10752 17558 10804
rect 18230 10752 18236 10804
rect 18288 10752 18294 10804
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 18877 10795 18935 10801
rect 18877 10792 18889 10795
rect 18748 10764 18889 10792
rect 18748 10752 18754 10764
rect 18877 10761 18889 10764
rect 18923 10761 18935 10795
rect 18877 10755 18935 10761
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10792 19671 10795
rect 20714 10792 20720 10804
rect 19659 10764 20720 10792
rect 19659 10761 19671 10764
rect 19613 10755 19671 10761
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 18506 10724 18512 10736
rect 16776 10696 18512 10724
rect 18506 10684 18512 10696
rect 18564 10724 18570 10736
rect 20165 10727 20223 10733
rect 18564 10696 20116 10724
rect 18564 10684 18570 10696
rect 15381 10619 15439 10625
rect 15764 10628 15884 10656
rect 15764 10597 15792 10628
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19392 10628 19564 10656
rect 19392 10616 19398 10628
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10557 14979 10591
rect 14921 10551 14979 10557
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10588 15531 10591
rect 15749 10591 15807 10597
rect 15749 10588 15761 10591
rect 15519 10560 15761 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 15749 10557 15761 10560
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 15841 10591 15899 10597
rect 15841 10557 15853 10591
rect 15887 10588 15899 10591
rect 16574 10588 16580 10600
rect 15887 10560 16580 10588
rect 15887 10557 15899 10560
rect 15841 10551 15899 10557
rect 12130 10523 12188 10529
rect 12130 10520 12142 10523
rect 11348 10492 12142 10520
rect 12130 10489 12142 10492
rect 12176 10489 12188 10523
rect 12130 10483 12188 10489
rect 13633 10523 13691 10529
rect 13633 10489 13645 10523
rect 13679 10489 13691 10523
rect 13633 10483 13691 10489
rect 11514 10452 11520 10464
rect 10980 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 13265 10455 13323 10461
rect 13265 10421 13277 10455
rect 13311 10452 13323 10455
rect 13648 10452 13676 10483
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 14476 10520 14504 10551
rect 13780 10492 14504 10520
rect 15212 10520 15240 10551
rect 16574 10548 16580 10560
rect 16632 10548 16638 10600
rect 17862 10548 17868 10600
rect 17920 10548 17926 10600
rect 17957 10591 18015 10597
rect 17957 10557 17969 10591
rect 18003 10588 18015 10591
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 18003 10560 18153 10588
rect 18003 10557 18015 10560
rect 17957 10551 18015 10557
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18656 10560 18797 10588
rect 18656 10548 18662 10560
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 18785 10551 18843 10557
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 19536 10597 19564 10628
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 18932 10560 19257 10588
rect 18932 10548 18938 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 19978 10588 19984 10600
rect 19843 10560 19984 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 15657 10523 15715 10529
rect 15657 10520 15669 10523
rect 15212 10492 15669 10520
rect 13780 10480 13786 10492
rect 15657 10489 15669 10492
rect 15703 10489 15715 10523
rect 15657 10483 15715 10489
rect 16108 10523 16166 10529
rect 16108 10489 16120 10523
rect 16154 10520 16166 10523
rect 16206 10520 16212 10532
rect 16154 10492 16212 10520
rect 16154 10489 16166 10492
rect 16108 10483 16166 10489
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 17405 10523 17463 10529
rect 17405 10489 17417 10523
rect 17451 10489 17463 10523
rect 19536 10520 19564 10551
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20088 10597 20116 10696
rect 20165 10693 20177 10727
rect 20211 10724 20223 10727
rect 21726 10724 21732 10736
rect 20211 10696 21732 10724
rect 20211 10693 20223 10696
rect 20165 10687 20223 10693
rect 21726 10684 21732 10696
rect 21784 10684 21790 10736
rect 20456 10628 20668 10656
rect 20073 10591 20131 10597
rect 20073 10557 20085 10591
rect 20119 10557 20131 10591
rect 20073 10551 20131 10557
rect 20456 10529 20484 10628
rect 20640 10597 20668 10628
rect 20916 10628 21496 10656
rect 20916 10597 20944 10628
rect 21468 10597 21496 10628
rect 20533 10591 20591 10597
rect 20533 10557 20545 10591
rect 20579 10557 20591 10591
rect 20533 10551 20591 10557
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10588 20683 10591
rect 20901 10591 20959 10597
rect 20901 10588 20913 10591
rect 20671 10560 20913 10588
rect 20671 10557 20683 10560
rect 20625 10551 20683 10557
rect 20901 10557 20913 10560
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10588 21051 10591
rect 21177 10591 21235 10597
rect 21177 10588 21189 10591
rect 21039 10560 21189 10588
rect 21039 10557 21051 10560
rect 20993 10551 21051 10557
rect 21177 10557 21189 10560
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21453 10591 21511 10597
rect 21453 10557 21465 10591
rect 21499 10588 21511 10591
rect 21634 10588 21640 10600
rect 21499 10560 21640 10588
rect 21499 10557 21511 10560
rect 21453 10551 21511 10557
rect 20441 10523 20499 10529
rect 20441 10520 20453 10523
rect 19536 10492 20453 10520
rect 17405 10483 17463 10489
rect 20441 10489 20453 10492
rect 20487 10489 20499 10523
rect 20548 10520 20576 10551
rect 21634 10548 21640 10560
rect 21692 10548 21698 10600
rect 22278 10520 22284 10532
rect 20548 10492 22284 10520
rect 20441 10483 20499 10489
rect 13311 10424 13676 10452
rect 13311 10421 13323 10424
rect 13265 10415 13323 10421
rect 14274 10412 14280 10464
rect 14332 10412 14338 10464
rect 14550 10412 14556 10464
rect 14608 10412 14614 10464
rect 14826 10412 14832 10464
rect 14884 10412 14890 10464
rect 15102 10412 15108 10464
rect 15160 10412 15166 10464
rect 17221 10455 17279 10461
rect 17221 10421 17233 10455
rect 17267 10452 17279 10455
rect 17420 10452 17448 10483
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 17267 10424 17448 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 18966 10412 18972 10464
rect 19024 10452 19030 10464
rect 19337 10455 19395 10461
rect 19337 10452 19349 10455
rect 19024 10424 19349 10452
rect 19024 10412 19030 10424
rect 19337 10421 19349 10424
rect 19383 10421 19395 10455
rect 19337 10415 19395 10421
rect 19886 10412 19892 10464
rect 19944 10412 19950 10464
rect 20717 10455 20775 10461
rect 20717 10421 20729 10455
rect 20763 10452 20775 10455
rect 21174 10452 21180 10464
rect 20763 10424 21180 10452
rect 20763 10421 20775 10424
rect 20717 10415 20775 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 21542 10412 21548 10464
rect 21600 10412 21606 10464
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 10226 10248 10232 10260
rect 8168 10220 10232 10248
rect 8168 10208 8174 10220
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10781 10251 10839 10257
rect 10781 10217 10793 10251
rect 10827 10248 10839 10251
rect 11054 10248 11060 10260
rect 10827 10220 11060 10248
rect 10827 10217 10839 10220
rect 10781 10211 10839 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11330 10208 11336 10260
rect 11388 10208 11394 10260
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12216 10220 13676 10248
rect 12216 10208 12222 10220
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 9646 10183 9704 10189
rect 9646 10180 9658 10183
rect 8536 10152 9658 10180
rect 8536 10140 8542 10152
rect 9646 10149 9658 10152
rect 9692 10149 9704 10183
rect 9646 10143 9704 10149
rect 10318 10140 10324 10192
rect 10376 10140 10382 10192
rect 10870 10140 10876 10192
rect 10928 10140 10934 10192
rect 11146 10140 11152 10192
rect 11204 10140 11210 10192
rect 12360 10152 13124 10180
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8757 10115 8815 10121
rect 8757 10112 8769 10115
rect 8444 10084 8769 10112
rect 8444 10072 8450 10084
rect 8757 10081 8769 10084
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 8849 10115 8907 10121
rect 8849 10081 8861 10115
rect 8895 10112 8907 10115
rect 9214 10112 9220 10124
rect 8895 10084 9220 10112
rect 8895 10081 8907 10084
rect 8849 10075 8907 10081
rect 9214 10072 9220 10084
rect 9272 10112 9278 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 9272 10084 9321 10112
rect 9272 10072 9278 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 10336 10112 10364 10140
rect 9548 10084 10364 10112
rect 9548 10072 9554 10084
rect 9401 10047 9459 10053
rect 9401 10044 9413 10047
rect 8864 10016 9260 10044
rect 8202 9936 8208 9988
rect 8260 9976 8266 9988
rect 8864 9976 8892 10016
rect 9232 9985 9260 10016
rect 9324 10016 9413 10044
rect 9324 9988 9352 10016
rect 9401 10013 9413 10016
rect 9447 10013 9459 10047
rect 10888 10044 10916 10140
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11164 10112 11192 10140
rect 11103 10084 11192 10112
rect 11701 10115 11759 10121
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11701 10081 11713 10115
rect 11747 10112 11759 10115
rect 11790 10112 11796 10124
rect 11747 10084 11796 10112
rect 11747 10081 11759 10084
rect 11701 10075 11759 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 12158 10072 12164 10124
rect 12216 10072 12222 10124
rect 12250 10072 12256 10124
rect 12308 10072 12314 10124
rect 12360 10121 12388 10152
rect 13096 10121 13124 10152
rect 13648 10121 13676 10220
rect 13722 10208 13728 10260
rect 13780 10208 13786 10260
rect 14274 10208 14280 10260
rect 14332 10208 14338 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14884 10220 15332 10248
rect 14884 10208 14890 10220
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 14001 10183 14059 10189
rect 14001 10180 14013 10183
rect 13872 10152 14013 10180
rect 13872 10140 13878 10152
rect 14001 10149 14013 10152
rect 14047 10149 14059 10183
rect 14292 10180 14320 10208
rect 14737 10183 14795 10189
rect 14737 10180 14749 10183
rect 14292 10152 14749 10180
rect 14001 10143 14059 10149
rect 14737 10149 14749 10152
rect 14783 10149 14795 10183
rect 14737 10143 14795 10149
rect 15102 10140 15108 10192
rect 15160 10140 15166 10192
rect 15304 10189 15332 10220
rect 16206 10208 16212 10260
rect 16264 10208 16270 10260
rect 17034 10248 17040 10260
rect 16868 10220 17040 10248
rect 15289 10183 15347 10189
rect 15289 10149 15301 10183
rect 15335 10149 15347 10183
rect 15289 10143 15347 10149
rect 15841 10183 15899 10189
rect 15841 10149 15853 10183
rect 15887 10180 15899 10183
rect 16224 10180 16252 10208
rect 15887 10152 16252 10180
rect 15887 10149 15899 10152
rect 15841 10143 15899 10149
rect 12345 10115 12403 10121
rect 12345 10081 12357 10115
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 12529 10115 12587 10121
rect 12529 10081 12541 10115
rect 12575 10112 12587 10115
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12575 10084 12817 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 13424 10115 13482 10121
rect 13424 10081 13436 10115
rect 13470 10112 13482 10115
rect 13633 10115 13691 10121
rect 13470 10084 13584 10112
rect 13470 10081 13482 10084
rect 13424 10075 13482 10081
rect 12268 10044 12296 10072
rect 10888 10016 12296 10044
rect 9401 10007 9459 10013
rect 8260 9948 8892 9976
rect 8941 9979 8999 9985
rect 8260 9936 8266 9948
rect 8941 9945 8953 9979
rect 8987 9976 8999 9979
rect 9217 9979 9275 9985
rect 8987 9948 9168 9976
rect 8987 9945 8999 9948
rect 8941 9939 8999 9945
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 7984 9880 8677 9908
rect 7984 9868 7990 9880
rect 8665 9877 8677 9880
rect 8711 9877 8723 9911
rect 9140 9908 9168 9948
rect 9217 9945 9229 9979
rect 9263 9945 9275 9979
rect 9217 9939 9275 9945
rect 9306 9936 9312 9988
rect 9364 9936 9370 9988
rect 11514 9936 11520 9988
rect 11572 9976 11578 9988
rect 12069 9979 12127 9985
rect 12069 9976 12081 9979
rect 11572 9948 12081 9976
rect 11572 9936 11578 9948
rect 12069 9945 12081 9948
rect 12115 9976 12127 9979
rect 12342 9976 12348 9988
rect 12115 9948 12348 9976
rect 12115 9945 12127 9948
rect 12069 9939 12127 9945
rect 12342 9936 12348 9948
rect 12400 9976 12406 9988
rect 12544 9976 12572 10075
rect 13556 10044 13584 10084
rect 13633 10081 13645 10115
rect 13679 10112 13691 10115
rect 14090 10112 14096 10124
rect 13679 10084 14096 10112
rect 13679 10081 13691 10084
rect 13633 10075 13691 10081
rect 14090 10072 14096 10084
rect 14148 10112 14154 10124
rect 15120 10112 15148 10140
rect 14148 10084 15148 10112
rect 15749 10115 15807 10121
rect 14148 10072 14154 10084
rect 15749 10081 15761 10115
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 16761 10115 16819 10121
rect 16761 10081 16773 10115
rect 16807 10112 16819 10115
rect 16868 10112 16896 10220
rect 17034 10208 17040 10220
rect 17092 10248 17098 10260
rect 17862 10248 17868 10260
rect 17092 10220 17868 10248
rect 17092 10208 17098 10220
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 20625 10251 20683 10257
rect 20625 10217 20637 10251
rect 20671 10248 20683 10251
rect 20671 10220 21404 10248
rect 20671 10217 20683 10220
rect 20625 10211 20683 10217
rect 19512 10183 19570 10189
rect 17696 10152 19288 10180
rect 17696 10124 17724 10152
rect 16807 10084 16896 10112
rect 16807 10081 16819 10084
rect 16761 10075 16819 10081
rect 14182 10044 14188 10056
rect 13556 10016 14188 10044
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14366 10004 14372 10056
rect 14424 10044 14430 10056
rect 14734 10044 14740 10056
rect 14424 10016 14740 10044
rect 14424 10004 14430 10016
rect 14734 10004 14740 10016
rect 14792 10044 14798 10056
rect 15764 10044 15792 10075
rect 16942 10072 16948 10124
rect 17000 10072 17006 10124
rect 17126 10072 17132 10124
rect 17184 10072 17190 10124
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 14792 10016 15792 10044
rect 14792 10004 14798 10016
rect 12400 9948 12572 9976
rect 12621 9979 12679 9985
rect 12400 9936 12406 9948
rect 12621 9945 12633 9979
rect 12667 9976 12679 9979
rect 13173 9979 13231 9985
rect 13173 9976 13185 9979
rect 12667 9948 13185 9976
rect 12667 9945 12679 9948
rect 12621 9939 12679 9945
rect 13173 9945 13185 9948
rect 13219 9945 13231 9979
rect 13173 9939 13231 9945
rect 13495 9979 13553 9985
rect 13495 9945 13507 9979
rect 13541 9976 13553 9979
rect 15194 9976 15200 9988
rect 13541 9948 15200 9976
rect 13541 9945 13553 9948
rect 13495 9939 13553 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 15764 9976 15792 10016
rect 16298 10004 16304 10056
rect 16356 10004 16362 10056
rect 17218 9976 17224 9988
rect 15764 9948 17224 9976
rect 17218 9936 17224 9948
rect 17276 9936 17282 9988
rect 9766 9908 9772 9920
rect 9140 9880 9772 9908
rect 8665 9871 8723 9877
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 11330 9908 11336 9920
rect 10192 9880 11336 9908
rect 10192 9868 10198 9880
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 11793 9911 11851 9917
rect 11793 9877 11805 9911
rect 11839 9908 11851 9911
rect 12710 9908 12716 9920
rect 11839 9880 12716 9908
rect 11839 9877 11851 9880
rect 11793 9871 11851 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 12897 9911 12955 9917
rect 12897 9877 12909 9911
rect 12943 9908 12955 9911
rect 13814 9908 13820 9920
rect 12943 9880 13820 9908
rect 12943 9877 12955 9880
rect 12897 9871 12955 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 14056 9880 14105 9908
rect 14056 9868 14062 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 14826 9868 14832 9920
rect 14884 9868 14890 9920
rect 15565 9911 15623 9917
rect 15565 9877 15577 9911
rect 15611 9908 15623 9911
rect 16482 9908 16488 9920
rect 15611 9880 16488 9908
rect 15611 9877 15623 9880
rect 15565 9871 15623 9877
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17037 9911 17095 9917
rect 17037 9908 17049 9911
rect 16724 9880 17049 9908
rect 16724 9868 16730 9880
rect 17037 9877 17049 9880
rect 17083 9877 17095 9911
rect 17037 9871 17095 9877
rect 17310 9868 17316 9920
rect 17368 9868 17374 9920
rect 17420 9908 17448 10075
rect 17678 10072 17684 10124
rect 17736 10072 17742 10124
rect 17948 10115 18006 10121
rect 17948 10081 17960 10115
rect 17994 10112 18006 10115
rect 18966 10112 18972 10124
rect 17994 10084 18972 10112
rect 17994 10081 18006 10084
rect 17948 10075 18006 10081
rect 18966 10072 18972 10084
rect 19024 10072 19030 10124
rect 19260 10121 19288 10152
rect 19512 10149 19524 10183
rect 19558 10180 19570 10183
rect 21266 10180 21272 10192
rect 19558 10152 21272 10180
rect 19558 10149 19570 10152
rect 19512 10143 19570 10149
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 21376 10189 21404 10220
rect 21542 10208 21548 10260
rect 21600 10208 21606 10260
rect 21637 10251 21695 10257
rect 21637 10217 21649 10251
rect 21683 10248 21695 10251
rect 31662 10248 31668 10260
rect 21683 10220 31668 10248
rect 21683 10217 21695 10220
rect 21637 10211 21695 10217
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 21361 10183 21419 10189
rect 21361 10149 21373 10183
rect 21407 10149 21419 10183
rect 21560 10180 21588 10208
rect 21560 10152 22140 10180
rect 21361 10143 21419 10149
rect 19245 10115 19303 10121
rect 19245 10081 19257 10115
rect 19291 10081 19303 10115
rect 19245 10075 19303 10081
rect 19886 10072 19892 10124
rect 19944 10112 19950 10124
rect 22112 10121 22140 10152
rect 20717 10115 20775 10121
rect 20717 10112 20729 10115
rect 19944 10084 20729 10112
rect 19944 10072 19950 10084
rect 20717 10081 20729 10084
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 21821 10115 21879 10121
rect 21821 10081 21833 10115
rect 21867 10081 21879 10115
rect 21821 10075 21879 10081
rect 22097 10115 22155 10121
rect 22097 10081 22109 10115
rect 22143 10081 22155 10115
rect 22097 10075 22155 10081
rect 18616 9948 19196 9976
rect 18414 9908 18420 9920
rect 17420 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9908 18478 9920
rect 18616 9908 18644 9948
rect 18472 9880 18644 9908
rect 18472 9868 18478 9880
rect 19058 9868 19064 9920
rect 19116 9868 19122 9920
rect 19168 9908 19196 9948
rect 20254 9936 20260 9988
rect 20312 9976 20318 9988
rect 21542 9976 21548 9988
rect 20312 9948 21548 9976
rect 20312 9936 20318 9948
rect 21542 9936 21548 9948
rect 21600 9976 21606 9988
rect 21836 9976 21864 10075
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 22186 10044 22192 10056
rect 21959 10016 22192 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 22186 10004 22192 10016
rect 22244 10004 22250 10056
rect 22554 9976 22560 9988
rect 21600 9948 22560 9976
rect 21600 9936 21606 9948
rect 22554 9936 22560 9948
rect 22612 9936 22618 9988
rect 20809 9911 20867 9917
rect 20809 9908 20821 9911
rect 19168 9880 20821 9908
rect 20809 9877 20821 9880
rect 20855 9877 20867 9911
rect 20809 9871 20867 9877
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22189 9911 22247 9917
rect 22189 9908 22201 9911
rect 22060 9880 22201 9908
rect 22060 9868 22066 9880
rect 22189 9877 22201 9880
rect 22235 9877 22247 9911
rect 22189 9871 22247 9877
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 9398 9664 9404 9716
rect 9456 9664 9462 9716
rect 9490 9664 9496 9716
rect 9548 9664 9554 9716
rect 9953 9707 10011 9713
rect 9953 9673 9965 9707
rect 9999 9704 10011 9707
rect 10778 9704 10784 9716
rect 9999 9676 10784 9704
rect 9999 9673 10011 9676
rect 9953 9667 10011 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 10873 9707 10931 9713
rect 10873 9673 10885 9707
rect 10919 9704 10931 9707
rect 13630 9704 13636 9716
rect 10919 9676 13636 9704
rect 10919 9673 10931 9676
rect 10873 9667 10931 9673
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 14461 9707 14519 9713
rect 14461 9673 14473 9707
rect 14507 9704 14519 9707
rect 14550 9704 14556 9716
rect 14507 9676 14556 9704
rect 14507 9673 14519 9676
rect 14461 9667 14519 9673
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 20533 9707 20591 9713
rect 20533 9673 20545 9707
rect 20579 9704 20591 9707
rect 22005 9707 22063 9713
rect 20579 9676 21956 9704
rect 20579 9673 20591 9676
rect 20533 9667 20591 9673
rect 7837 9639 7895 9645
rect 7837 9605 7849 9639
rect 7883 9636 7895 9639
rect 8570 9636 8576 9648
rect 7883 9608 8576 9636
rect 7883 9605 7895 9608
rect 7837 9599 7895 9605
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 8662 9596 8668 9648
rect 8720 9596 8726 9648
rect 8941 9639 8999 9645
rect 8941 9605 8953 9639
rect 8987 9636 8999 9639
rect 9122 9636 9128 9648
rect 8987 9608 9128 9636
rect 8987 9605 8999 9608
rect 8941 9599 8999 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 9217 9639 9275 9645
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 9416 9636 9444 9664
rect 10134 9636 10140 9648
rect 9263 9608 9444 9636
rect 9784 9608 10140 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 9009 9513 9067 9519
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7392 9472 7757 9500
rect 7392 9376 7420 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 8202 9460 8208 9512
rect 8260 9460 8266 9512
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 8588 9432 8616 9463
rect 8846 9460 8852 9512
rect 8904 9500 8910 9512
rect 9009 9500 9021 9513
rect 8904 9479 9021 9500
rect 9055 9510 9067 9513
rect 9125 9513 9183 9519
rect 9055 9479 9076 9510
rect 8904 9472 9076 9479
rect 9125 9479 9137 9513
rect 9171 9500 9183 9513
rect 9585 9503 9643 9509
rect 9171 9479 9536 9500
rect 9125 9473 9536 9479
rect 9140 9472 9536 9473
rect 8904 9460 8910 9472
rect 9140 9432 9168 9472
rect 8588 9404 9168 9432
rect 9508 9376 9536 9472
rect 9585 9469 9597 9503
rect 9631 9469 9643 9503
rect 9784 9500 9812 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 12069 9639 12127 9645
rect 12069 9605 12081 9639
rect 12115 9636 12127 9639
rect 12526 9636 12532 9648
rect 12115 9608 12532 9636
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 16298 9636 16304 9648
rect 13964 9608 16304 9636
rect 13964 9596 13970 9608
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 10284 9540 10333 9568
rect 10284 9528 10290 9540
rect 10321 9537 10333 9540
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 11425 9571 11483 9577
rect 11425 9537 11437 9571
rect 11471 9568 11483 9571
rect 11606 9568 11612 9580
rect 11471 9540 11612 9568
rect 11471 9537 11483 9540
rect 11425 9531 11483 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 14274 9528 14280 9580
rect 14332 9528 14338 9580
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9784 9472 9873 9500
rect 9585 9463 9643 9469
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9600 9432 9628 9463
rect 9950 9460 9956 9512
rect 10008 9509 10014 9512
rect 10008 9500 10017 9509
rect 10008 9472 10053 9500
rect 10008 9463 10017 9472
rect 10008 9460 10014 9463
rect 10134 9460 10140 9512
rect 10192 9460 10198 9512
rect 10410 9460 10416 9512
rect 10468 9460 10474 9512
rect 10502 9460 10508 9512
rect 10560 9460 10566 9512
rect 10962 9460 10968 9512
rect 11020 9460 11026 9512
rect 11238 9460 11244 9512
rect 11296 9460 11302 9512
rect 11330 9460 11336 9512
rect 11388 9460 11394 9512
rect 14144 9503 14202 9509
rect 14144 9469 14156 9503
rect 14190 9500 14202 9503
rect 14292 9500 14320 9528
rect 14384 9509 14412 9608
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 17218 9596 17224 9648
rect 17276 9636 17282 9648
rect 18785 9639 18843 9645
rect 18785 9636 18797 9639
rect 17276 9608 18797 9636
rect 17276 9596 17282 9608
rect 18785 9605 18797 9608
rect 18831 9605 18843 9639
rect 18785 9599 18843 9605
rect 19518 9596 19524 9648
rect 19576 9596 19582 9648
rect 21928 9636 21956 9676
rect 22005 9673 22017 9707
rect 22051 9704 22063 9707
rect 22094 9704 22100 9716
rect 22051 9676 22100 9704
rect 22051 9673 22063 9676
rect 22005 9667 22063 9673
rect 22094 9664 22100 9676
rect 22152 9664 22158 9716
rect 22278 9664 22284 9716
rect 22336 9664 22342 9716
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 23385 9707 23443 9713
rect 23385 9704 23397 9707
rect 22428 9676 23397 9704
rect 22428 9664 22434 9676
rect 23385 9673 23397 9676
rect 23431 9673 23443 9707
rect 23385 9667 23443 9673
rect 28258 9636 28264 9648
rect 21928 9608 28264 9636
rect 28258 9596 28264 9608
rect 28316 9596 28322 9648
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22244 9540 22508 9568
rect 22244 9528 22250 9540
rect 14190 9472 14320 9500
rect 14369 9503 14427 9509
rect 14190 9469 14202 9472
rect 14144 9463 14202 9469
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 14369 9463 14427 9469
rect 18524 9472 18889 9500
rect 10226 9432 10232 9444
rect 9600 9404 10232 9432
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 10928 9404 11161 9432
rect 10928 9392 10934 9404
rect 11149 9401 11161 9404
rect 11195 9401 11207 9435
rect 11348 9432 11376 9460
rect 18524 9444 18552 9472
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 19116 9472 19257 9500
rect 19116 9460 19122 9472
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 20809 9503 20867 9509
rect 20809 9500 20821 9503
rect 20772 9472 20821 9500
rect 20772 9460 20778 9472
rect 20809 9469 20821 9472
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 21082 9460 21088 9512
rect 21140 9460 21146 9512
rect 21450 9460 21456 9512
rect 21508 9460 21514 9512
rect 21542 9460 21548 9512
rect 21600 9460 21606 9512
rect 21634 9460 21640 9512
rect 21692 9460 21698 9512
rect 21726 9460 21732 9512
rect 21784 9500 21790 9512
rect 21913 9503 21971 9509
rect 21913 9500 21925 9503
rect 21784 9472 21925 9500
rect 21784 9460 21790 9472
rect 21913 9469 21925 9472
rect 21959 9469 21971 9503
rect 21913 9463 21971 9469
rect 22002 9460 22008 9512
rect 22060 9460 22066 9512
rect 22370 9460 22376 9512
rect 22428 9460 22434 9512
rect 22480 9509 22508 9540
rect 22554 9528 22560 9580
rect 22612 9568 22618 9580
rect 22612 9540 22968 9568
rect 22612 9528 22618 9540
rect 22940 9509 22968 9540
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9469 22523 9503
rect 22465 9463 22523 9469
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23017 9503 23075 9509
rect 23017 9500 23029 9503
rect 22971 9472 23029 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23017 9469 23029 9472
rect 23063 9469 23075 9503
rect 23017 9463 23075 9469
rect 23109 9503 23167 9509
rect 23109 9469 23121 9503
rect 23155 9500 23167 9503
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 23155 9472 23305 9500
rect 23155 9469 23167 9472
rect 23109 9463 23167 9469
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 12066 9432 12072 9444
rect 11348 9404 12072 9432
rect 11149 9395 11207 9401
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 13354 9392 13360 9444
rect 13412 9392 13418 9444
rect 13446 9392 13452 9444
rect 13504 9432 13510 9444
rect 13633 9435 13691 9441
rect 13633 9432 13645 9435
rect 13504 9404 13645 9432
rect 13504 9392 13510 9404
rect 13633 9401 13645 9404
rect 13679 9401 13691 9435
rect 13633 9395 13691 9401
rect 13998 9392 14004 9444
rect 14056 9392 14062 9444
rect 14231 9435 14289 9441
rect 14231 9401 14243 9435
rect 14277 9432 14289 9435
rect 14829 9435 14887 9441
rect 14829 9432 14841 9435
rect 14277 9404 14841 9432
rect 14277 9401 14289 9404
rect 14231 9395 14289 9401
rect 14829 9401 14841 9404
rect 14875 9401 14887 9435
rect 16761 9435 16819 9441
rect 16761 9432 16773 9435
rect 14829 9395 14887 9401
rect 15488 9404 16773 9432
rect 15488 9376 15516 9404
rect 16761 9401 16773 9404
rect 16807 9401 16819 9435
rect 16761 9395 16819 9401
rect 18506 9392 18512 9444
rect 18564 9392 18570 9444
rect 19702 9392 19708 9444
rect 19760 9392 19766 9444
rect 20070 9392 20076 9444
rect 20128 9392 20134 9444
rect 20625 9435 20683 9441
rect 20625 9401 20637 9435
rect 20671 9432 20683 9435
rect 22020 9432 22048 9460
rect 20671 9404 22048 9432
rect 20671 9401 20683 9404
rect 20625 9395 20683 9401
rect 22094 9392 22100 9444
rect 22152 9432 22158 9444
rect 22152 9404 22876 9432
rect 22152 9392 22158 9404
rect 7374 9324 7380 9376
rect 7432 9324 7438 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 9398 9364 9404 9376
rect 8536 9336 9404 9364
rect 8536 9324 8542 9336
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9490 9324 9496 9376
rect 9548 9324 9554 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 10042 9364 10048 9376
rect 9815 9336 10048 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10594 9324 10600 9376
rect 10652 9324 10658 9376
rect 15470 9324 15476 9376
rect 15528 9324 15534 9376
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 16117 9367 16175 9373
rect 16117 9364 16129 9367
rect 15712 9336 16129 9364
rect 15712 9324 15718 9336
rect 16117 9333 16129 9336
rect 16163 9333 16175 9367
rect 16117 9327 16175 9333
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 17678 9364 17684 9376
rect 16632 9336 17684 9364
rect 16632 9324 16638 9336
rect 17678 9324 17684 9336
rect 17736 9364 17742 9376
rect 18049 9367 18107 9373
rect 18049 9364 18061 9367
rect 17736 9336 18061 9364
rect 17736 9324 17742 9336
rect 18049 9333 18061 9336
rect 18095 9333 18107 9367
rect 18049 9327 18107 9333
rect 20898 9324 20904 9376
rect 20956 9324 20962 9376
rect 21174 9324 21180 9376
rect 21232 9324 21238 9376
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 21729 9367 21787 9373
rect 21729 9364 21741 9367
rect 21416 9336 21741 9364
rect 21416 9324 21422 9336
rect 21729 9333 21741 9336
rect 21775 9333 21787 9367
rect 21729 9327 21787 9333
rect 22554 9324 22560 9376
rect 22612 9324 22618 9376
rect 22848 9373 22876 9404
rect 22833 9367 22891 9373
rect 22833 9333 22845 9367
rect 22879 9333 22891 9367
rect 22833 9327 22891 9333
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 7834 9120 7840 9172
rect 7892 9120 7898 9172
rect 7926 9120 7932 9172
rect 7984 9120 7990 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8294 9160 8300 9172
rect 8159 9132 8300 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8754 9120 8760 9172
rect 8812 9120 8818 9172
rect 8938 9120 8944 9172
rect 8996 9120 9002 9172
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 9548 9132 9720 9160
rect 9548 9120 9554 9132
rect 7374 9024 7380 9036
rect 7208 8996 7380 9024
rect 7208 8820 7236 8996
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 7650 8984 7656 9036
rect 7708 8984 7714 9036
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 9024 7803 9027
rect 7852 9024 7880 9120
rect 7791 8996 7880 9024
rect 7791 8993 7803 8996
rect 7745 8987 7803 8993
rect 7926 8984 7932 9036
rect 7984 8984 7990 9036
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 8076 8996 8217 9024
rect 8076 8984 8082 8996
rect 8205 8993 8217 8996
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 8481 8987 8539 8993
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 8772 9024 8800 9120
rect 9508 9092 9536 9120
rect 9140 9064 9536 9092
rect 8849 9027 8907 9033
rect 8849 9024 8861 9027
rect 8772 8996 8861 9024
rect 8573 8987 8631 8993
rect 8849 8993 8861 8996
rect 8895 8993 8907 9027
rect 8849 8987 8907 8993
rect 7558 8916 7564 8968
rect 7616 8916 7622 8968
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8888 7343 8891
rect 7926 8888 7932 8900
rect 7331 8860 7932 8888
rect 7331 8857 7343 8860
rect 7285 8851 7343 8857
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 8496 8888 8524 8987
rect 8588 8956 8616 8987
rect 9140 8956 9168 9064
rect 9582 9052 9588 9104
rect 9640 9052 9646 9104
rect 9692 9092 9720 9132
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10502 9160 10508 9172
rect 10100 9132 10508 9160
rect 10100 9120 10106 9132
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 10612 9092 10640 9123
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 11020 9132 11805 9160
rect 11020 9120 11026 9132
rect 11793 9129 11805 9132
rect 11839 9129 11851 9163
rect 11793 9123 11851 9129
rect 12066 9120 12072 9172
rect 12124 9120 12130 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 15470 9160 15476 9172
rect 13412 9132 15476 9160
rect 13412 9120 13418 9132
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 16942 9120 16948 9172
rect 17000 9120 17006 9172
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 17184 9132 17233 9160
rect 17184 9120 17190 9132
rect 17221 9129 17233 9132
rect 17267 9129 17279 9163
rect 19334 9160 19340 9172
rect 17221 9123 17279 9129
rect 19168 9132 19340 9160
rect 11057 9095 11115 9101
rect 11057 9092 11069 9095
rect 9692 9064 10456 9092
rect 10612 9064 11069 9092
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9306 9024 9312 9036
rect 9263 8996 9312 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 9484 9027 9542 9033
rect 9484 8993 9496 9027
rect 9530 9024 9542 9027
rect 9600 9024 9628 9052
rect 9530 8996 9628 9024
rect 9530 8993 9542 8996
rect 9484 8987 9542 8993
rect 10428 8968 10456 9064
rect 11057 9061 11069 9064
rect 11103 9061 11115 9095
rect 11057 9055 11115 9061
rect 11238 9052 11244 9104
rect 11296 9092 11302 9104
rect 11698 9092 11704 9104
rect 11296 9064 11704 9092
rect 11296 9052 11302 9064
rect 11698 9052 11704 9064
rect 11756 9092 11762 9104
rect 13906 9092 13912 9104
rect 11756 9064 13912 9092
rect 11756 9052 11762 9064
rect 12176 9033 12204 9064
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 14001 9095 14059 9101
rect 14001 9061 14013 9095
rect 14047 9092 14059 9095
rect 15654 9092 15660 9104
rect 14047 9064 15660 9092
rect 14047 9061 14059 9064
rect 14001 9055 14059 9061
rect 15654 9052 15660 9064
rect 15712 9092 15718 9104
rect 17405 9095 17463 9101
rect 17405 9092 17417 9095
rect 15712 9064 17417 9092
rect 15712 9052 15718 9064
rect 17405 9061 17417 9064
rect 17451 9061 17463 9095
rect 17405 9055 17463 9061
rect 17954 9052 17960 9104
rect 18012 9092 18018 9104
rect 19168 9101 19196 9132
rect 19334 9120 19340 9132
rect 19392 9160 19398 9172
rect 21082 9160 21088 9172
rect 19392 9132 21088 9160
rect 19392 9120 19398 9132
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 21174 9120 21180 9172
rect 21232 9120 21238 9172
rect 21266 9120 21272 9172
rect 21324 9120 21330 9172
rect 21913 9163 21971 9169
rect 21913 9129 21925 9163
rect 21959 9160 21971 9163
rect 22554 9160 22560 9172
rect 21959 9132 22560 9160
rect 21959 9129 21971 9132
rect 21913 9123 21971 9129
rect 22554 9120 22560 9132
rect 22612 9120 22618 9172
rect 19153 9095 19211 9101
rect 19153 9092 19165 9095
rect 18012 9064 19165 9092
rect 18012 9052 18018 9064
rect 19153 9061 19165 9064
rect 19199 9061 19211 9095
rect 19153 9055 19211 9061
rect 19444 9064 20760 9092
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 12161 9027 12219 9033
rect 12161 8993 12173 9027
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 8588 8928 9168 8956
rect 10410 8916 10416 8968
rect 10468 8956 10474 8968
rect 11790 8956 11796 8968
rect 10468 8928 11796 8956
rect 10468 8916 10474 8928
rect 11790 8916 11796 8928
rect 11848 8956 11854 8968
rect 11900 8956 11928 8987
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 13538 9024 13544 9036
rect 12676 8996 13544 9024
rect 12676 8984 12682 8996
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13872 8996 14197 9024
rect 13872 8984 13878 8996
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 8993 16451 9027
rect 16393 8987 16451 8993
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 9024 16635 9027
rect 16853 9027 16911 9033
rect 16623 8996 16804 9024
rect 16623 8993 16635 8996
rect 16577 8987 16635 8993
rect 11848 8928 11928 8956
rect 11848 8916 11854 8928
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 13906 8956 13912 8968
rect 12584 8928 13912 8956
rect 12584 8916 12590 8928
rect 13906 8916 13912 8928
rect 13964 8916 13970 8968
rect 16408 8956 16436 8987
rect 16776 8956 16804 8996
rect 16853 8993 16865 9027
rect 16899 9024 16911 9027
rect 16942 9024 16948 9036
rect 16899 8996 16948 9024
rect 16899 8993 16911 8996
rect 16853 8987 16911 8993
rect 16942 8984 16948 8996
rect 17000 9024 17006 9036
rect 17000 8996 17264 9024
rect 17000 8984 17006 8996
rect 17034 8956 17040 8968
rect 16408 8928 16620 8956
rect 16776 8928 17040 8956
rect 16592 8900 16620 8928
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 17236 8956 17264 8996
rect 17310 8984 17316 9036
rect 17368 8984 17374 9036
rect 17972 8956 18000 9052
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 19444 9024 19472 9064
rect 20732 9033 20760 9064
rect 18840 8996 19472 9024
rect 19512 9027 19570 9033
rect 18840 8984 18846 8996
rect 19512 8993 19524 9027
rect 19558 9024 19570 9027
rect 20717 9027 20775 9033
rect 19558 8996 20576 9024
rect 19558 8993 19570 8996
rect 19512 8987 19570 8993
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 17236 8928 18000 8956
rect 18708 8928 19257 8956
rect 8496 8860 8800 8888
rect 8386 8820 8392 8832
rect 7208 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 8772 8820 8800 8860
rect 12986 8848 12992 8900
rect 13044 8888 13050 8900
rect 14642 8888 14648 8900
rect 13044 8860 14648 8888
rect 13044 8848 13050 8860
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 16574 8848 16580 8900
rect 16632 8848 16638 8900
rect 18708 8832 18736 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 9858 8820 9864 8832
rect 8772 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 12529 8823 12587 8829
rect 12529 8820 12541 8823
rect 12492 8792 12541 8820
rect 12492 8780 12498 8792
rect 12529 8789 12541 8792
rect 12575 8789 12587 8823
rect 12529 8783 12587 8789
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 15562 8820 15568 8832
rect 13412 8792 15568 8820
rect 13412 8780 13418 8792
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 18690 8780 18696 8832
rect 18748 8780 18754 8832
rect 20548 8820 20576 8996
rect 20717 8993 20729 9027
rect 20763 8993 20775 9027
rect 20717 8987 20775 8993
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 21192 9024 21220 9120
rect 21284 9092 21312 9120
rect 21284 9064 21864 9092
rect 21836 9033 21864 9064
rect 22278 9052 22284 9104
rect 22336 9052 22342 9104
rect 22370 9052 22376 9104
rect 22428 9052 22434 9104
rect 20947 8996 21220 9024
rect 21361 9027 21419 9033
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 21361 8993 21373 9027
rect 21407 8993 21419 9027
rect 21361 8987 21419 8993
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 8993 21879 9027
rect 21821 8987 21879 8993
rect 21376 8956 21404 8987
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22097 9027 22155 9033
rect 22097 9024 22109 9027
rect 22060 8996 22109 9024
rect 22060 8984 22066 8996
rect 22097 8993 22109 8996
rect 22143 8993 22155 9027
rect 22097 8987 22155 8993
rect 22296 8956 22324 9052
rect 22388 9023 22416 9052
rect 22373 9017 22431 9023
rect 22373 8983 22385 9017
rect 22419 8983 22431 9017
rect 22373 8977 22431 8983
rect 20640 8928 21404 8956
rect 21468 8928 22324 8956
rect 20640 8897 20668 8928
rect 20625 8891 20683 8897
rect 20625 8857 20637 8891
rect 20671 8857 20683 8891
rect 21468 8888 21496 8928
rect 20625 8851 20683 8857
rect 20732 8860 21496 8888
rect 21637 8891 21695 8897
rect 20732 8820 20760 8860
rect 21637 8857 21649 8891
rect 21683 8888 21695 8891
rect 28258 8888 28264 8900
rect 21683 8860 28264 8888
rect 21683 8857 21695 8860
rect 21637 8851 21695 8857
rect 28258 8848 28264 8860
rect 28316 8848 28322 8900
rect 20548 8792 20760 8820
rect 20806 8780 20812 8832
rect 20864 8780 20870 8832
rect 20990 8780 20996 8832
rect 21048 8820 21054 8832
rect 22002 8820 22008 8832
rect 21048 8792 22008 8820
rect 21048 8780 21054 8792
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 22186 8780 22192 8832
rect 22244 8780 22250 8832
rect 22462 8780 22468 8832
rect 22520 8780 22526 8832
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 9214 8616 9220 8628
rect 8444 8588 9220 8616
rect 8444 8576 8450 8588
rect 9214 8576 9220 8588
rect 9272 8616 9278 8628
rect 10686 8616 10692 8628
rect 9272 8588 10692 8616
rect 9272 8576 9278 8588
rect 10686 8576 10692 8588
rect 10744 8616 10750 8628
rect 11054 8616 11060 8628
rect 10744 8588 11060 8616
rect 10744 8576 10750 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 12526 8616 12532 8628
rect 11287 8588 12532 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 12713 8619 12771 8625
rect 12713 8585 12725 8619
rect 12759 8616 12771 8619
rect 13446 8616 13452 8628
rect 12759 8588 13452 8616
rect 12759 8585 12771 8588
rect 12713 8579 12771 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 16715 8619 16773 8625
rect 16715 8616 16727 8619
rect 14332 8588 16727 8616
rect 14332 8576 14338 8588
rect 16715 8585 16727 8588
rect 16761 8585 16773 8619
rect 18322 8616 18328 8628
rect 16715 8579 16773 8585
rect 17420 8588 18328 8616
rect 8113 8551 8171 8557
rect 8113 8517 8125 8551
rect 8159 8548 8171 8551
rect 8570 8548 8576 8560
rect 8159 8520 8576 8548
rect 8159 8517 8171 8520
rect 8113 8511 8171 8517
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 8662 8508 8668 8560
rect 8720 8508 8726 8560
rect 8757 8551 8815 8557
rect 8757 8517 8769 8551
rect 8803 8548 8815 8551
rect 11146 8548 11152 8560
rect 8803 8520 11152 8548
rect 8803 8517 8815 8520
rect 8757 8511 8815 8517
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 13170 8548 13176 8560
rect 11348 8520 13176 8548
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8478 8412 8484 8424
rect 8251 8384 8484 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 8680 8421 8708 8508
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 11238 8480 11244 8492
rect 8996 8452 9352 8480
rect 8996 8440 9002 8452
rect 9324 8421 9352 8452
rect 9600 8452 11244 8480
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8381 8723 8415
rect 8665 8375 8723 8381
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 8588 8344 8616 8375
rect 9033 8347 9091 8353
rect 9033 8344 9045 8347
rect 8588 8316 9045 8344
rect 9033 8313 9045 8316
rect 9079 8313 9091 8347
rect 9140 8344 9168 8375
rect 9600 8344 9628 8452
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 9950 8412 9956 8424
rect 9723 8384 9956 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 11348 8421 11376 8520
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 13265 8551 13323 8557
rect 13265 8517 13277 8551
rect 13311 8548 13323 8551
rect 13354 8548 13360 8560
rect 13311 8520 13360 8548
rect 13311 8517 13323 8520
rect 13265 8511 13323 8517
rect 13354 8508 13360 8520
rect 13412 8508 13418 8560
rect 14921 8551 14979 8557
rect 14921 8517 14933 8551
rect 14967 8517 14979 8551
rect 14921 8511 14979 8517
rect 11624 8452 12848 8480
rect 11624 8421 11652 8452
rect 11333 8415 11391 8421
rect 11333 8381 11345 8415
rect 11379 8381 11391 8415
rect 11333 8375 11391 8381
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12342 8412 12348 8424
rect 12299 8384 12348 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 9140 8316 9628 8344
rect 9033 8307 9091 8313
rect 9858 8304 9864 8356
rect 9916 8304 9922 8356
rect 10226 8304 10232 8356
rect 10284 8304 10290 8356
rect 10594 8304 10600 8356
rect 10652 8304 10658 8356
rect 11514 8304 11520 8356
rect 11572 8304 11578 8356
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 8481 8279 8539 8285
rect 8481 8276 8493 8279
rect 8444 8248 8493 8276
rect 8444 8236 8450 8248
rect 8481 8245 8493 8248
rect 8527 8245 8539 8279
rect 8481 8239 8539 8245
rect 10686 8236 10692 8288
rect 10744 8236 10750 8288
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 11330 8276 11336 8288
rect 10836 8248 11336 8276
rect 10836 8236 10842 8248
rect 11330 8236 11336 8248
rect 11388 8276 11394 8288
rect 11716 8276 11744 8375
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 12526 8372 12532 8424
rect 12584 8372 12590 8424
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8412 12679 8415
rect 12710 8412 12716 8424
rect 12667 8384 12716 8412
rect 12667 8381 12679 8384
rect 12621 8375 12679 8381
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 11790 8304 11796 8356
rect 11848 8304 11854 8356
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 12161 8347 12219 8353
rect 12161 8344 12173 8347
rect 11940 8316 12173 8344
rect 11940 8304 11946 8316
rect 12161 8313 12173 8316
rect 12207 8313 12219 8347
rect 12161 8307 12219 8313
rect 12437 8347 12495 8353
rect 12437 8313 12449 8347
rect 12483 8344 12495 8347
rect 12483 8316 12756 8344
rect 12483 8313 12495 8316
rect 12437 8307 12495 8313
rect 12728 8288 12756 8316
rect 11388 8248 11744 8276
rect 11388 8236 11394 8248
rect 12710 8236 12716 8288
rect 12768 8236 12774 8288
rect 12820 8276 12848 8452
rect 12894 8440 12900 8492
rect 12952 8480 12958 8492
rect 12952 8452 13216 8480
rect 12952 8440 12958 8452
rect 13078 8372 13084 8424
rect 13136 8372 13142 8424
rect 13188 8421 13216 8452
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 13797 8415 13855 8421
rect 13797 8412 13809 8415
rect 13688 8384 13809 8412
rect 13688 8372 13694 8384
rect 13797 8381 13809 8384
rect 13843 8381 13855 8415
rect 14936 8412 14964 8511
rect 15194 8508 15200 8560
rect 15252 8508 15258 8560
rect 16546 8520 16758 8548
rect 15212 8480 15240 8508
rect 16546 8480 16574 8520
rect 15212 8452 16574 8480
rect 15105 8415 15163 8421
rect 15105 8412 15117 8415
rect 14936 8384 15117 8412
rect 13797 8375 13855 8381
rect 15105 8381 15117 8384
rect 15151 8381 15163 8415
rect 15105 8375 15163 8381
rect 15841 8415 15899 8421
rect 15841 8381 15853 8415
rect 15887 8412 15899 8415
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15887 8384 16037 8412
rect 15887 8381 15899 8384
rect 15841 8375 15899 8381
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 16117 8415 16175 8421
rect 16117 8381 16129 8415
rect 16163 8412 16175 8415
rect 16553 8415 16611 8421
rect 16553 8412 16565 8415
rect 16163 8384 16565 8412
rect 16163 8381 16175 8384
rect 16117 8375 16175 8381
rect 16546 8381 16565 8384
rect 16599 8381 16611 8415
rect 16730 8412 16758 8520
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 16786 8423 16844 8429
rect 16786 8412 16798 8423
rect 16730 8389 16798 8412
rect 16832 8389 16844 8423
rect 16730 8384 16844 8389
rect 16786 8383 16844 8384
rect 16546 8375 16611 8381
rect 13081 8369 13139 8372
rect 12986 8304 12992 8356
rect 13044 8304 13050 8356
rect 15470 8304 15476 8356
rect 15528 8304 15534 8356
rect 15654 8304 15660 8356
rect 15712 8344 15718 8356
rect 16132 8344 16160 8375
rect 15712 8316 16160 8344
rect 16546 8344 16574 8375
rect 16960 8344 16988 8440
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 17218 8372 17224 8424
rect 17276 8412 17282 8424
rect 17420 8421 17448 8588
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 22097 8619 22155 8625
rect 22097 8616 22109 8619
rect 20456 8588 22109 8616
rect 18340 8520 18736 8548
rect 17589 8483 17647 8489
rect 17589 8449 17601 8483
rect 17635 8480 17647 8483
rect 18340 8480 18368 8520
rect 17635 8452 18368 8480
rect 17635 8449 17647 8452
rect 17589 8443 17647 8449
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 17276 8384 17325 8412
rect 17276 8372 17282 8384
rect 17313 8381 17325 8384
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 17405 8415 17463 8421
rect 17773 8415 17831 8421
rect 17405 8381 17417 8415
rect 17451 8381 17463 8415
rect 17405 8375 17463 8381
rect 17681 8409 17739 8415
rect 17681 8375 17693 8409
rect 17727 8375 17739 8409
rect 17773 8381 17785 8415
rect 17819 8412 17831 8415
rect 17954 8412 17960 8424
rect 17819 8384 17960 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 17681 8369 17739 8375
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18708 8421 18736 8520
rect 18782 8508 18788 8560
rect 18840 8508 18846 8560
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 19153 8415 19211 8421
rect 19153 8381 19165 8415
rect 19199 8381 19211 8415
rect 19153 8375 19211 8381
rect 19420 8415 19478 8421
rect 19420 8381 19432 8415
rect 19466 8412 19478 8415
rect 20456 8412 20484 8588
rect 22097 8585 22109 8588
rect 22143 8585 22155 8619
rect 22097 8579 22155 8585
rect 20533 8551 20591 8557
rect 20533 8517 20545 8551
rect 20579 8517 20591 8551
rect 22370 8548 22376 8560
rect 20533 8511 20591 8517
rect 21376 8520 22376 8548
rect 19466 8384 20484 8412
rect 20548 8412 20576 8511
rect 21376 8424 21404 8520
rect 22370 8508 22376 8520
rect 22428 8508 22434 8560
rect 31662 8480 31668 8492
rect 21652 8452 31668 8480
rect 20717 8415 20775 8421
rect 20717 8412 20729 8415
rect 20548 8384 20729 8412
rect 19466 8381 19478 8384
rect 19420 8375 19478 8381
rect 20717 8381 20729 8384
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 16546 8316 16988 8344
rect 15712 8304 15718 8316
rect 14550 8276 14556 8288
rect 12820 8248 14556 8276
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 15562 8276 15568 8288
rect 15252 8248 15568 8276
rect 15252 8236 15258 8248
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 16485 8279 16543 8285
rect 16485 8276 16497 8279
rect 16264 8248 16497 8276
rect 16264 8236 16270 8248
rect 16485 8245 16497 8248
rect 16531 8245 16543 8279
rect 16485 8239 16543 8245
rect 17034 8236 17040 8288
rect 17092 8236 17098 8288
rect 17696 8276 17724 8369
rect 17862 8304 17868 8356
rect 17920 8304 17926 8356
rect 18049 8347 18107 8353
rect 18049 8313 18061 8347
rect 18095 8344 18107 8347
rect 18322 8344 18328 8356
rect 18095 8316 18328 8344
rect 18095 8313 18107 8316
rect 18049 8307 18107 8313
rect 18322 8304 18328 8316
rect 18380 8304 18386 8356
rect 18417 8347 18475 8353
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 18598 8344 18604 8356
rect 18463 8316 18604 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 19168 8344 19196 8375
rect 21358 8372 21364 8424
rect 21416 8372 21422 8424
rect 21450 8372 21456 8424
rect 21508 8372 21514 8424
rect 18708 8316 19196 8344
rect 18708 8288 18736 8316
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 20036 8316 21281 8344
rect 20036 8304 20042 8316
rect 21269 8313 21281 8316
rect 21315 8313 21327 8347
rect 21269 8307 21327 8313
rect 21542 8304 21548 8356
rect 21600 8304 21606 8356
rect 18138 8276 18144 8288
rect 17696 8248 18144 8276
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 18690 8236 18696 8288
rect 18748 8236 18754 8288
rect 20993 8279 21051 8285
rect 20993 8245 21005 8279
rect 21039 8276 21051 8279
rect 21652 8276 21680 8452
rect 31662 8440 31668 8452
rect 31720 8440 31726 8492
rect 21726 8372 21732 8424
rect 21784 8372 21790 8424
rect 22002 8372 22008 8424
rect 22060 8372 22066 8424
rect 21039 8248 21680 8276
rect 21039 8245 21051 8248
rect 20993 8239 21051 8245
rect 21818 8236 21824 8288
rect 21876 8236 21882 8288
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8478 8072 8484 8084
rect 8435 8044 8484 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 10594 8032 10600 8084
rect 10652 8032 10658 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12584 8044 13001 8072
rect 12584 8032 12590 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13817 8075 13875 8081
rect 13817 8072 13829 8075
rect 13679 8044 13829 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13817 8041 13829 8044
rect 13863 8041 13875 8075
rect 13817 8035 13875 8041
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14967 8075 15025 8081
rect 14967 8072 14979 8075
rect 14240 8044 14979 8072
rect 14240 8032 14246 8044
rect 14967 8041 14979 8044
rect 15013 8041 15025 8075
rect 14967 8035 15025 8041
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 17405 8075 17463 8081
rect 17405 8072 17417 8075
rect 15703 8044 17417 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 17405 8041 17417 8044
rect 17451 8041 17463 8075
rect 17405 8035 17463 8041
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 20806 8072 20812 8084
rect 17727 8044 20812 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 20806 8032 20812 8044
rect 20864 8032 20870 8084
rect 8570 7964 8576 8016
rect 8628 8004 8634 8016
rect 9462 8007 9520 8013
rect 9462 8004 9474 8007
rect 8628 7976 9474 8004
rect 8628 7964 8634 7976
rect 9462 7973 9474 7976
rect 9508 7973 9520 8007
rect 9462 7967 9520 7973
rect 11238 7964 11244 8016
rect 11296 7964 11302 8016
rect 12253 8007 12311 8013
rect 11992 7976 12204 8004
rect 8481 7939 8539 7945
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 8662 7936 8668 7948
rect 8527 7908 8668 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 8846 7936 8852 7948
rect 8803 7908 8852 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 9030 7896 9036 7948
rect 9088 7896 9094 7948
rect 9214 7896 9220 7948
rect 9272 7896 9278 7948
rect 10410 7896 10416 7948
rect 10468 7936 10474 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10468 7908 11161 7936
rect 10468 7896 10474 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11256 7936 11284 7964
rect 11992 7945 12020 7976
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11256 7908 11621 7936
rect 11149 7899 11207 7905
rect 11609 7905 11621 7908
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7905 12035 7939
rect 11977 7899 12035 7905
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7905 12127 7939
rect 12176 7936 12204 7976
rect 12253 7973 12265 8007
rect 12299 8004 12311 8007
rect 12342 8004 12348 8016
rect 12299 7976 12348 8004
rect 12299 7973 12311 7976
rect 12253 7967 12311 7973
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 12768 7976 13277 8004
rect 12768 7964 12774 7976
rect 13265 7973 13277 7976
rect 13311 7973 13323 8007
rect 13265 7967 13323 7973
rect 13538 7964 13544 8016
rect 13596 8004 13602 8016
rect 16206 8004 16212 8016
rect 13596 7976 14964 8004
rect 13596 7964 13602 7976
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 12176 7908 13093 7936
rect 12069 7899 12127 7905
rect 13081 7905 13093 7908
rect 13127 7936 13139 7939
rect 13127 7908 13308 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 12084 7868 12112 7899
rect 13170 7868 13176 7880
rect 12084 7840 13176 7868
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 8711 7772 9260 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 9232 7732 9260 7772
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 11664 7772 12388 7800
rect 11664 7760 11670 7772
rect 9858 7732 9864 7744
rect 9232 7704 9864 7732
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11241 7735 11299 7741
rect 11241 7732 11253 7735
rect 11020 7704 11253 7732
rect 11020 7692 11026 7704
rect 11241 7701 11253 7704
rect 11287 7701 11299 7735
rect 11241 7695 11299 7701
rect 11698 7692 11704 7744
rect 11756 7692 11762 7744
rect 12360 7741 12388 7772
rect 12434 7760 12440 7812
rect 12492 7800 12498 7812
rect 12710 7800 12716 7812
rect 12492 7772 12716 7800
rect 12492 7760 12498 7772
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7701 12403 7735
rect 13280 7732 13308 7908
rect 13354 7896 13360 7948
rect 13412 7896 13418 7948
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 13814 7936 13820 7948
rect 13679 7908 13820 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 13464 7800 13492 7899
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 13909 7939 13967 7945
rect 13909 7905 13921 7939
rect 13955 7936 13967 7939
rect 14090 7936 14096 7948
rect 13955 7908 14096 7936
rect 13955 7905 13967 7908
rect 13909 7899 13967 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7936 14243 7939
rect 14274 7936 14280 7948
rect 14231 7908 14280 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7936 14427 7939
rect 14458 7936 14464 7948
rect 14415 7908 14464 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 14792 7908 14841 7936
rect 14792 7896 14798 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14936 7936 14964 7976
rect 15672 7976 16212 8004
rect 15038 7945 15096 7951
rect 15672 7945 15700 7976
rect 16206 7964 16212 7976
rect 16264 7964 16270 8016
rect 17034 8004 17040 8016
rect 16500 7976 17040 8004
rect 16500 7945 16528 7976
rect 17034 7964 17040 7976
rect 17092 7964 17098 8016
rect 18414 8004 18420 8016
rect 17788 7976 18420 8004
rect 15038 7936 15050 7945
rect 14936 7911 15050 7936
rect 15084 7911 15096 7945
rect 14936 7908 15096 7911
rect 15038 7905 15096 7908
rect 15197 7939 15255 7945
rect 15197 7905 15209 7939
rect 15243 7905 15255 7939
rect 14829 7899 14887 7905
rect 15197 7899 15255 7905
rect 15473 7939 15531 7945
rect 15473 7905 15485 7939
rect 15519 7905 15531 7939
rect 15473 7899 15531 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15749 7939 15807 7945
rect 15749 7905 15761 7939
rect 15795 7936 15807 7939
rect 16485 7939 16543 7945
rect 15795 7908 16436 7936
rect 15795 7905 15807 7908
rect 15749 7899 15807 7905
rect 14461 7803 14519 7809
rect 13464 7772 14228 7800
rect 13722 7732 13728 7744
rect 13280 7704 13728 7732
rect 12345 7695 12403 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14090 7692 14096 7744
rect 14148 7692 14154 7744
rect 14200 7732 14228 7772
rect 14461 7769 14473 7803
rect 14507 7800 14519 7803
rect 15212 7800 15240 7899
rect 14507 7772 15240 7800
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 14737 7735 14795 7741
rect 14737 7732 14749 7735
rect 14200 7704 14749 7732
rect 14737 7701 14749 7704
rect 14783 7701 14795 7735
rect 14737 7695 14795 7701
rect 15289 7735 15347 7741
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 15378 7732 15384 7744
rect 15335 7704 15384 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 15488 7732 15516 7899
rect 16408 7880 16436 7908
rect 16485 7905 16497 7939
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 16574 7896 16580 7948
rect 16632 7896 16638 7948
rect 17126 7896 17132 7948
rect 17184 7896 17190 7948
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7936 17555 7939
rect 17678 7936 17684 7948
rect 17543 7908 17684 7936
rect 17543 7905 17555 7908
rect 17497 7899 17555 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17788 7945 17816 7976
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 18509 8007 18567 8013
rect 18509 7973 18521 8007
rect 18555 8004 18567 8007
rect 21818 8004 21824 8016
rect 18555 7976 21824 8004
rect 18555 7973 18567 7976
rect 18509 7967 18567 7973
rect 21818 7964 21824 7976
rect 21876 7964 21882 8016
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 18049 7939 18107 7945
rect 18049 7905 18061 7939
rect 18095 7936 18107 7939
rect 18138 7936 18144 7948
rect 18095 7908 18144 7936
rect 18095 7905 18107 7908
rect 18049 7899 18107 7905
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 18960 7939 19018 7945
rect 18960 7905 18972 7939
rect 19006 7936 19018 7939
rect 19426 7936 19432 7948
rect 19006 7908 19432 7936
rect 19006 7905 19018 7908
rect 18960 7899 19018 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 20257 7939 20315 7945
rect 20257 7936 20269 7939
rect 20088 7908 20269 7936
rect 16390 7828 16396 7880
rect 16448 7828 16454 7880
rect 16592 7868 16620 7896
rect 18690 7868 18696 7880
rect 16592 7840 18696 7868
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 15841 7803 15899 7809
rect 15841 7769 15853 7803
rect 15887 7800 15899 7803
rect 16666 7800 16672 7812
rect 15887 7772 16672 7800
rect 15887 7769 15899 7772
rect 15841 7763 15899 7769
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 20088 7809 20116 7908
rect 20257 7905 20269 7908
rect 20303 7905 20315 7939
rect 20257 7899 20315 7905
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 20990 7936 20996 7948
rect 20763 7908 20996 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 21726 7868 21732 7880
rect 20855 7840 21732 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 20073 7803 20131 7809
rect 20073 7769 20085 7803
rect 20119 7769 20131 7803
rect 21266 7800 21272 7812
rect 20073 7763 20131 7769
rect 20456 7772 21272 7800
rect 16393 7735 16451 7741
rect 16393 7732 16405 7735
rect 15488 7704 16405 7732
rect 16393 7701 16405 7704
rect 16439 7701 16451 7735
rect 16393 7695 16451 7701
rect 17037 7735 17095 7741
rect 17037 7701 17049 7735
rect 17083 7732 17095 7735
rect 17402 7732 17408 7744
rect 17083 7704 17408 7732
rect 17083 7701 17095 7704
rect 17037 7695 17095 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 18417 7735 18475 7741
rect 18417 7701 18429 7735
rect 18463 7732 18475 7735
rect 20456 7732 20484 7772
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 18463 7704 20484 7732
rect 18463 7701 18475 7704
rect 18417 7695 18475 7701
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 9677 7531 9735 7537
rect 7708 7500 8984 7528
rect 7708 7488 7714 7500
rect 8956 7460 8984 7500
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 10410 7528 10416 7540
rect 9723 7500 10416 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 12618 7528 12624 7540
rect 10704 7500 12624 7528
rect 10229 7463 10287 7469
rect 10229 7460 10241 7463
rect 8956 7432 10241 7460
rect 10229 7429 10241 7432
rect 10275 7429 10287 7463
rect 10229 7423 10287 7429
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9401 7395 9459 7401
rect 9088 7364 9352 7392
rect 9088 7352 9094 7364
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 9324 7333 9352 7364
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 10134 7392 10140 7404
rect 9447 7364 10140 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10594 7392 10600 7404
rect 10244 7364 10600 7392
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8720 7296 8953 7324
rect 8720 7284 8726 7296
rect 8941 7293 8953 7296
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7326 9827 7327
rect 9953 7327 10011 7333
rect 9953 7326 9965 7327
rect 9815 7298 9965 7326
rect 9815 7293 9827 7298
rect 9769 7287 9827 7293
rect 9953 7293 9965 7298
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7324 10103 7327
rect 10244 7324 10272 7364
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10704 7401 10732 7500
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 12710 7488 12716 7540
rect 12768 7488 12774 7540
rect 13170 7488 13176 7540
rect 13228 7488 13234 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13354 7528 13360 7540
rect 13311 7500 13360 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 14458 7528 14464 7540
rect 13780 7500 14464 7528
rect 13780 7488 13786 7500
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 15378 7488 15384 7540
rect 15436 7528 15442 7540
rect 16206 7528 16212 7540
rect 15436 7500 16212 7528
rect 15436 7488 15442 7500
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 16390 7488 16396 7540
rect 16448 7528 16454 7540
rect 17678 7528 17684 7540
rect 16448 7500 17684 7528
rect 16448 7488 16454 7500
rect 17678 7488 17684 7500
rect 17736 7528 17742 7540
rect 17736 7500 17908 7528
rect 17736 7488 17742 7500
rect 12069 7463 12127 7469
rect 12069 7429 12081 7463
rect 12115 7460 12127 7463
rect 12342 7460 12348 7472
rect 12115 7432 12348 7460
rect 12115 7429 12127 7432
rect 12069 7423 12127 7429
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 12526 7460 12532 7472
rect 12452 7432 12532 7460
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 10091 7296 10272 7324
rect 10321 7327 10379 7333
rect 10091 7293 10103 7296
rect 10045 7287 10103 7293
rect 10321 7293 10333 7327
rect 10367 7324 10379 7327
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10367 7296 10425 7324
rect 10367 7293 10379 7296
rect 10321 7287 10379 7293
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 12452 7324 12480 7432
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 12728 7460 12756 7488
rect 12636 7432 12756 7460
rect 13188 7460 13216 7488
rect 13817 7463 13875 7469
rect 13817 7460 13829 7463
rect 13188 7432 13829 7460
rect 10551 7296 12480 7324
rect 12529 7327 12587 7333
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 12529 7293 12541 7327
rect 12575 7324 12587 7327
rect 12636 7324 12664 7432
rect 13817 7429 13829 7432
rect 13863 7429 13875 7463
rect 17880 7460 17908 7500
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 19242 7528 19248 7540
rect 18472 7500 19248 7528
rect 18472 7488 18478 7500
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19889 7531 19947 7537
rect 19889 7497 19901 7531
rect 19935 7528 19947 7531
rect 20070 7528 20076 7540
rect 19935 7500 20076 7528
rect 19935 7497 19947 7500
rect 19889 7491 19947 7497
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20165 7531 20223 7537
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 20254 7528 20260 7540
rect 20211 7500 20260 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 20254 7488 20260 7500
rect 20312 7488 20318 7540
rect 20441 7531 20499 7537
rect 20441 7497 20453 7531
rect 20487 7528 20499 7531
rect 22002 7528 22008 7540
rect 20487 7500 22008 7528
rect 20487 7497 20499 7500
rect 20441 7491 20499 7497
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 17880 7432 19380 7460
rect 13817 7423 13875 7429
rect 12575 7296 12664 7324
rect 12820 7364 13952 7392
rect 12575 7293 12587 7296
rect 12529 7287 12587 7293
rect 8956 7188 8984 7287
rect 9030 7216 9036 7268
rect 9088 7216 9094 7268
rect 9324 7256 9352 7287
rect 10060 7256 10088 7287
rect 9324 7228 10088 7256
rect 10428 7256 10456 7287
rect 10428 7228 10548 7256
rect 10520 7200 10548 7228
rect 10778 7216 10784 7268
rect 10836 7256 10842 7268
rect 10934 7259 10992 7265
rect 10934 7256 10946 7259
rect 10836 7228 10946 7256
rect 10836 7216 10842 7228
rect 10934 7225 10946 7228
rect 10980 7225 10992 7259
rect 10934 7219 10992 7225
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 12342 7256 12348 7268
rect 11296 7228 12348 7256
rect 11296 7216 11302 7228
rect 12342 7216 12348 7228
rect 12400 7256 12406 7268
rect 12820 7256 12848 7364
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13078 7324 13084 7336
rect 12952 7296 13084 7324
rect 12952 7284 12958 7296
rect 13078 7284 13084 7296
rect 13136 7324 13142 7336
rect 13924 7333 13952 7364
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16632 7364 16957 7392
rect 16632 7352 16638 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 18598 7352 18604 7404
rect 18656 7352 18662 7404
rect 19352 7392 19380 7432
rect 19426 7420 19432 7472
rect 19484 7460 19490 7472
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 19484 7432 20729 7460
rect 19484 7420 19490 7432
rect 20717 7429 20729 7432
rect 20763 7429 20775 7463
rect 20717 7423 20775 7429
rect 21358 7420 21364 7472
rect 21416 7420 21422 7472
rect 19610 7392 19616 7404
rect 19352 7364 19616 7392
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 20070 7392 20076 7404
rect 19996 7364 20076 7392
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 13136 7296 13185 7324
rect 13136 7284 13142 7296
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7324 13967 7327
rect 13998 7324 14004 7336
rect 13955 7296 14004 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7324 15255 7327
rect 16592 7324 16620 7352
rect 15243 7296 16620 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 18616 7324 18644 7352
rect 18616 7296 18920 7324
rect 12400 7228 12848 7256
rect 12400 7216 12406 7228
rect 12986 7216 12992 7268
rect 13044 7216 13050 7268
rect 13538 7216 13544 7268
rect 13596 7256 13602 7268
rect 13596 7228 13952 7256
rect 13596 7216 13602 7228
rect 10502 7188 10508 7200
rect 8956 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 12308 7160 12449 7188
rect 12308 7148 12314 7160
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 12894 7148 12900 7200
rect 12952 7148 12958 7200
rect 13924 7188 13952 7228
rect 14090 7216 14096 7268
rect 14148 7216 14154 7268
rect 15013 7259 15071 7265
rect 15013 7225 15025 7259
rect 15059 7256 15071 7259
rect 15286 7256 15292 7268
rect 15059 7228 15292 7256
rect 15059 7225 15071 7228
rect 15013 7219 15071 7225
rect 15286 7216 15292 7228
rect 15344 7216 15350 7268
rect 15470 7265 15476 7268
rect 15464 7219 15476 7265
rect 15470 7216 15476 7219
rect 15528 7216 15534 7268
rect 16942 7216 16948 7268
rect 17000 7256 17006 7268
rect 17190 7259 17248 7265
rect 17190 7256 17202 7259
rect 17000 7228 17202 7256
rect 17000 7216 17006 7228
rect 17190 7225 17202 7228
rect 17236 7225 17248 7259
rect 17190 7219 17248 7225
rect 18785 7259 18843 7265
rect 18785 7225 18797 7259
rect 18831 7225 18843 7259
rect 18892 7256 18920 7296
rect 18966 7284 18972 7336
rect 19024 7324 19030 7336
rect 19245 7327 19303 7333
rect 19245 7324 19257 7327
rect 19024 7296 19257 7324
rect 19024 7284 19030 7296
rect 19245 7293 19257 7296
rect 19291 7293 19303 7327
rect 19245 7287 19303 7293
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19996 7333 20024 7364
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 21376 7392 21404 7420
rect 20364 7364 21404 7392
rect 20257 7337 20315 7343
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 19392 7296 19717 7324
rect 19392 7284 19398 7296
rect 19705 7293 19717 7296
rect 19751 7293 19763 7327
rect 19705 7287 19763 7293
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7293 20039 7327
rect 20257 7324 20269 7337
rect 19981 7287 20039 7293
rect 20180 7303 20269 7324
rect 20303 7303 20315 7337
rect 20364 7336 20392 7364
rect 20180 7297 20315 7303
rect 20180 7296 20300 7297
rect 20070 7256 20076 7268
rect 18892 7228 20076 7256
rect 18785 7219 18843 7225
rect 14185 7191 14243 7197
rect 14185 7188 14197 7191
rect 13924 7160 14197 7188
rect 14185 7157 14197 7160
rect 14231 7157 14243 7191
rect 14185 7151 14243 7157
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 14734 7188 14740 7200
rect 14516 7160 14740 7188
rect 14516 7148 14522 7160
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 14921 7191 14979 7197
rect 14921 7157 14933 7191
rect 14967 7188 14979 7191
rect 15378 7188 15384 7200
rect 14967 7160 15384 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 16574 7148 16580 7200
rect 16632 7148 16638 7200
rect 16761 7191 16819 7197
rect 16761 7157 16773 7191
rect 16807 7188 16819 7191
rect 17034 7188 17040 7200
rect 16807 7160 17040 7188
rect 16807 7157 16819 7160
rect 16761 7151 16819 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 18325 7191 18383 7197
rect 18325 7157 18337 7191
rect 18371 7188 18383 7191
rect 18800 7188 18828 7219
rect 20070 7216 20076 7228
rect 20128 7216 20134 7268
rect 18371 7160 18828 7188
rect 18371 7157 18383 7160
rect 18325 7151 18383 7157
rect 18874 7148 18880 7200
rect 18932 7148 18938 7200
rect 19334 7148 19340 7200
rect 19392 7148 19398 7200
rect 19426 7148 19432 7200
rect 19484 7188 19490 7200
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 19484 7160 19625 7188
rect 19484 7148 19490 7160
rect 19613 7157 19625 7160
rect 19659 7157 19671 7191
rect 19613 7151 19671 7157
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 20180 7188 20208 7296
rect 20346 7284 20352 7336
rect 20404 7284 20410 7336
rect 20622 7284 20628 7336
rect 20680 7284 20686 7336
rect 19944 7160 20208 7188
rect 19944 7148 19950 7160
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 7558 6944 7564 6996
rect 7616 6944 7622 6996
rect 7926 6944 7932 6996
rect 7984 6984 7990 6996
rect 7984 6956 8708 6984
rect 7984 6944 7990 6956
rect 7576 6916 7604 6944
rect 7576 6888 8616 6916
rect 8018 6808 8024 6860
rect 8076 6808 8082 6860
rect 8036 6712 8064 6808
rect 8588 6780 8616 6888
rect 8680 6848 8708 6956
rect 9030 6944 9036 6996
rect 9088 6944 9094 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 11330 6984 11336 6996
rect 10560 6956 11336 6984
rect 10560 6944 10566 6956
rect 11330 6944 11336 6956
rect 11388 6944 11394 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 11885 6987 11943 6993
rect 11885 6984 11897 6987
rect 11756 6956 11897 6984
rect 11756 6944 11762 6956
rect 11885 6953 11897 6956
rect 11931 6953 11943 6987
rect 11885 6947 11943 6953
rect 11992 6956 12434 6984
rect 9048 6916 9076 6944
rect 11992 6916 12020 6956
rect 12253 6919 12311 6925
rect 12253 6916 12265 6919
rect 9048 6888 10088 6916
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 8680 6820 9781 6848
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6848 9919 6851
rect 9950 6848 9956 6860
rect 9907 6820 9956 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10060 6857 10088 6888
rect 10980 6888 11284 6916
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10226 6848 10232 6860
rect 10183 6820 10232 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 10502 6808 10508 6860
rect 10560 6808 10566 6860
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 10980 6848 11008 6888
rect 10827 6820 11008 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11149 6851 11207 6857
rect 11149 6848 11161 6851
rect 11112 6820 11161 6848
rect 11112 6808 11118 6820
rect 11149 6817 11161 6820
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 8588 6752 10425 6780
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 8036 6684 10824 6712
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 9456 6616 10701 6644
rect 9456 6604 9462 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10796 6644 10824 6684
rect 11057 6647 11115 6653
rect 11057 6644 11069 6647
rect 10796 6616 11069 6644
rect 10689 6607 10747 6613
rect 11057 6613 11069 6616
rect 11103 6613 11115 6647
rect 11164 6644 11192 6811
rect 11256 6712 11284 6888
rect 11532 6888 12020 6916
rect 12084 6888 12265 6916
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11532 6848 11560 6888
rect 11471 6820 11560 6848
rect 11609 6851 11667 6857
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 11609 6817 11621 6851
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11624 6780 11652 6811
rect 11698 6808 11704 6860
rect 11756 6808 11762 6860
rect 12084 6857 12112 6888
rect 12253 6885 12265 6888
rect 12299 6885 12311 6919
rect 12406 6916 12434 6956
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 13872 6956 14657 6984
rect 13872 6944 13878 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 14645 6947 14703 6953
rect 15473 6987 15531 6993
rect 15473 6953 15485 6987
rect 15519 6984 15531 6987
rect 16390 6984 16396 6996
rect 15519 6956 16396 6984
rect 15519 6953 15531 6956
rect 15473 6947 15531 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 17034 6944 17040 6996
rect 17092 6984 17098 6996
rect 17221 6987 17279 6993
rect 17221 6984 17233 6987
rect 17092 6956 17233 6984
rect 17092 6944 17098 6956
rect 17221 6953 17233 6956
rect 17267 6953 17279 6987
rect 17221 6947 17279 6953
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 18690 6984 18696 6996
rect 18196 6956 18696 6984
rect 18196 6944 18202 6956
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 18966 6944 18972 6996
rect 19024 6944 19030 6996
rect 19245 6987 19303 6993
rect 19245 6953 19257 6987
rect 19291 6984 19303 6987
rect 19334 6984 19340 6996
rect 19291 6956 19340 6984
rect 19291 6953 19303 6956
rect 19245 6947 19303 6953
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 19610 6984 19616 6996
rect 19444 6956 19616 6984
rect 13078 6916 13084 6928
rect 12406 6888 13084 6916
rect 12253 6879 12311 6885
rect 13078 6876 13084 6888
rect 13136 6876 13142 6928
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 14792 6888 15884 6916
rect 14792 6876 14798 6888
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6817 11943 6851
rect 11885 6811 11943 6817
rect 12069 6851 12127 6857
rect 12069 6817 12081 6851
rect 12115 6817 12127 6851
rect 12069 6811 12127 6817
rect 11379 6752 11652 6780
rect 11716 6780 11744 6808
rect 11900 6780 11928 6811
rect 12158 6808 12164 6860
rect 12216 6808 12222 6860
rect 12618 6808 12624 6860
rect 12676 6808 12682 6860
rect 12894 6857 12900 6860
rect 12888 6811 12900 6857
rect 12894 6808 12900 6811
rect 12952 6808 12958 6860
rect 14458 6808 14464 6860
rect 14516 6808 14522 6860
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 12250 6780 12256 6792
rect 11716 6752 11836 6780
rect 11900 6752 12256 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11422 6712 11428 6724
rect 11256 6684 11428 6712
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 11701 6715 11759 6721
rect 11701 6712 11713 6715
rect 11572 6684 11713 6712
rect 11572 6672 11578 6684
rect 11701 6681 11713 6684
rect 11747 6681 11759 6715
rect 11701 6675 11759 6681
rect 11808 6644 11836 6752
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14568 6780 14596 6811
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 14829 6851 14887 6857
rect 14829 6848 14841 6851
rect 14700 6820 14841 6848
rect 14700 6808 14706 6820
rect 14829 6817 14841 6820
rect 14875 6817 14887 6851
rect 14829 6811 14887 6817
rect 15010 6808 15016 6860
rect 15068 6808 15074 6860
rect 15304 6857 15332 6888
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15381 6851 15439 6857
rect 15381 6817 15393 6851
rect 15427 6817 15439 6851
rect 15381 6811 15439 6817
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 13780 6752 14596 6780
rect 13780 6740 13786 6752
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 15396 6780 15424 6811
rect 15252 6752 15424 6780
rect 15252 6740 15258 6752
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 15672 6780 15700 6811
rect 15580 6752 15700 6780
rect 15856 6780 15884 6888
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16408 6848 16436 6944
rect 16574 6876 16580 6928
rect 16632 6916 16638 6928
rect 16669 6919 16727 6925
rect 16669 6916 16681 6919
rect 16632 6888 16681 6916
rect 16632 6876 16638 6888
rect 16669 6885 16681 6888
rect 16715 6885 16727 6919
rect 16669 6879 16727 6885
rect 16776 6888 17448 6916
rect 16347 6820 16436 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16776 6780 16804 6888
rect 17420 6857 17448 6888
rect 17313 6851 17371 6857
rect 17313 6817 17325 6851
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 17405 6851 17463 6857
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 17494 6848 17500 6860
rect 17451 6820 17500 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 15856 6752 16804 6780
rect 17328 6780 17356 6811
rect 17494 6808 17500 6820
rect 17552 6848 17558 6860
rect 17678 6848 17684 6860
rect 17552 6820 17684 6848
rect 17552 6808 17558 6820
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 17862 6808 17868 6860
rect 17920 6808 17926 6860
rect 18049 6851 18107 6857
rect 18049 6817 18061 6851
rect 18095 6848 18107 6851
rect 18095 6820 18368 6848
rect 18095 6817 18107 6820
rect 18049 6811 18107 6817
rect 18340 6792 18368 6820
rect 18506 6808 18512 6860
rect 18564 6808 18570 6860
rect 18601 6851 18659 6857
rect 18601 6817 18613 6851
rect 18647 6817 18659 6851
rect 18601 6811 18659 6817
rect 18877 6851 18935 6857
rect 18877 6817 18889 6851
rect 18923 6848 18935 6851
rect 19242 6848 19248 6860
rect 18923 6820 19248 6848
rect 18923 6817 18935 6820
rect 18877 6811 18935 6817
rect 17954 6780 17960 6792
rect 17328 6752 17960 6780
rect 14001 6715 14059 6721
rect 14001 6681 14013 6715
rect 14047 6712 14059 6715
rect 14090 6712 14096 6724
rect 14047 6684 14096 6712
rect 14047 6681 14059 6684
rect 14001 6675 14059 6681
rect 14090 6672 14096 6684
rect 14148 6672 14154 6724
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6712 14427 6715
rect 15488 6712 15516 6740
rect 14415 6684 15516 6712
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 15580 6656 15608 6752
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18322 6740 18328 6792
rect 18380 6740 18386 6792
rect 15749 6715 15807 6721
rect 15749 6681 15761 6715
rect 15795 6712 15807 6715
rect 16298 6712 16304 6724
rect 15795 6684 16304 6712
rect 15795 6681 15807 6684
rect 15749 6675 15807 6681
rect 16298 6672 16304 6684
rect 16356 6672 16362 6724
rect 16850 6672 16856 6724
rect 16908 6672 16914 6724
rect 17497 6715 17555 6721
rect 17497 6681 17509 6715
rect 17543 6712 17555 6715
rect 18616 6712 18644 6811
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19444 6857 19472 6956
rect 19610 6944 19616 6956
rect 19668 6984 19674 6996
rect 20349 6987 20407 6993
rect 19668 6956 20300 6984
rect 19668 6944 19674 6956
rect 20070 6876 20076 6928
rect 20128 6876 20134 6928
rect 19337 6851 19395 6857
rect 19337 6817 19349 6851
rect 19383 6817 19395 6851
rect 19337 6811 19395 6817
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 19352 6780 19380 6811
rect 19702 6808 19708 6860
rect 19760 6808 19766 6860
rect 19978 6808 19984 6860
rect 20036 6808 20042 6860
rect 20272 6857 20300 6956
rect 20349 6953 20361 6987
rect 20395 6984 20407 6987
rect 20622 6984 20628 6996
rect 20395 6956 20628 6984
rect 20395 6953 20407 6956
rect 20349 6947 20407 6953
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 20990 6944 20996 6996
rect 21048 6944 21054 6996
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 20257 6851 20315 6857
rect 20257 6817 20269 6851
rect 20303 6848 20315 6851
rect 21008 6848 21036 6944
rect 20303 6820 21036 6848
rect 20303 6817 20315 6820
rect 20257 6811 20315 6817
rect 19996 6780 20024 6808
rect 19352 6752 20024 6780
rect 17543 6684 18644 6712
rect 17543 6681 17555 6684
rect 17497 6675 17555 6681
rect 18782 6672 18788 6724
rect 18840 6712 18846 6724
rect 19797 6715 19855 6721
rect 19797 6712 19809 6715
rect 18840 6684 19809 6712
rect 18840 6672 18846 6684
rect 19797 6681 19809 6684
rect 19843 6681 19855 6715
rect 20180 6712 20208 6811
rect 22462 6712 22468 6724
rect 20180 6684 22468 6712
rect 19797 6675 19855 6681
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 11164 6616 11836 6644
rect 14921 6647 14979 6653
rect 11057 6607 11115 6613
rect 14921 6613 14933 6647
rect 14967 6644 14979 6647
rect 15197 6647 15255 6653
rect 15197 6644 15209 6647
rect 14967 6616 15209 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 15197 6613 15209 6616
rect 15243 6613 15255 6647
rect 15197 6607 15255 6613
rect 15562 6604 15568 6656
rect 15620 6604 15626 6656
rect 16390 6604 16396 6656
rect 16448 6604 16454 6656
rect 17957 6647 18015 6653
rect 17957 6613 17969 6647
rect 18003 6644 18015 6647
rect 18417 6647 18475 6653
rect 18417 6644 18429 6647
rect 18003 6616 18429 6644
rect 18003 6613 18015 6616
rect 17957 6607 18015 6613
rect 18417 6613 18429 6616
rect 18463 6613 18475 6647
rect 18417 6607 18475 6613
rect 19521 6647 19579 6653
rect 19521 6613 19533 6647
rect 19567 6644 19579 6647
rect 21450 6644 21456 6656
rect 19567 6616 21456 6644
rect 19567 6613 19579 6616
rect 19521 6607 19579 6613
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 10502 6400 10508 6452
rect 10560 6400 10566 6452
rect 10778 6400 10784 6452
rect 10836 6400 10842 6452
rect 11333 6443 11391 6449
rect 11333 6440 11345 6443
rect 10980 6412 11345 6440
rect 10520 6372 10548 6400
rect 10980 6372 11008 6412
rect 11333 6409 11345 6412
rect 11379 6409 11391 6443
rect 11333 6403 11391 6409
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 11480 6412 11621 6440
rect 11480 6400 11486 6412
rect 11609 6409 11621 6412
rect 11655 6409 11667 6443
rect 11609 6403 11667 6409
rect 11882 6400 11888 6452
rect 11940 6400 11946 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6440 12219 6443
rect 12342 6440 12348 6452
rect 12207 6412 12348 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 13722 6440 13728 6452
rect 12492 6412 13728 6440
rect 12492 6400 12498 6412
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 14645 6443 14703 6449
rect 14645 6440 14657 6443
rect 14608 6412 14657 6440
rect 14608 6400 14614 6412
rect 14645 6409 14657 6412
rect 14691 6409 14703 6443
rect 14645 6403 14703 6409
rect 15010 6400 15016 6452
rect 15068 6440 15074 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15068 6412 15577 6440
rect 15068 6400 15074 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 16390 6400 16396 6452
rect 16448 6400 16454 6452
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6440 16911 6443
rect 16942 6440 16948 6452
rect 16899 6412 16948 6440
rect 16899 6409 16911 6412
rect 16853 6403 16911 6409
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 17126 6400 17132 6452
rect 17184 6440 17190 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17184 6412 17417 6440
rect 17184 6400 17190 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17405 6403 17463 6409
rect 17770 6400 17776 6452
rect 17828 6400 17834 6452
rect 18782 6400 18788 6452
rect 18840 6400 18846 6452
rect 19426 6400 19432 6452
rect 19484 6400 19490 6452
rect 10520 6344 11008 6372
rect 11054 6332 11060 6384
rect 11112 6332 11118 6384
rect 12618 6372 12624 6384
rect 11164 6344 12624 6372
rect 8938 6196 8944 6248
rect 8996 6196 9002 6248
rect 9858 6196 9864 6248
rect 9916 6196 9922 6248
rect 10134 6196 10140 6248
rect 10192 6236 10198 6248
rect 11164 6245 11192 6344
rect 12618 6332 12624 6344
rect 12676 6332 12682 6384
rect 12710 6332 12716 6384
rect 12768 6332 12774 6384
rect 12989 6375 13047 6381
rect 12989 6341 13001 6375
rect 13035 6372 13047 6375
rect 13078 6372 13084 6384
rect 13035 6344 13084 6372
rect 13035 6341 13047 6344
rect 12989 6335 13047 6341
rect 13078 6332 13084 6344
rect 13136 6332 13142 6384
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 14277 6375 14335 6381
rect 14277 6372 14289 6375
rect 13320 6344 14289 6372
rect 13320 6332 13326 6344
rect 14277 6341 14289 6344
rect 14323 6341 14335 6375
rect 14277 6335 14335 6341
rect 15286 6332 15292 6384
rect 15344 6332 15350 6384
rect 11238 6264 11244 6316
rect 11296 6264 11302 6316
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11388 6276 12112 6304
rect 11388 6264 11394 6276
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 10192 6208 10701 6236
rect 10192 6196 10198 6208
rect 10689 6205 10701 6208
rect 10735 6205 10747 6239
rect 10689 6199 10747 6205
rect 10965 6239 11023 6245
rect 10965 6205 10977 6239
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 11149 6239 11207 6245
rect 11149 6205 11161 6239
rect 11195 6205 11207 6239
rect 11256 6236 11284 6264
rect 11716 6245 11744 6276
rect 11425 6239 11483 6245
rect 11425 6236 11437 6239
rect 11256 6208 11437 6236
rect 11149 6199 11207 6205
rect 11425 6205 11437 6208
rect 11471 6236 11483 6239
rect 11701 6239 11759 6245
rect 11471 6208 11652 6236
rect 11471 6205 11483 6208
rect 11425 6199 11483 6205
rect 8956 6100 8984 6196
rect 9876 6168 9904 6196
rect 10980 6168 11008 6199
rect 9876 6140 11008 6168
rect 11624 6168 11652 6208
rect 11701 6205 11713 6239
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11974 6196 11980 6248
rect 12032 6196 12038 6248
rect 12084 6238 12112 6276
rect 12268 6276 12449 6304
rect 12158 6238 12164 6248
rect 12084 6210 12164 6238
rect 12158 6196 12164 6210
rect 12216 6196 12222 6248
rect 12268 6245 12296 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 13096 6304 13124 6332
rect 15562 6304 15568 6316
rect 13096 6276 15568 6304
rect 12437 6267 12495 6273
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 12342 6196 12348 6248
rect 12400 6196 12406 6248
rect 13648 6245 13676 6276
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12544 6208 12633 6236
rect 12066 6168 12072 6180
rect 11624 6140 12072 6168
rect 12066 6128 12072 6140
rect 12124 6128 12130 6180
rect 12544 6100 12572 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6236 13231 6239
rect 13633 6239 13691 6245
rect 13219 6208 13400 6236
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 12710 6128 12716 6180
rect 12768 6128 12774 6180
rect 13096 6168 13124 6199
rect 13265 6171 13323 6177
rect 13265 6168 13277 6171
rect 13096 6140 13277 6168
rect 13265 6137 13277 6140
rect 13311 6137 13323 6171
rect 13265 6131 13323 6137
rect 8956 6072 12572 6100
rect 12728 6100 12756 6128
rect 13372 6100 13400 6208
rect 13633 6205 13645 6239
rect 13679 6205 13691 6239
rect 13633 6199 13691 6205
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13872 6208 13921 6236
rect 13872 6196 13878 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 13998 6196 14004 6248
rect 14056 6236 14062 6248
rect 14936 6245 14964 6276
rect 15562 6264 15568 6276
rect 15620 6304 15626 6316
rect 15620 6276 15792 6304
rect 15620 6264 15626 6276
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14056 6208 14381 6236
rect 14056 6196 14062 6208
rect 14369 6205 14381 6208
rect 14415 6236 14427 6239
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14415 6208 14565 6236
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6205 14979 6239
rect 14921 6199 14979 6205
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6236 15071 6239
rect 15197 6239 15255 6245
rect 15197 6236 15209 6239
rect 15059 6208 15209 6236
rect 15059 6205 15071 6208
rect 15013 6199 15071 6205
rect 15197 6205 15209 6208
rect 15243 6205 15255 6239
rect 15197 6199 15255 6205
rect 15654 6196 15660 6248
rect 15712 6196 15718 6248
rect 15764 6245 15792 6276
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 16206 6196 16212 6248
rect 16264 6196 16270 6248
rect 16408 6236 16436 6400
rect 18800 6372 18828 6400
rect 16960 6344 18828 6372
rect 16485 6239 16543 6245
rect 16485 6236 16497 6239
rect 16408 6208 16497 6236
rect 16485 6205 16497 6208
rect 16531 6205 16543 6239
rect 16485 6199 16543 6205
rect 16758 6196 16764 6248
rect 16816 6196 16822 6248
rect 16960 6245 16988 6344
rect 17494 6304 17500 6316
rect 17052 6276 17500 6304
rect 17052 6245 17080 6276
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 18046 6304 18052 6316
rect 17880 6276 18052 6304
rect 17880 6245 17908 6276
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 18138 6264 18144 6316
rect 18196 6264 18202 6316
rect 19444 6304 19472 6400
rect 18248 6276 19472 6304
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6205 17003 6239
rect 16945 6199 17003 6205
rect 17037 6239 17095 6245
rect 17037 6205 17049 6239
rect 17083 6205 17095 6239
rect 17037 6199 17095 6205
rect 17129 6239 17187 6245
rect 17129 6205 17141 6239
rect 17175 6236 17187 6239
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 17175 6208 17325 6236
rect 17175 6205 17187 6208
rect 17129 6199 17187 6205
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 17681 6239 17739 6245
rect 17681 6205 17693 6239
rect 17727 6205 17739 6239
rect 17681 6199 17739 6205
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6205 17923 6239
rect 17865 6199 17923 6205
rect 17957 6239 18015 6245
rect 17957 6205 17969 6239
rect 18003 6236 18015 6239
rect 18156 6236 18184 6264
rect 18248 6245 18276 6276
rect 18003 6208 18184 6236
rect 18233 6239 18291 6245
rect 18003 6205 18015 6208
rect 17957 6199 18015 6205
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6236 18475 6239
rect 21542 6236 21548 6248
rect 18463 6208 21548 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 13725 6171 13783 6177
rect 13725 6137 13737 6171
rect 13771 6168 13783 6171
rect 14090 6168 14096 6180
rect 13771 6140 14096 6168
rect 13771 6137 13783 6140
rect 13725 6131 13783 6137
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 14458 6128 14464 6180
rect 14516 6128 14522 6180
rect 16224 6168 16252 6196
rect 16393 6171 16451 6177
rect 16393 6168 16405 6171
rect 16224 6140 16405 6168
rect 16393 6137 16405 6140
rect 16439 6137 16451 6171
rect 16776 6168 16804 6196
rect 17696 6168 17724 6199
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 16776 6140 17724 6168
rect 16393 6131 16451 6137
rect 18322 6128 18328 6180
rect 18380 6168 18386 6180
rect 20898 6168 20904 6180
rect 18380 6140 20904 6168
rect 18380 6128 18386 6140
rect 20898 6128 20904 6140
rect 20956 6128 20962 6180
rect 12728 6072 13400 6100
rect 13998 6060 14004 6112
rect 14056 6060 14062 6112
rect 14476 6100 14504 6128
rect 15841 6103 15899 6109
rect 15841 6100 15853 6103
rect 14476 6072 15853 6100
rect 15841 6069 15853 6072
rect 15887 6069 15899 6103
rect 15841 6063 15899 6069
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6100 18107 6103
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 18095 6072 18245 6100
rect 18095 6069 18107 6072
rect 18049 6063 18107 6069
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 18233 6063 18291 6069
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 9674 5856 9680 5908
rect 9732 5856 9738 5908
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 9824 5868 11897 5896
rect 9824 5856 9830 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12529 5899 12587 5905
rect 12529 5896 12541 5899
rect 12124 5868 12541 5896
rect 12124 5856 12130 5868
rect 12529 5865 12541 5868
rect 12575 5896 12587 5899
rect 12710 5896 12716 5908
rect 12575 5868 12716 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 13044 5868 13553 5896
rect 13044 5856 13050 5868
rect 13541 5865 13553 5868
rect 13587 5865 13599 5899
rect 13541 5859 13599 5865
rect 13998 5856 14004 5908
rect 14056 5856 14062 5908
rect 14090 5856 14096 5908
rect 14148 5856 14154 5908
rect 9692 5760 9720 5856
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11204 5800 12112 5828
rect 11204 5788 11210 5800
rect 12084 5769 12112 5800
rect 11885 5763 11943 5769
rect 11885 5760 11897 5763
rect 9692 5732 11897 5760
rect 11885 5729 11897 5732
rect 11931 5729 11943 5763
rect 11885 5723 11943 5729
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 12161 5763 12219 5769
rect 12161 5729 12173 5763
rect 12207 5729 12219 5763
rect 12161 5723 12219 5729
rect 12253 5763 12311 5769
rect 12253 5729 12265 5763
rect 12299 5760 12311 5763
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 12299 5732 12449 5760
rect 12299 5729 12311 5732
rect 12253 5723 12311 5729
rect 12437 5729 12449 5732
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 13081 5763 13139 5769
rect 13081 5729 13093 5763
rect 13127 5760 13139 5763
rect 13173 5763 13231 5769
rect 13173 5760 13185 5763
rect 13127 5732 13185 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 13173 5729 13185 5732
rect 13219 5729 13231 5763
rect 13173 5723 13231 5729
rect 13265 5763 13323 5769
rect 13265 5729 13277 5763
rect 13311 5760 13323 5763
rect 13449 5763 13507 5769
rect 13449 5760 13461 5763
rect 13311 5732 13461 5760
rect 13311 5729 13323 5732
rect 13265 5723 13323 5729
rect 13449 5729 13461 5732
rect 13495 5729 13507 5763
rect 13449 5723 13507 5729
rect 11698 5652 11704 5704
rect 11756 5692 11762 5704
rect 12176 5692 12204 5723
rect 13096 5692 13124 5723
rect 13906 5720 13912 5772
rect 13964 5720 13970 5772
rect 14016 5760 14044 5856
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 14016 5732 14105 5760
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 11756 5664 12204 5692
rect 12452 5664 13124 5692
rect 11756 5652 11762 5664
rect 12452 5636 12480 5664
rect 12434 5584 12440 5636
rect 12492 5584 12498 5636
rect 12986 5516 12992 5568
rect 13044 5516 13050 5568
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 12345 5355 12403 5361
rect 12345 5352 12357 5355
rect 11112 5324 12357 5352
rect 11112 5312 11118 5324
rect 12345 5321 12357 5324
rect 12391 5321 12403 5355
rect 12345 5315 12403 5321
rect 12618 5312 12624 5364
rect 12676 5312 12682 5364
rect 12894 5312 12900 5364
rect 12952 5352 12958 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12952 5324 13001 5352
rect 12952 5312 12958 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12452 5080 12480 5111
rect 12526 5108 12532 5160
rect 12584 5108 12590 5160
rect 12710 5108 12716 5160
rect 12768 5108 12774 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 12986 5148 12992 5160
rect 12943 5120 12992 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 12728 5080 12756 5108
rect 12452 5052 12756 5080
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 18046 4128 18052 4140
rect 14424 4100 18052 4128
rect 14424 4088 14430 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 14090 3516 14096 3528
rect 12400 3488 14096 3516
rect 12400 3476 12406 3488
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
rect 16022 416 16028 468
rect 16080 456 16086 468
rect 16482 456 16488 468
rect 16080 428 16488 456
rect 16080 416 16086 428
rect 16482 416 16488 428
rect 16540 416 16546 468
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 12256 18912 12308 18964
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 15016 12724 15068 12776
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 21272 12724 21324 12776
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 16304 12588 16356 12640
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 22008 12588 22060 12640
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 11888 12291 11940 12300
rect 11888 12257 11897 12291
rect 11897 12257 11931 12291
rect 11931 12257 11940 12291
rect 11888 12248 11940 12257
rect 12348 12248 12400 12300
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 12716 12248 12768 12300
rect 12992 12291 13044 12300
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 16764 12384 16816 12436
rect 19340 12384 19392 12436
rect 15016 12316 15068 12368
rect 17592 12359 17644 12368
rect 17592 12325 17604 12359
rect 17604 12325 17644 12359
rect 17592 12316 17644 12325
rect 17776 12316 17828 12368
rect 18052 12316 18104 12368
rect 14832 12248 14884 12300
rect 12532 12180 12584 12232
rect 8852 12112 8904 12164
rect 16764 12291 16816 12300
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 15568 12180 15620 12232
rect 19248 12248 19300 12300
rect 17132 12180 17184 12232
rect 10876 12044 10928 12096
rect 11612 12044 11664 12096
rect 12900 12044 12952 12096
rect 14372 12044 14424 12096
rect 14924 12087 14976 12096
rect 14924 12053 14933 12087
rect 14933 12053 14967 12087
rect 14967 12053 14976 12087
rect 14924 12044 14976 12053
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 17040 12044 17092 12096
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 17684 12044 17736 12096
rect 19432 12044 19484 12096
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 9128 11840 9180 11892
rect 11244 11772 11296 11824
rect 8668 11704 8720 11756
rect 11520 11840 11572 11892
rect 12440 11840 12492 11892
rect 12992 11840 13044 11892
rect 11428 11772 11480 11824
rect 12808 11772 12860 11824
rect 13912 11772 13964 11824
rect 10600 11679 10652 11688
rect 10600 11645 10618 11679
rect 10618 11645 10652 11679
rect 10600 11636 10652 11645
rect 10692 11636 10744 11688
rect 11612 11704 11664 11756
rect 8944 11568 8996 11620
rect 11980 11636 12032 11688
rect 11336 11568 11388 11620
rect 12532 11636 12584 11688
rect 14004 11636 14056 11688
rect 16764 11840 16816 11892
rect 17224 11840 17276 11892
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 20628 11840 20680 11892
rect 14832 11636 14884 11688
rect 15752 11636 15804 11688
rect 12256 11568 12308 11620
rect 13544 11568 13596 11620
rect 14372 11611 14424 11620
rect 14372 11577 14381 11611
rect 14381 11577 14415 11611
rect 14415 11577 14424 11611
rect 14372 11568 14424 11577
rect 17040 11636 17092 11688
rect 17316 11636 17368 11688
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 10140 11500 10192 11552
rect 10968 11500 11020 11552
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 12440 11500 12492 11552
rect 12716 11500 12768 11552
rect 16304 11500 16356 11552
rect 16488 11543 16540 11552
rect 16488 11509 16497 11543
rect 16497 11509 16531 11543
rect 16531 11509 16540 11543
rect 16488 11500 16540 11509
rect 17684 11772 17736 11824
rect 17776 11772 17828 11824
rect 19156 11772 19208 11824
rect 18420 11636 18472 11688
rect 17868 11568 17920 11620
rect 19064 11636 19116 11688
rect 19432 11679 19484 11688
rect 19432 11645 19466 11679
rect 19466 11645 19484 11679
rect 19432 11636 19484 11645
rect 21456 11636 21508 11688
rect 18052 11500 18104 11552
rect 18512 11500 18564 11552
rect 18880 11500 18932 11552
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 10600 11296 10652 11348
rect 10968 11296 11020 11348
rect 8576 11160 8628 11212
rect 9588 11203 9640 11212
rect 9588 11169 9597 11203
rect 9597 11169 9631 11203
rect 9631 11169 9640 11203
rect 9588 11160 9640 11169
rect 10048 11160 10100 11212
rect 9312 11092 9364 11144
rect 10876 11160 10928 11212
rect 11152 11296 11204 11348
rect 11520 11296 11572 11348
rect 11612 11296 11664 11348
rect 12532 11296 12584 11348
rect 14188 11296 14240 11348
rect 14924 11296 14976 11348
rect 11244 11201 11296 11212
rect 11244 11167 11253 11201
rect 11253 11167 11287 11201
rect 11287 11167 11296 11201
rect 11244 11160 11296 11167
rect 11428 11203 11480 11212
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 11980 11160 12032 11212
rect 12440 11160 12492 11212
rect 13544 11271 13596 11280
rect 13544 11237 13553 11271
rect 13553 11237 13587 11271
rect 13587 11237 13596 11271
rect 13544 11228 13596 11237
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 16212 11339 16264 11348
rect 16212 11305 16221 11339
rect 16221 11305 16255 11339
rect 16255 11305 16264 11339
rect 16212 11296 16264 11305
rect 16488 11296 16540 11348
rect 18236 11296 18288 11348
rect 16856 11160 16908 11212
rect 17132 11228 17184 11280
rect 9036 11024 9088 11076
rect 11152 11024 11204 11076
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 12992 11092 13044 11144
rect 16580 11092 16632 11144
rect 19064 11228 19116 11280
rect 19248 11271 19300 11280
rect 19248 11237 19282 11271
rect 19282 11237 19300 11271
rect 19248 11228 19300 11237
rect 17316 11160 17368 11212
rect 18420 11160 18472 11212
rect 11980 11024 12032 11076
rect 16764 11067 16816 11076
rect 16764 11033 16773 11067
rect 16773 11033 16807 11067
rect 16807 11033 16816 11067
rect 16764 11024 16816 11033
rect 18328 11024 18380 11076
rect 9680 10956 9732 11008
rect 11704 10999 11756 11008
rect 11704 10965 11713 10999
rect 11713 10965 11747 10999
rect 11747 10965 11756 10999
rect 11704 10956 11756 10965
rect 18604 10999 18656 11008
rect 18604 10965 18613 10999
rect 18613 10965 18647 10999
rect 18647 10965 18656 10999
rect 18604 10956 18656 10965
rect 28264 11024 28316 11076
rect 19340 10956 19392 11008
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 8484 10548 8536 10600
rect 9680 10752 9732 10804
rect 10140 10752 10192 10804
rect 11060 10752 11112 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 9680 10548 9732 10600
rect 8760 10480 8812 10532
rect 10140 10548 10192 10600
rect 11428 10684 11480 10736
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 7840 10412 7892 10464
rect 9404 10412 9456 10464
rect 9864 10412 9916 10464
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 10324 10412 10376 10464
rect 10784 10455 10836 10464
rect 10784 10421 10793 10455
rect 10793 10421 10827 10455
rect 10827 10421 10836 10455
rect 10784 10412 10836 10421
rect 11060 10523 11112 10532
rect 11060 10489 11069 10523
rect 11069 10489 11103 10523
rect 11103 10489 11112 10523
rect 11060 10480 11112 10489
rect 12900 10752 12952 10804
rect 13820 10727 13872 10736
rect 13820 10693 13829 10727
rect 13829 10693 13863 10727
rect 13863 10693 13872 10727
rect 13820 10684 13872 10693
rect 12992 10616 13044 10668
rect 12532 10548 12584 10600
rect 14004 10548 14056 10600
rect 14372 10548 14424 10600
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 18236 10795 18288 10804
rect 18236 10761 18245 10795
rect 18245 10761 18279 10795
rect 18279 10761 18288 10795
rect 18236 10752 18288 10761
rect 18696 10752 18748 10804
rect 20720 10752 20772 10804
rect 18512 10684 18564 10736
rect 19340 10616 19392 10668
rect 11520 10412 11572 10464
rect 13728 10480 13780 10532
rect 16580 10548 16632 10600
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 18604 10548 18656 10600
rect 18880 10548 18932 10600
rect 16212 10480 16264 10532
rect 19984 10548 20036 10600
rect 21732 10684 21784 10736
rect 21640 10548 21692 10600
rect 14280 10455 14332 10464
rect 14280 10421 14289 10455
rect 14289 10421 14323 10455
rect 14323 10421 14332 10455
rect 14280 10412 14332 10421
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 15108 10455 15160 10464
rect 15108 10421 15117 10455
rect 15117 10421 15151 10455
rect 15151 10421 15160 10455
rect 15108 10412 15160 10421
rect 22284 10480 22336 10532
rect 18972 10412 19024 10464
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 21180 10412 21232 10464
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 21548 10455 21600 10464
rect 21548 10421 21557 10455
rect 21557 10421 21591 10455
rect 21591 10421 21600 10455
rect 21548 10412 21600 10421
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 8116 10208 8168 10260
rect 10232 10208 10284 10260
rect 11060 10208 11112 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 12164 10208 12216 10260
rect 8484 10140 8536 10192
rect 10324 10140 10376 10192
rect 10876 10140 10928 10192
rect 11152 10140 11204 10192
rect 8392 10072 8444 10124
rect 9220 10072 9272 10124
rect 9496 10072 9548 10124
rect 8208 9936 8260 9988
rect 11796 10072 11848 10124
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12256 10115 12308 10124
rect 12256 10081 12265 10115
rect 12265 10081 12299 10115
rect 12299 10081 12308 10115
rect 12256 10072 12308 10081
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 14280 10208 14332 10260
rect 14832 10208 14884 10260
rect 13820 10140 13872 10192
rect 15108 10140 15160 10192
rect 16212 10208 16264 10260
rect 7932 9868 7984 9920
rect 9312 9936 9364 9988
rect 11520 9936 11572 9988
rect 12348 9936 12400 9988
rect 14096 10072 14148 10124
rect 17040 10208 17092 10260
rect 17868 10208 17920 10260
rect 14188 10004 14240 10056
rect 14372 10004 14424 10056
rect 14740 10004 14792 10056
rect 16948 10115 17000 10124
rect 16948 10081 16957 10115
rect 16957 10081 16991 10115
rect 16991 10081 17000 10115
rect 16948 10072 17000 10081
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 15200 9936 15252 9988
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 17224 9936 17276 9988
rect 9772 9868 9824 9920
rect 10140 9868 10192 9920
rect 11336 9868 11388 9920
rect 12716 9868 12768 9920
rect 13820 9868 13872 9920
rect 14004 9868 14056 9920
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 16488 9868 16540 9920
rect 16672 9868 16724 9920
rect 17316 9911 17368 9920
rect 17316 9877 17325 9911
rect 17325 9877 17359 9911
rect 17359 9877 17368 9911
rect 17316 9868 17368 9877
rect 17684 10115 17736 10124
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 18972 10072 19024 10124
rect 21272 10140 21324 10192
rect 21548 10208 21600 10260
rect 31668 10208 31720 10260
rect 19892 10072 19944 10124
rect 18420 9868 18472 9920
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 20260 9936 20312 9988
rect 21548 9936 21600 9988
rect 22192 10004 22244 10056
rect 22560 9936 22612 9988
rect 22008 9868 22060 9920
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 9404 9664 9456 9716
rect 9496 9707 9548 9716
rect 9496 9673 9505 9707
rect 9505 9673 9539 9707
rect 9539 9673 9548 9707
rect 9496 9664 9548 9673
rect 10784 9664 10836 9716
rect 13636 9664 13688 9716
rect 14556 9664 14608 9716
rect 8576 9596 8628 9648
rect 8668 9639 8720 9648
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 9128 9596 9180 9648
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 8852 9460 8904 9512
rect 10140 9596 10192 9648
rect 12532 9596 12584 9648
rect 13912 9596 13964 9648
rect 10232 9528 10284 9580
rect 11612 9528 11664 9580
rect 14280 9528 14332 9580
rect 9956 9503 10008 9512
rect 9956 9469 9971 9503
rect 9971 9469 10005 9503
rect 10005 9469 10008 9503
rect 9956 9460 10008 9469
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 10416 9503 10468 9512
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 10508 9503 10560 9512
rect 10508 9469 10517 9503
rect 10517 9469 10551 9503
rect 10551 9469 10560 9503
rect 10508 9460 10560 9469
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 11244 9503 11296 9512
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 11336 9503 11388 9512
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 16304 9596 16356 9648
rect 17224 9596 17276 9648
rect 19524 9639 19576 9648
rect 19524 9605 19533 9639
rect 19533 9605 19567 9639
rect 19567 9605 19576 9639
rect 19524 9596 19576 9605
rect 22100 9664 22152 9716
rect 22284 9707 22336 9716
rect 22284 9673 22293 9707
rect 22293 9673 22327 9707
rect 22327 9673 22336 9707
rect 22284 9664 22336 9673
rect 22376 9664 22428 9716
rect 28264 9596 28316 9648
rect 22192 9528 22244 9580
rect 10232 9392 10284 9444
rect 10876 9392 10928 9444
rect 19064 9460 19116 9512
rect 20720 9460 20772 9512
rect 21088 9503 21140 9512
rect 21088 9469 21097 9503
rect 21097 9469 21131 9503
rect 21131 9469 21140 9503
rect 21088 9460 21140 9469
rect 21456 9503 21508 9512
rect 21456 9469 21465 9503
rect 21465 9469 21499 9503
rect 21499 9469 21508 9503
rect 21456 9460 21508 9469
rect 21548 9503 21600 9512
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 21548 9460 21600 9469
rect 21640 9503 21692 9512
rect 21640 9469 21649 9503
rect 21649 9469 21683 9503
rect 21683 9469 21692 9503
rect 21640 9460 21692 9469
rect 21732 9460 21784 9512
rect 22008 9460 22060 9512
rect 22376 9503 22428 9512
rect 22376 9469 22385 9503
rect 22385 9469 22419 9503
rect 22419 9469 22428 9503
rect 22376 9460 22428 9469
rect 22560 9528 22612 9580
rect 12072 9392 12124 9444
rect 13360 9435 13412 9444
rect 13360 9401 13369 9435
rect 13369 9401 13403 9435
rect 13403 9401 13412 9435
rect 13360 9392 13412 9401
rect 13452 9392 13504 9444
rect 14004 9435 14056 9444
rect 14004 9401 14013 9435
rect 14013 9401 14047 9435
rect 14047 9401 14056 9435
rect 14004 9392 14056 9401
rect 18512 9392 18564 9444
rect 19708 9435 19760 9444
rect 19708 9401 19717 9435
rect 19717 9401 19751 9435
rect 19751 9401 19760 9435
rect 19708 9392 19760 9401
rect 20076 9435 20128 9444
rect 20076 9401 20085 9435
rect 20085 9401 20119 9435
rect 20119 9401 20128 9435
rect 20076 9392 20128 9401
rect 22100 9392 22152 9444
rect 7380 9324 7432 9376
rect 8484 9324 8536 9376
rect 9404 9324 9456 9376
rect 9496 9324 9548 9376
rect 10048 9324 10100 9376
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 15476 9324 15528 9376
rect 15660 9324 15712 9376
rect 16580 9324 16632 9376
rect 17684 9324 17736 9376
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 21180 9367 21232 9376
rect 21180 9333 21189 9367
rect 21189 9333 21223 9367
rect 21223 9333 21232 9367
rect 21180 9324 21232 9333
rect 21364 9324 21416 9376
rect 22560 9367 22612 9376
rect 22560 9333 22569 9367
rect 22569 9333 22603 9367
rect 22603 9333 22612 9367
rect 22560 9324 22612 9333
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 7840 9120 7892 9172
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 8300 9120 8352 9172
rect 8760 9120 8812 9172
rect 8944 9163 8996 9172
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 9496 9120 9548 9172
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 7932 9027 7984 9036
rect 7932 8993 7941 9027
rect 7941 8993 7975 9027
rect 7975 8993 7984 9027
rect 7932 8984 7984 8993
rect 8024 8984 8076 9036
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 7932 8848 7984 8900
rect 9588 9052 9640 9104
rect 10048 9120 10100 9172
rect 10508 9120 10560 9172
rect 10968 9120 11020 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 13360 9120 13412 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 17132 9120 17184 9172
rect 9312 8984 9364 9036
rect 11244 9052 11296 9104
rect 11704 9052 11756 9104
rect 13912 9052 13964 9104
rect 15660 9052 15712 9104
rect 17960 9052 18012 9104
rect 19340 9120 19392 9172
rect 21088 9120 21140 9172
rect 21180 9120 21232 9172
rect 21272 9120 21324 9172
rect 22560 9120 22612 9172
rect 10416 8916 10468 8968
rect 11796 8916 11848 8968
rect 12624 8984 12676 9036
rect 13544 8984 13596 9036
rect 13820 8984 13872 9036
rect 12532 8916 12584 8968
rect 13912 8916 13964 8968
rect 16948 8984 17000 9036
rect 17040 8916 17092 8968
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 18788 8984 18840 9036
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 12992 8848 13044 8900
rect 14648 8848 14700 8900
rect 16580 8848 16632 8900
rect 9864 8780 9916 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 12440 8780 12492 8832
rect 13360 8780 13412 8832
rect 15568 8780 15620 8832
rect 18696 8780 18748 8832
rect 22284 9052 22336 9104
rect 22376 9052 22428 9104
rect 22008 8984 22060 9036
rect 28264 8848 28316 8900
rect 20812 8823 20864 8832
rect 20812 8789 20821 8823
rect 20821 8789 20855 8823
rect 20855 8789 20864 8823
rect 20812 8780 20864 8789
rect 20996 8780 21048 8832
rect 22008 8780 22060 8832
rect 22192 8823 22244 8832
rect 22192 8789 22201 8823
rect 22201 8789 22235 8823
rect 22235 8789 22244 8823
rect 22192 8780 22244 8789
rect 22468 8823 22520 8832
rect 22468 8789 22477 8823
rect 22477 8789 22511 8823
rect 22511 8789 22520 8823
rect 22468 8780 22520 8789
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 8392 8576 8444 8628
rect 9220 8576 9272 8628
rect 10692 8576 10744 8628
rect 11060 8576 11112 8628
rect 12532 8576 12584 8628
rect 13452 8576 13504 8628
rect 14280 8576 14332 8628
rect 8576 8508 8628 8560
rect 8668 8508 8720 8560
rect 11152 8508 11204 8560
rect 8484 8372 8536 8424
rect 8944 8440 8996 8492
rect 11244 8440 11296 8492
rect 9956 8372 10008 8424
rect 13176 8508 13228 8560
rect 13360 8508 13412 8560
rect 9864 8347 9916 8356
rect 9864 8313 9873 8347
rect 9873 8313 9907 8347
rect 9907 8313 9916 8347
rect 9864 8304 9916 8313
rect 10232 8347 10284 8356
rect 10232 8313 10241 8347
rect 10241 8313 10275 8347
rect 10275 8313 10284 8347
rect 10232 8304 10284 8313
rect 10600 8347 10652 8356
rect 10600 8313 10609 8347
rect 10609 8313 10643 8347
rect 10643 8313 10652 8347
rect 10600 8304 10652 8313
rect 11520 8347 11572 8356
rect 11520 8313 11529 8347
rect 11529 8313 11563 8347
rect 11563 8313 11572 8347
rect 11520 8304 11572 8313
rect 8392 8236 8444 8288
rect 10692 8279 10744 8288
rect 10692 8245 10701 8279
rect 10701 8245 10735 8279
rect 10735 8245 10744 8279
rect 10692 8236 10744 8245
rect 10784 8236 10836 8288
rect 11336 8236 11388 8288
rect 12348 8372 12400 8424
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 12716 8372 12768 8424
rect 11796 8347 11848 8356
rect 11796 8313 11805 8347
rect 11805 8313 11839 8347
rect 11839 8313 11848 8347
rect 11796 8304 11848 8313
rect 11888 8304 11940 8356
rect 12716 8236 12768 8288
rect 12900 8440 12952 8492
rect 13084 8409 13136 8424
rect 13084 8375 13093 8409
rect 13093 8375 13127 8409
rect 13127 8375 13136 8409
rect 13084 8372 13136 8375
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13636 8372 13688 8424
rect 15200 8508 15252 8560
rect 16948 8440 17000 8492
rect 12992 8347 13044 8356
rect 12992 8313 13001 8347
rect 13001 8313 13035 8347
rect 13035 8313 13044 8347
rect 12992 8304 13044 8313
rect 15476 8347 15528 8356
rect 15476 8313 15485 8347
rect 15485 8313 15519 8347
rect 15519 8313 15528 8347
rect 15476 8304 15528 8313
rect 15660 8304 15712 8356
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17224 8372 17276 8424
rect 18328 8576 18380 8628
rect 17960 8372 18012 8424
rect 18788 8551 18840 8560
rect 18788 8517 18797 8551
rect 18797 8517 18831 8551
rect 18831 8517 18840 8551
rect 18788 8508 18840 8517
rect 22376 8508 22428 8560
rect 14556 8236 14608 8288
rect 15200 8236 15252 8288
rect 15568 8236 15620 8288
rect 16212 8236 16264 8288
rect 17040 8279 17092 8288
rect 17040 8245 17049 8279
rect 17049 8245 17083 8279
rect 17083 8245 17092 8279
rect 17040 8236 17092 8245
rect 17868 8347 17920 8356
rect 17868 8313 17877 8347
rect 17877 8313 17911 8347
rect 17911 8313 17920 8347
rect 17868 8304 17920 8313
rect 18328 8304 18380 8356
rect 18604 8304 18656 8356
rect 21364 8415 21416 8424
rect 21364 8381 21373 8415
rect 21373 8381 21407 8415
rect 21407 8381 21416 8415
rect 21364 8372 21416 8381
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 19984 8304 20036 8356
rect 21548 8347 21600 8356
rect 21548 8313 21557 8347
rect 21557 8313 21591 8347
rect 21591 8313 21600 8347
rect 21548 8304 21600 8313
rect 18144 8236 18196 8288
rect 18696 8236 18748 8288
rect 31668 8440 31720 8492
rect 21732 8415 21784 8424
rect 21732 8381 21741 8415
rect 21741 8381 21775 8415
rect 21775 8381 21784 8415
rect 21732 8372 21784 8381
rect 22008 8415 22060 8424
rect 22008 8381 22017 8415
rect 22017 8381 22051 8415
rect 22051 8381 22060 8415
rect 22008 8372 22060 8381
rect 21824 8279 21876 8288
rect 21824 8245 21833 8279
rect 21833 8245 21867 8279
rect 21867 8245 21876 8279
rect 21824 8236 21876 8245
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 8484 8032 8536 8084
rect 10600 8075 10652 8084
rect 10600 8041 10609 8075
rect 10609 8041 10643 8075
rect 10643 8041 10652 8075
rect 10600 8032 10652 8041
rect 12532 8032 12584 8084
rect 14188 8032 14240 8084
rect 20812 8032 20864 8084
rect 8576 7964 8628 8016
rect 11244 7964 11296 8016
rect 8668 7896 8720 7948
rect 8852 7896 8904 7948
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 9036 7896 9088 7905
rect 9220 7939 9272 7948
rect 9220 7905 9229 7939
rect 9229 7905 9263 7939
rect 9263 7905 9272 7939
rect 9220 7896 9272 7905
rect 10416 7896 10468 7948
rect 12348 7964 12400 8016
rect 12716 7964 12768 8016
rect 13544 7964 13596 8016
rect 13176 7828 13228 7880
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 11612 7760 11664 7812
rect 9864 7692 9916 7744
rect 10968 7692 11020 7744
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 12440 7760 12492 7812
rect 12716 7760 12768 7812
rect 13360 7939 13412 7948
rect 13360 7905 13369 7939
rect 13369 7905 13403 7939
rect 13403 7905 13412 7939
rect 13360 7896 13412 7905
rect 13820 7896 13872 7948
rect 14096 7896 14148 7948
rect 14280 7896 14332 7948
rect 14464 7896 14516 7948
rect 14740 7896 14792 7948
rect 16212 7964 16264 8016
rect 17040 7964 17092 8016
rect 13728 7692 13780 7744
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 15384 7692 15436 7744
rect 16580 7896 16632 7948
rect 17132 7939 17184 7948
rect 17132 7905 17141 7939
rect 17141 7905 17175 7939
rect 17175 7905 17184 7939
rect 17132 7896 17184 7905
rect 17684 7896 17736 7948
rect 18420 7964 18472 8016
rect 21824 7964 21876 8016
rect 18144 7896 18196 7948
rect 19432 7896 19484 7948
rect 16396 7828 16448 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 16672 7760 16724 7812
rect 20996 7896 21048 7948
rect 21732 7828 21784 7880
rect 17408 7692 17460 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 21272 7760 21324 7812
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 7656 7488 7708 7540
rect 10416 7488 10468 7540
rect 9036 7352 9088 7404
rect 8668 7284 8720 7336
rect 10140 7352 10192 7404
rect 10600 7352 10652 7404
rect 12624 7488 12676 7540
rect 12716 7488 12768 7540
rect 13176 7488 13228 7540
rect 13360 7488 13412 7540
rect 13728 7488 13780 7540
rect 14464 7488 14516 7540
rect 15384 7488 15436 7540
rect 16212 7488 16264 7540
rect 16396 7488 16448 7540
rect 17684 7488 17736 7540
rect 12348 7420 12400 7472
rect 12532 7420 12584 7472
rect 18420 7488 18472 7540
rect 19248 7488 19300 7540
rect 20076 7488 20128 7540
rect 20260 7488 20312 7540
rect 22008 7488 22060 7540
rect 9036 7259 9088 7268
rect 9036 7225 9045 7259
rect 9045 7225 9079 7259
rect 9079 7225 9088 7259
rect 9036 7216 9088 7225
rect 10784 7216 10836 7268
rect 11244 7216 11296 7268
rect 12348 7216 12400 7268
rect 12900 7284 12952 7336
rect 13084 7284 13136 7336
rect 16580 7352 16632 7404
rect 18604 7352 18656 7404
rect 19432 7420 19484 7472
rect 21364 7420 21416 7472
rect 19616 7352 19668 7404
rect 14004 7284 14056 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 12992 7259 13044 7268
rect 12992 7225 13001 7259
rect 13001 7225 13035 7259
rect 13035 7225 13044 7259
rect 12992 7216 13044 7225
rect 13544 7216 13596 7268
rect 10508 7148 10560 7200
rect 12256 7148 12308 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 14096 7259 14148 7268
rect 14096 7225 14105 7259
rect 14105 7225 14139 7259
rect 14139 7225 14148 7259
rect 14096 7216 14148 7225
rect 15292 7216 15344 7268
rect 15476 7259 15528 7268
rect 15476 7225 15510 7259
rect 15510 7225 15528 7259
rect 15476 7216 15528 7225
rect 16948 7216 17000 7268
rect 18972 7284 19024 7336
rect 19340 7284 19392 7336
rect 20076 7352 20128 7404
rect 14464 7148 14516 7200
rect 14740 7148 14792 7200
rect 15384 7148 15436 7200
rect 16580 7191 16632 7200
rect 16580 7157 16589 7191
rect 16589 7157 16623 7191
rect 16623 7157 16632 7191
rect 16580 7148 16632 7157
rect 17040 7148 17092 7200
rect 20076 7216 20128 7268
rect 18880 7191 18932 7200
rect 18880 7157 18889 7191
rect 18889 7157 18923 7191
rect 18923 7157 18932 7191
rect 18880 7148 18932 7157
rect 19340 7191 19392 7200
rect 19340 7157 19349 7191
rect 19349 7157 19383 7191
rect 19383 7157 19392 7191
rect 19340 7148 19392 7157
rect 19432 7148 19484 7200
rect 19892 7148 19944 7200
rect 20352 7327 20404 7336
rect 20352 7293 20361 7327
rect 20361 7293 20395 7327
rect 20395 7293 20404 7327
rect 20352 7284 20404 7293
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 7564 6944 7616 6996
rect 7932 6944 7984 6996
rect 8024 6808 8076 6860
rect 9036 6944 9088 6996
rect 10508 6944 10560 6996
rect 11336 6944 11388 6996
rect 11704 6944 11756 6996
rect 9956 6808 10008 6860
rect 10232 6808 10284 6860
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 11060 6808 11112 6860
rect 9404 6604 9456 6656
rect 11704 6808 11756 6860
rect 13820 6944 13872 6996
rect 16396 6944 16448 6996
rect 17040 6944 17092 6996
rect 18144 6944 18196 6996
rect 18696 6987 18748 6996
rect 18696 6953 18705 6987
rect 18705 6953 18739 6987
rect 18739 6953 18748 6987
rect 18696 6944 18748 6953
rect 18972 6987 19024 6996
rect 18972 6953 18981 6987
rect 18981 6953 19015 6987
rect 19015 6953 19024 6987
rect 18972 6944 19024 6953
rect 19340 6944 19392 6996
rect 13084 6876 13136 6928
rect 14740 6876 14792 6928
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 12900 6851 12952 6860
rect 12900 6817 12934 6851
rect 12934 6817 12952 6851
rect 12900 6808 12952 6817
rect 14464 6851 14516 6860
rect 14464 6817 14473 6851
rect 14473 6817 14507 6851
rect 14507 6817 14516 6851
rect 14464 6808 14516 6817
rect 11428 6672 11480 6724
rect 11520 6672 11572 6724
rect 12256 6740 12308 6792
rect 13728 6740 13780 6792
rect 14648 6808 14700 6860
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 15200 6740 15252 6792
rect 15476 6740 15528 6792
rect 16580 6876 16632 6928
rect 17500 6808 17552 6860
rect 17684 6808 17736 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 14096 6672 14148 6724
rect 17960 6740 18012 6792
rect 18328 6740 18380 6792
rect 16304 6672 16356 6724
rect 16856 6715 16908 6724
rect 16856 6681 16865 6715
rect 16865 6681 16899 6715
rect 16899 6681 16908 6715
rect 16856 6672 16908 6681
rect 19248 6808 19300 6860
rect 19616 6944 19668 6996
rect 20076 6919 20128 6928
rect 20076 6885 20085 6919
rect 20085 6885 20119 6919
rect 20119 6885 20128 6919
rect 20076 6876 20128 6885
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 19984 6808 20036 6860
rect 20628 6944 20680 6996
rect 20996 6944 21048 6996
rect 18788 6672 18840 6724
rect 22468 6672 22520 6724
rect 15568 6604 15620 6656
rect 16396 6647 16448 6656
rect 16396 6613 16405 6647
rect 16405 6613 16439 6647
rect 16439 6613 16448 6647
rect 16396 6604 16448 6613
rect 21456 6604 21508 6656
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 10508 6400 10560 6452
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 11428 6400 11480 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 12348 6400 12400 6452
rect 12440 6400 12492 6452
rect 13728 6400 13780 6452
rect 14556 6400 14608 6452
rect 15016 6400 15068 6452
rect 16396 6400 16448 6452
rect 16948 6400 17000 6452
rect 17132 6400 17184 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18788 6400 18840 6452
rect 19432 6400 19484 6452
rect 11060 6375 11112 6384
rect 11060 6341 11069 6375
rect 11069 6341 11103 6375
rect 11103 6341 11112 6375
rect 11060 6332 11112 6341
rect 8944 6196 8996 6248
rect 9864 6196 9916 6248
rect 10140 6196 10192 6248
rect 12624 6332 12676 6384
rect 12716 6375 12768 6384
rect 12716 6341 12725 6375
rect 12725 6341 12759 6375
rect 12759 6341 12768 6375
rect 12716 6332 12768 6341
rect 13084 6332 13136 6384
rect 13268 6332 13320 6384
rect 15292 6375 15344 6384
rect 15292 6341 15301 6375
rect 15301 6341 15335 6375
rect 15335 6341 15344 6375
rect 15292 6332 15344 6341
rect 11244 6264 11296 6316
rect 11336 6264 11388 6316
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 12164 6196 12216 6248
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 12072 6128 12124 6180
rect 12716 6128 12768 6180
rect 13820 6196 13872 6248
rect 14004 6196 14056 6248
rect 15568 6264 15620 6316
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 16212 6196 16264 6248
rect 16764 6196 16816 6248
rect 17500 6264 17552 6316
rect 18052 6264 18104 6316
rect 18144 6264 18196 6316
rect 14096 6128 14148 6180
rect 14464 6128 14516 6180
rect 21548 6196 21600 6248
rect 18328 6128 18380 6180
rect 20904 6128 20956 6180
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 9680 5856 9732 5908
rect 9772 5856 9824 5908
rect 12072 5856 12124 5908
rect 12716 5856 12768 5908
rect 12992 5856 13044 5908
rect 14004 5856 14056 5908
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 11152 5788 11204 5840
rect 11704 5652 11756 5704
rect 13912 5763 13964 5772
rect 13912 5729 13921 5763
rect 13921 5729 13955 5763
rect 13955 5729 13964 5763
rect 13912 5720 13964 5729
rect 12440 5584 12492 5636
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 11060 5312 11112 5364
rect 12624 5355 12676 5364
rect 12624 5321 12633 5355
rect 12633 5321 12667 5355
rect 12667 5321 12676 5355
rect 12624 5312 12676 5321
rect 12900 5312 12952 5364
rect 12532 5151 12584 5160
rect 12532 5117 12541 5151
rect 12541 5117 12575 5151
rect 12575 5117 12584 5151
rect 12532 5108 12584 5117
rect 12716 5108 12768 5160
rect 12992 5108 13044 5160
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 14372 4088 14424 4140
rect 18052 4088 18104 4140
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 12348 3476 12400 3528
rect 14096 3476 14148 3528
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
rect 16028 416 16080 468
rect 16488 416 16540 468
<< metal2 >>
rect 12254 19600 12310 20000
rect 13542 19600 13598 20000
rect 14186 19600 14242 20000
rect 15474 19600 15530 20000
rect 16118 19600 16174 20000
rect 17406 19600 17462 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 19338 19600 19394 20000
rect 19536 19638 19932 19666
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 12268 18970 12296 19600
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 4250 18459 4558 18468
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 4250 15260 4558 15269
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 11888 12300 11940 12306
rect 11808 12260 11888 12288
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 9042 7420 9318
rect 7852 9178 7880 10406
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 8102 10299 8410 10308
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7944 9178 7972 9862
rect 8128 9586 8156 10202
rect 8496 10198 8524 10542
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8404 10033 8432 10066
rect 8390 10024 8446 10033
rect 8208 9988 8260 9994
rect 8390 9959 8446 9968
rect 8208 9930 8260 9936
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8220 9518 8248 9930
rect 8588 9654 8616 11154
rect 8680 9654 8708 11698
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 8300 9172 8352 9178
rect 8496 9160 8524 9318
rect 8772 9178 8800 10474
rect 8864 9518 8892 12106
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8956 9178 8984 11562
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8352 9132 8524 9160
rect 8760 9172 8812 9178
rect 8300 9114 8352 9120
rect 8760 9114 8812 9120
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 7930 9072 7986 9081
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7656 9036 7708 9042
rect 7930 9007 7932 9016
rect 7656 8978 7708 8984
rect 7984 9007 7986 9016
rect 8024 9036 8076 9042
rect 7932 8978 7984 8984
rect 8024 8978 8076 8984
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 7576 7002 7604 8910
rect 7668 7546 7696 8978
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7944 7002 7972 8842
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 8036 6866 8064 8978
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8404 8634 8432 8774
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8680 8566 8708 8774
rect 8576 8560 8628 8566
rect 8390 8528 8446 8537
rect 8576 8502 8628 8508
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8390 8463 8446 8472
rect 8404 8294 8432 8463
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 8496 8090 8524 8366
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8588 8022 8616 8502
rect 8772 8294 8800 9114
rect 9048 9081 9076 11018
rect 9140 9654 9168 11834
rect 10600 11688 10652 11694
rect 9954 11656 10010 11665
rect 10600 11630 10652 11636
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 9954 11591 10010 11600
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9324 10606 9352 11086
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9310 10160 9366 10169
rect 9220 10124 9272 10130
rect 9310 10095 9366 10104
rect 9220 10066 9272 10072
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9034 9072 9090 9081
rect 9034 9007 9090 9016
rect 8942 8936 8998 8945
rect 8942 8871 8998 8880
rect 8956 8498 8984 8871
rect 9232 8634 9260 10066
rect 9324 9994 9352 10095
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9324 9042 9352 9930
rect 9416 9722 9444 10406
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9508 10033 9536 10066
rect 9494 10024 9550 10033
rect 9494 9959 9550 9968
rect 9494 9752 9550 9761
rect 9404 9716 9456 9722
rect 9494 9687 9496 9696
rect 9404 9658 9456 9664
rect 9548 9687 9550 9696
rect 9496 9658 9548 9664
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9324 8294 9352 8978
rect 8772 8266 8892 8294
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8864 7954 8892 8266
rect 9232 8266 9352 8294
rect 9232 7954 9260 8266
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 8680 7342 8708 7890
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 8956 6254 8984 7686
rect 9048 7410 9076 7890
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9048 7002 9076 7210
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9416 6662 9444 9318
rect 9508 9178 9536 9318
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9600 9110 9628 11154
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10810 9720 10950
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 9692 5914 9720 10542
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 5914 9812 9862
rect 9876 8838 9904 10406
rect 9968 9518 9996 11591
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10588 10088 11154
rect 10152 10810 10180 11494
rect 10612 11354 10640 11630
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10140 10600 10192 10606
rect 10060 10560 10140 10588
rect 10140 10542 10192 10548
rect 10152 9926 10180 10542
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10244 10266 10272 10406
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10336 10198 10364 10406
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 10152 9654 10180 9862
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 9956 9512 10008 9518
rect 10140 9512 10192 9518
rect 9956 9454 10008 9460
rect 10138 9480 10140 9489
rect 10192 9480 10194 9489
rect 10244 9450 10272 9522
rect 10138 9415 10194 9424
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 9178 10088 9318
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9876 7993 9904 8298
rect 9862 7984 9918 7993
rect 9862 7919 9918 7928
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 6254 9904 7686
rect 9968 6866 9996 8366
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 10152 6254 10180 7346
rect 10244 6866 10272 8298
rect 10336 8294 10364 10134
rect 10598 9752 10654 9761
rect 10598 9687 10654 9696
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10428 8974 10456 9454
rect 10520 9178 10548 9454
rect 10612 9382 10640 9687
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10704 8634 10732 11630
rect 10888 11218 10916 12038
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11244 11824 11296 11830
rect 11428 11824 11480 11830
rect 11296 11784 11428 11812
rect 11244 11766 11296 11772
rect 11428 11766 11480 11772
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10980 11354 11008 11494
rect 11242 11384 11298 11393
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11152 11348 11204 11354
rect 11242 11319 11298 11328
rect 11152 11290 11204 11296
rect 11164 11257 11192 11290
rect 11150 11248 11206 11257
rect 10876 11212 10928 11218
rect 11256 11218 11284 11319
rect 11150 11183 11206 11192
rect 11244 11212 11296 11218
rect 10876 11154 10928 11160
rect 11244 11154 11296 11160
rect 11348 11098 11376 11562
rect 11532 11354 11560 11834
rect 11624 11762 11652 12038
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11610 11656 11666 11665
rect 11610 11591 11666 11600
rect 11624 11354 11652 11591
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11393 11744 11494
rect 11702 11384 11758 11393
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11612 11348 11664 11354
rect 11702 11319 11758 11328
rect 11612 11290 11664 11296
rect 11426 11248 11482 11257
rect 11426 11183 11428 11192
rect 11480 11183 11482 11192
rect 11520 11212 11572 11218
rect 11428 11154 11480 11160
rect 11520 11154 11572 11160
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11256 11070 11376 11098
rect 11058 10840 11114 10849
rect 11058 10775 11060 10784
rect 11112 10775 11114 10784
rect 11060 10746 11112 10752
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 9722 10824 10406
rect 10888 10198 10916 10542
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10266 11100 10474
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11164 10198 11192 11018
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11256 9908 11284 11070
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 11334 10296 11390 10305
rect 11334 10231 11336 10240
rect 11388 10231 11390 10240
rect 11336 10202 11388 10208
rect 11336 9920 11388 9926
rect 11256 9880 11336 9908
rect 11336 9862 11388 9868
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 10968 9512 11020 9518
rect 10874 9480 10930 9489
rect 10968 9454 11020 9460
rect 10874 9415 10876 9424
rect 10928 9415 10930 9424
rect 10876 9386 10928 9392
rect 10980 9178 11008 9454
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11164 8838 11192 9551
rect 11348 9518 11376 9862
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11256 9110 11284 9454
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10336 8266 10548 8294
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10428 7546 10456 7890
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10520 7206 10548 8266
rect 10612 8090 10640 8298
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10704 7585 10732 8230
rect 10690 7576 10746 7585
rect 10690 7511 10746 7520
rect 10600 7404 10652 7410
rect 10796 7392 10824 8230
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10652 7364 10824 7392
rect 10600 7346 10652 7352
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 7002 10548 7142
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10520 6458 10548 6802
rect 10796 6458 10824 7210
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 10322 3768 10378 3777
rect 10322 3703 10378 3712
rect 9678 3496 9734 3505
rect 9678 3431 9734 3440
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 9692 400 9720 3431
rect 10336 400 10364 3703
rect 10980 400 11008 7686
rect 11072 6866 11100 8570
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11072 5370 11100 6326
rect 11164 5846 11192 8502
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11256 8022 11284 8434
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11256 7274 11284 7958
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11348 7154 11376 8230
rect 11256 7126 11376 7154
rect 11256 6322 11284 7126
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11348 6322 11376 6938
rect 11440 6905 11468 10678
rect 11532 10470 11560 11154
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 9994 11560 10406
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11624 9586 11652 11154
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10810 11744 10950
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11808 10690 11836 12260
rect 11888 12242 11940 12248
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11992 11218 12020 11630
rect 12256 11620 12308 11626
rect 12360 11608 12388 12242
rect 12452 11898 12480 12242
rect 12544 12238 12572 18566
rect 13556 16574 13584 19600
rect 13556 16546 13860 16574
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12544 11694 12572 12174
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12308 11580 12388 11608
rect 12256 11562 12308 11568
rect 12440 11552 12492 11558
rect 12360 11512 12440 11540
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11992 11082 12020 11154
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11955 10843 12263 10852
rect 11716 10662 11836 10690
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11716 9110 11744 10662
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12176 10130 12204 10202
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12256 10124 12308 10130
rect 12360 10112 12388 11512
rect 12440 11494 12492 11500
rect 12544 11354 12572 11630
rect 12728 11558 12756 12242
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12308 10084 12388 10112
rect 12256 10066 12308 10072
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11808 8974 11836 10066
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 9178 12112 9386
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11808 8650 11836 8910
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 11808 8622 11928 8650
rect 11900 8362 11928 8622
rect 12360 8430 12388 9930
rect 12452 8838 12480 11154
rect 12820 11150 12848 11766
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12912 10810 12940 12038
rect 13004 11898 13032 12242
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13556 11286 13584 11562
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13004 10674 13032 11086
rect 13832 10742 13860 16546
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 11830 13952 12582
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 14016 10606 14044 11630
rect 14200 11354 14228 19600
rect 15488 16574 15516 19600
rect 16132 19258 16160 19600
rect 16132 19230 16252 19258
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 15488 16546 15700 16574
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15028 12374 15056 12718
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14372 12096 14424 12102
rect 14844 12073 14872 12242
rect 15580 12238 15608 12582
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 14924 12096 14976 12102
rect 14372 12038 14424 12044
rect 14830 12064 14886 12073
rect 14384 11626 14412 12038
rect 14924 12038 14976 12044
rect 14830 11999 14886 12008
rect 14844 11694 14872 11999
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14936 11354 14964 12038
rect 15672 11354 15700 16546
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15764 11694 15792 12038
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15807 11452 16115 11461
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15807 11387 16115 11396
rect 16224 11354 16252 19230
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 11558 16344 12582
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16776 12306 16804 12378
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11898 16804 12242
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17040 12096 17092 12102
rect 17144 12073 17172 12174
rect 17224 12096 17276 12102
rect 17040 12038 17092 12044
rect 17130 12064 17186 12073
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 17052 11694 17080 12038
rect 17224 12038 17276 12044
rect 17130 11999 17186 12008
rect 17236 11898 17264 12038
rect 17328 11898 17356 12718
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 12544 10169 12572 10542
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13740 10266 13768 10474
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14292 10266 14320 10406
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 13820 10192 13872 10198
rect 12530 10160 12586 10169
rect 13820 10134 13872 10140
rect 12530 10095 12586 10104
rect 12544 9654 12572 10095
rect 13832 9926 13860 10134
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14002 10024 14058 10033
rect 14002 9959 14058 9968
rect 14016 9926 14044 9959
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 12532 9648 12584 9654
rect 12584 9608 12664 9636
rect 12532 9590 12584 9596
rect 12636 9042 12664 9608
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11426 6896 11482 6905
rect 11426 6831 11482 6840
rect 11532 6730 11560 8298
rect 11808 7857 11836 8298
rect 11794 7848 11850 7857
rect 11612 7812 11664 7818
rect 11794 7783 11850 7792
rect 11612 7754 11664 7760
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11440 6458 11468 6666
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11624 400 11652 7754
rect 11704 7744 11756 7750
rect 11900 7698 11928 8298
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 11704 7686 11756 7692
rect 11716 7002 11744 7686
rect 11808 7670 11928 7698
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11716 5710 11744 6802
rect 11808 6236 11836 7670
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 12360 7478 12388 7958
rect 12452 7818 12480 8774
rect 12544 8634 12572 8910
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12544 8090 12572 8366
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12348 7472 12400 7478
rect 12162 7440 12218 7449
rect 12348 7414 12400 7420
rect 12162 7375 12218 7384
rect 12176 6866 12204 7375
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12268 6798 12296 7142
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11955 6491 12263 6500
rect 12360 6458 12388 7210
rect 12452 6458 12480 7754
rect 12636 7546 12664 8978
rect 12728 8430 12756 9862
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13372 9178 13400 9386
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12806 8528 12862 8537
rect 12806 8463 12862 8472
rect 12900 8492 12952 8498
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 8022 12756 8230
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 7546 12756 7754
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 11900 6361 11928 6394
rect 11886 6352 11942 6361
rect 12360 6338 12388 6394
rect 12360 6310 12480 6338
rect 11886 6287 11942 6296
rect 11980 6248 12032 6254
rect 11808 6208 11980 6236
rect 11980 6190 12032 6196
rect 12164 6248 12216 6254
rect 12348 6248 12400 6254
rect 12216 6208 12348 6236
rect 12164 6190 12216 6196
rect 12348 6190 12400 6196
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12084 5914 12112 6122
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 12452 5642 12480 6310
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 12544 5166 12572 7414
rect 12636 6866 12664 7482
rect 12820 7290 12848 8463
rect 12900 8434 12952 8440
rect 12912 7342 12940 8434
rect 13004 8362 13032 8842
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8566 13400 8774
rect 13464 8634 13492 9386
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13176 8560 13228 8566
rect 13082 8528 13138 8537
rect 13176 8502 13228 8508
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13082 8463 13138 8472
rect 13096 8430 13124 8463
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 13188 7970 13216 8502
rect 13556 8498 13584 8978
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13556 8022 13584 8434
rect 13648 8430 13676 9658
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13924 9110 13952 9590
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13636 8424 13688 8430
rect 13832 8401 13860 8978
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13636 8366 13688 8372
rect 13818 8392 13874 8401
rect 13818 8327 13874 8336
rect 13544 8016 13596 8022
rect 13188 7942 13308 7970
rect 13544 7958 13596 7964
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 7546 13216 7822
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 12728 7262 12848 7290
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12992 7268 13044 7274
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12728 6390 12756 7262
rect 12992 7210 13044 7216
rect 12900 7200 12952 7206
rect 12820 7160 12900 7188
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12636 5370 12664 6326
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12728 5914 12756 6122
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12728 5166 12756 5850
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 12360 898 12388 3470
rect 12820 2774 12848 7160
rect 12900 7142 12952 7148
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 5370 12940 6802
rect 13004 5914 13032 7210
rect 13096 6934 13124 7278
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 13096 6390 13124 6870
rect 13280 6390 13308 7942
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13372 7546 13400 7890
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13740 7546 13768 7686
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 13004 5166 13032 5510
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12820 2746 12940 2774
rect 12268 870 12388 898
rect 12268 400 12296 870
rect 12912 400 12940 2746
rect 13556 400 13584 7210
rect 13832 7002 13860 7890
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6458 13768 6734
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13740 6236 13768 6394
rect 13820 6248 13872 6254
rect 13740 6208 13820 6236
rect 13820 6190 13872 6196
rect 13924 5778 13952 8910
rect 14016 7426 14044 9386
rect 14108 7954 14136 10066
rect 14384 10062 14412 10542
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14200 8090 14228 9998
rect 14568 9722 14596 10406
rect 14844 10266 14872 10406
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 15120 10198 15148 10406
rect 15807 10364 16115 10373
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 16224 10266 16252 10474
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 16316 10062 16344 11494
rect 16500 11354 16528 11494
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 17132 11280 17184 11286
rect 17184 11228 17264 11234
rect 17132 11222 17264 11228
rect 16856 11212 16908 11218
rect 17144 11206 17264 11222
rect 17328 11218 17356 11630
rect 17420 11506 17448 19600
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12434 17540 12582
rect 17512 12406 17632 12434
rect 17604 12374 17632 12406
rect 18064 12374 18092 19600
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17696 11830 17724 12038
rect 17788 11830 17816 12310
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17500 11688 17552 11694
rect 17788 11676 17816 11766
rect 17552 11648 17816 11676
rect 18420 11688 18472 11694
rect 17500 11630 17552 11636
rect 18420 11630 18472 11636
rect 17868 11620 17920 11626
rect 17788 11580 17868 11608
rect 17420 11478 17540 11506
rect 16856 11154 16908 11160
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16592 10606 16620 11086
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14292 8634 14320 9522
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14462 8120 14518 8129
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14292 8078 14462 8106
rect 14292 7954 14320 8078
rect 14462 8055 14518 8064
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7562 14136 7686
rect 14108 7534 14412 7562
rect 14476 7546 14504 7890
rect 14016 7398 14228 7426
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 6254 14044 7278
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 6730 14136 7210
rect 14096 6724 14148 6730
rect 14096 6666 14148 6672
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5914 14044 6054
rect 14108 5914 14136 6122
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 14200 4162 14228 7398
rect 14108 4134 14228 4162
rect 14384 4146 14412 7534
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14476 7206 14504 7482
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14476 6186 14504 6802
rect 14568 6458 14596 8230
rect 14660 6866 14688 8842
rect 14752 7954 14780 9998
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 6934 14780 7142
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14372 4140 14424 4146
rect 14108 3534 14136 4134
rect 14372 4082 14424 4088
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14108 462 14228 490
rect 9678 0 9734 400
rect 10322 0 10378 400
rect 10966 0 11022 400
rect 11610 0 11666 400
rect 12254 0 12310 400
rect 12898 0 12954 400
rect 13542 0 13598 400
rect 14108 377 14136 462
rect 14200 400 14228 462
rect 14844 400 14872 9862
rect 15212 8566 15240 9930
rect 16316 9654 16344 9998
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15488 9178 15516 9318
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15672 9110 15700 9318
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15474 8392 15530 8401
rect 15474 8327 15476 8336
rect 15528 8327 15530 8336
rect 15476 8298 15528 8304
rect 15580 8294 15608 8774
rect 16302 8528 16358 8537
rect 16302 8463 16358 8472
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15568 8288 15620 8294
rect 15672 8265 15700 8298
rect 16212 8288 16264 8294
rect 15568 8230 15620 8236
rect 15658 8256 15714 8265
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15028 6458 15056 6802
rect 15212 6798 15240 8230
rect 16212 8230 16264 8236
rect 15658 8191 15714 8200
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15658 8120 15714 8129
rect 15807 8123 16115 8132
rect 15658 8055 15714 8064
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7546 15424 7686
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15304 6390 15332 7210
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15396 5534 15424 7142
rect 15488 6798 15516 7210
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15580 6322 15608 6598
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15672 6254 15700 8055
rect 16224 8022 16252 8230
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 16224 6254 16252 7482
rect 16316 6730 16344 8463
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16408 7546 16436 7822
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16408 7002 16436 7482
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6458 16436 6598
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 15396 5506 15516 5534
rect 15488 400 15516 5506
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 16500 474 16528 9862
rect 16592 9382 16620 10542
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8906 16620 9318
rect 16684 9178 16712 9862
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16592 7954 16620 8842
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16592 7410 16620 7890
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16684 7342 16712 7754
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16592 6934 16620 7142
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16776 6254 16804 11018
rect 16868 9024 16896 11154
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16960 9178 16988 10066
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16948 9036 17000 9042
rect 16868 8996 16948 9024
rect 16948 8978 17000 8984
rect 16960 8498 16988 8978
rect 17052 8974 17080 10202
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17144 9178 17172 10066
rect 17236 9994 17264 11206
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17512 10810 17540 11478
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 17236 9654 17264 9930
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17328 9042 17356 9862
rect 17696 9382 17724 10066
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8514 17080 8910
rect 17788 8673 17816 11580
rect 17868 11562 17920 11568
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17880 10266 17908 10542
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17774 8664 17830 8673
rect 17774 8599 17830 8608
rect 16948 8492 17000 8498
rect 17052 8486 17264 8514
rect 16948 8434 17000 8440
rect 17236 8430 17264 8486
rect 17972 8430 18000 9046
rect 17132 8424 17184 8430
rect 17130 8392 17132 8401
rect 17224 8424 17276 8430
rect 17184 8392 17186 8401
rect 17960 8424 18012 8430
rect 17224 8366 17276 8372
rect 17498 8392 17554 8401
rect 17130 8327 17186 8336
rect 17960 8366 18012 8372
rect 17498 8327 17554 8336
rect 17868 8356 17920 8362
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 17052 8022 17080 8230
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16868 5534 16896 6666
rect 16960 6458 16988 7210
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 7002 17080 7142
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 17144 6458 17172 7890
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 16776 5506 16896 5534
rect 16028 468 16080 474
rect 16488 468 16540 474
rect 16080 428 16160 456
rect 16028 410 16080 416
rect 16132 400 16160 428
rect 16488 410 16540 416
rect 16776 400 16804 5506
rect 17420 400 17448 7686
rect 17512 6866 17540 8327
rect 17774 8308 17830 8317
rect 17868 8298 17920 8304
rect 17774 8243 17830 8252
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17696 7546 17724 7890
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17682 6896 17738 6905
rect 17500 6860 17552 6866
rect 17682 6831 17684 6840
rect 17500 6802 17552 6808
rect 17736 6831 17738 6840
rect 17684 6802 17736 6808
rect 17512 6322 17540 6802
rect 17788 6458 17816 8243
rect 17880 6866 17908 8298
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17972 6798 18000 7686
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 18064 6322 18092 11494
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18248 10810 18276 11290
rect 18432 11218 18460 11630
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18340 8634 18368 11018
rect 18524 10742 18552 11494
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18420 9920 18472 9926
rect 18524 9908 18552 10678
rect 18616 10606 18644 10950
rect 18708 10810 18736 19600
rect 19352 12442 19380 19600
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19156 11824 19208 11830
rect 19260 11812 19288 12242
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19208 11784 19288 11812
rect 19156 11766 19208 11772
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18892 10606 18920 11494
rect 19076 11286 19104 11630
rect 19260 11286 19288 11784
rect 19444 11694 19472 12038
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10674 19380 10950
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 10130 19012 10406
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 18472 9880 18552 9908
rect 19064 9920 19116 9926
rect 18420 9862 18472 9868
rect 19064 9862 19116 9868
rect 18432 9432 18460 9862
rect 19076 9518 19104 9862
rect 19536 9654 19564 19638
rect 19904 19530 19932 19638
rect 19982 19600 20038 20000
rect 20626 19600 20682 20000
rect 19996 19530 20024 19600
rect 19904 19502 20024 19530
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 20640 11898 20668 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 31217 19068 31525 19077
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 31217 13628 31525 13637
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21284 12434 21312 12718
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 21284 12406 21404 12434
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 19984 10600 20036 10606
rect 20036 10548 20300 10554
rect 19984 10542 20300 10548
rect 19996 10526 20300 10542
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10130 19932 10406
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 20272 9994 20300 10526
rect 20260 9988 20312 9994
rect 20260 9930 20312 9936
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 18512 9444 18564 9450
rect 18432 9404 18512 9432
rect 19708 9444 19760 9450
rect 18512 9386 18564 9392
rect 19536 9404 19708 9432
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18326 8392 18382 8401
rect 18326 8327 18328 8336
rect 18380 8327 18382 8336
rect 18328 8298 18380 8304
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7954 18184 8230
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18156 7002 18184 7890
rect 18432 7546 18460 7958
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18156 6322 18184 6938
rect 18524 6866 18552 9386
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18616 7410 18644 8298
rect 18708 8294 18736 8774
rect 18800 8566 18828 8978
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 7886 18736 8230
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18972 7336 19024 7342
rect 19260 7313 19288 7482
rect 19352 7342 19380 9114
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19444 7478 19472 7890
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19340 7336 19392 7342
rect 18972 7278 19024 7284
rect 19246 7304 19302 7313
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18694 7032 18750 7041
rect 18694 6967 18696 6976
rect 18748 6967 18750 6976
rect 18696 6938 18748 6944
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18340 6186 18368 6734
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18800 6458 18828 6666
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18892 5534 18920 7142
rect 18984 7002 19012 7278
rect 19340 7278 19392 7284
rect 19246 7239 19302 7248
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 19260 6866 19288 7239
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19352 7002 19380 7142
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19444 6458 19472 7142
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19536 5534 19564 9404
rect 19708 9386 19760 9392
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19628 7002 19656 7346
rect 19892 7200 19944 7206
rect 19890 7168 19892 7177
rect 19944 7168 19946 7177
rect 19890 7103 19946 7112
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19706 6896 19762 6905
rect 19996 6866 20024 8298
rect 20088 7546 20116 9386
rect 20166 8392 20222 8401
rect 20166 8327 20222 8336
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20074 7440 20130 7449
rect 20074 7375 20076 7384
rect 20128 7375 20130 7384
rect 20076 7346 20128 7352
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 20088 6934 20116 7210
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 19706 6831 19708 6840
rect 19760 6831 19762 6840
rect 19984 6860 20036 6866
rect 19708 6802 19760 6808
rect 19984 6802 20036 6808
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 20180 5534 20208 8327
rect 20272 7546 20300 9930
rect 20732 9518 20760 10746
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21192 9466 21220 10406
rect 21284 10198 21312 10406
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20824 8090 20852 8774
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20272 7313 20300 7482
rect 20352 7336 20404 7342
rect 20258 7304 20314 7313
rect 20352 7278 20404 7284
rect 20258 7239 20314 7248
rect 20364 7041 20392 7278
rect 20350 7032 20406 7041
rect 20350 6967 20406 6976
rect 18708 5506 18920 5534
rect 19352 5506 19564 5534
rect 19996 5506 20208 5534
rect 20548 5534 20576 7686
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20640 7002 20668 7278
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20916 6186 20944 9318
rect 21100 9178 21128 9454
rect 21192 9438 21312 9466
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21192 9178 21220 9318
rect 21284 9178 21312 9438
rect 21376 9382 21404 12406
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21468 9518 21496 11630
rect 21732 10736 21784 10742
rect 21732 10678 21784 10684
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 10266 21588 10406
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21560 9518 21588 9930
rect 21652 9518 21680 10542
rect 21744 9518 21772 10678
rect 22020 10010 22048 12582
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28276 10985 28304 11018
rect 28262 10976 28318 10985
rect 27365 10908 27673 10917
rect 28262 10911 28318 10920
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 22192 10056 22244 10062
rect 22020 9982 22140 10010
rect 22192 9998 22244 10004
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22020 9518 22048 9862
rect 22112 9722 22140 9982
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22204 9586 22232 9998
rect 22296 9722 22324 10474
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31666 10296 31722 10305
rect 31666 10231 31668 10240
rect 31720 10231 31722 10240
rect 31668 10202 31720 10208
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22388 9602 22416 9658
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22296 9574 22416 9602
rect 22572 9586 22600 9930
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 28264 9648 28316 9654
rect 28262 9616 28264 9625
rect 28316 9616 28318 9625
rect 22560 9580 22612 9586
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 21364 9376 21416 9382
rect 22112 9330 22140 9386
rect 21364 9318 21416 9324
rect 21928 9302 22140 9330
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21008 7954 21036 8774
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 21008 7002 21036 7890
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20548 5506 20668 5534
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18064 400 18092 4082
rect 18708 400 18736 5506
rect 19352 400 19380 5506
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 19996 400 20024 5506
rect 20640 400 20668 5506
rect 21284 400 21312 7754
rect 21376 7478 21404 8366
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 21468 6662 21496 8366
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21560 6254 21588 8298
rect 21744 7886 21772 8366
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21836 8022 21864 8230
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21928 7449 21956 9302
rect 22296 9110 22324 9574
rect 28262 9551 28318 9560
rect 22560 9522 22612 9528
rect 22376 9512 22428 9518
rect 22376 9454 22428 9460
rect 22388 9110 22416 9454
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22572 9178 22600 9318
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 31217 9211 31525 9220
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22376 9104 22428 9110
rect 22376 9046 22428 9052
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 22020 8838 22048 8978
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22020 7546 22048 8366
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21914 7440 21970 7449
rect 21914 7375 21970 7384
rect 22204 7177 22232 8774
rect 22388 8566 22416 9046
rect 28262 8936 28318 8945
rect 28262 8871 28264 8880
rect 28316 8871 28318 8880
rect 28264 8842 28316 8848
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22190 7168 22246 7177
rect 22190 7103 22246 7112
rect 22480 6730 22508 8774
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31680 8265 31708 8434
rect 31666 8256 31722 8265
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 31217 8188 31525 8197
rect 31666 8191 31722 8200
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 31217 8123 31525 8132
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 27365 7579 27673 7588
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 27365 5468 27673 5477
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 31217 2748 31525 2757
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 14094 368 14150 377
rect 14094 303 14150 312
rect 14186 0 14242 400
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16118 0 16174 400
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 18050 0 18106 400
rect 18694 0 18750 400
rect 19338 0 19394 400
rect 19982 0 20038 400
rect 20626 0 20682 400
rect 21270 0 21326 400
<< via2 >>
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 8390 9968 8446 10024
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 7930 9036 7986 9072
rect 7930 9016 7932 9036
rect 7932 9016 7984 9036
rect 7984 9016 7986 9036
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 8390 8472 8446 8528
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 9954 11600 10010 11656
rect 9310 10104 9366 10160
rect 9034 9016 9090 9072
rect 8942 8880 8998 8936
rect 9494 9968 9550 10024
rect 9494 9716 9550 9752
rect 9494 9696 9496 9716
rect 9496 9696 9548 9716
rect 9548 9696 9550 9716
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 10138 9460 10140 9480
rect 10140 9460 10192 9480
rect 10192 9460 10194 9480
rect 10138 9424 10194 9460
rect 9862 7928 9918 7984
rect 10598 9696 10654 9752
rect 11242 11328 11298 11384
rect 11150 11192 11206 11248
rect 11610 11600 11666 11656
rect 11702 11328 11758 11384
rect 11426 11212 11482 11248
rect 11426 11192 11428 11212
rect 11428 11192 11480 11212
rect 11480 11192 11482 11212
rect 11058 10804 11114 10840
rect 11058 10784 11060 10804
rect 11060 10784 11112 10804
rect 11112 10784 11114 10804
rect 11334 10260 11390 10296
rect 11334 10240 11336 10260
rect 11336 10240 11388 10260
rect 11388 10240 11390 10260
rect 11150 9560 11206 9616
rect 10874 9444 10930 9480
rect 10874 9424 10876 9444
rect 10876 9424 10928 9444
rect 10928 9424 10930 9444
rect 10690 7520 10746 7576
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 10322 3712 10378 3768
rect 9678 3440 9734 3496
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 14830 12008 14886 12064
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 17130 12008 17186 12064
rect 12530 10104 12586 10160
rect 14002 9968 14058 10024
rect 11426 6840 11482 6896
rect 11794 7792 11850 7848
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 12162 7384 12218 7440
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 12806 8472 12862 8528
rect 11886 6296 11942 6352
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 13082 8472 13138 8528
rect 13818 8336 13874 8392
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 14462 8064 14518 8120
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 15474 8356 15530 8392
rect 15474 8336 15476 8356
rect 15476 8336 15528 8356
rect 15528 8336 15530 8356
rect 16302 8472 16358 8528
rect 15658 8200 15714 8256
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 15658 8064 15714 8120
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 17774 8608 17830 8664
rect 17130 8372 17132 8392
rect 17132 8372 17184 8392
rect 17184 8372 17186 8392
rect 17130 8336 17186 8372
rect 17498 8336 17554 8392
rect 17774 8252 17830 8308
rect 17682 6860 17738 6896
rect 17682 6840 17684 6860
rect 17684 6840 17736 6860
rect 17736 6840 17738 6860
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 18326 8356 18382 8392
rect 18326 8336 18328 8356
rect 18328 8336 18380 8356
rect 18380 8336 18382 8356
rect 18694 6996 18750 7032
rect 18694 6976 18696 6996
rect 18696 6976 18748 6996
rect 18748 6976 18750 6996
rect 19246 7248 19302 7304
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 19890 7148 19892 7168
rect 19892 7148 19944 7168
rect 19944 7148 19946 7168
rect 19890 7112 19946 7148
rect 19706 6860 19762 6896
rect 20166 8336 20222 8392
rect 20074 7404 20130 7440
rect 20074 7384 20076 7404
rect 20076 7384 20128 7404
rect 20128 7384 20130 7404
rect 19706 6840 19708 6860
rect 19708 6840 19760 6860
rect 19760 6840 19762 6860
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 20258 7248 20314 7304
rect 20350 6976 20406 7032
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 28262 10920 28318 10976
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10260 31722 10296
rect 31666 10240 31668 10260
rect 31668 10240 31720 10260
rect 31720 10240 31722 10260
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 28262 9596 28264 9616
rect 28264 9596 28316 9616
rect 28316 9596 28318 9616
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 28262 9560 28318 9596
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 21914 7384 21970 7440
rect 28262 8900 28318 8936
rect 28262 8880 28264 8900
rect 28264 8880 28316 8900
rect 28316 8880 28318 8900
rect 22190 7112 22246 7168
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 31666 8200 31722 8256
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
rect 14094 312 14150 368
<< metal3 >>
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31213 19007 31529 19008
rect 4246 18528 4562 18529
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31213 13567 31529 13568
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 14825 12066 14891 12069
rect 17125 12066 17191 12069
rect 14825 12064 17191 12066
rect 14825 12008 14830 12064
rect 14886 12008 17130 12064
rect 17186 12008 17191 12064
rect 14825 12006 17191 12008
rect 14825 12003 14891 12006
rect 17125 12003 17191 12006
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 0 11658 400 11688
rect 9949 11658 10015 11661
rect 11605 11658 11671 11661
rect 0 11656 11671 11658
rect 0 11600 9954 11656
rect 10010 11600 11610 11656
rect 11666 11600 11671 11656
rect 0 11598 11671 11600
rect 0 11568 400 11598
rect 9949 11595 10015 11598
rect 11605 11595 11671 11598
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 11237 11386 11303 11389
rect 11697 11386 11763 11389
rect 11237 11384 11763 11386
rect 11237 11328 11242 11384
rect 11298 11328 11702 11384
rect 11758 11328 11763 11384
rect 11237 11326 11763 11328
rect 11237 11323 11303 11326
rect 11697 11323 11763 11326
rect 11145 11250 11211 11253
rect 11421 11250 11487 11253
rect 11145 11248 11487 11250
rect 11145 11192 11150 11248
rect 11206 11192 11426 11248
rect 11482 11192 11487 11248
rect 11145 11190 11487 11192
rect 11145 11187 11211 11190
rect 11421 11187 11487 11190
rect 0 10978 400 11008
rect 28257 10978 28323 10981
rect 31600 10978 32000 11008
rect 0 10918 2790 10978
rect 0 10888 400 10918
rect 2730 10706 2790 10918
rect 28257 10976 32000 10978
rect 28257 10920 28262 10976
rect 28318 10920 32000 10976
rect 28257 10918 32000 10920
rect 28257 10915 28323 10918
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 31600 10888 32000 10918
rect 27361 10847 27677 10848
rect 11053 10842 11119 10845
rect 6870 10840 11119 10842
rect 6870 10784 11058 10840
rect 11114 10784 11119 10840
rect 6870 10782 11119 10784
rect 6870 10706 6930 10782
rect 11053 10779 11119 10782
rect 2730 10646 6930 10706
rect 8098 10368 8414 10369
rect 0 10298 400 10328
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 11329 10298 11395 10301
rect 0 10238 2790 10298
rect 0 10208 400 10238
rect 2730 10162 2790 10238
rect 8526 10296 11395 10298
rect 8526 10240 11334 10296
rect 11390 10240 11395 10296
rect 8526 10238 11395 10240
rect 8526 10162 8586 10238
rect 11329 10235 11395 10238
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 2730 10102 8586 10162
rect 9305 10162 9371 10165
rect 12525 10162 12591 10165
rect 9305 10160 12591 10162
rect 9305 10104 9310 10160
rect 9366 10104 12530 10160
rect 12586 10104 12591 10160
rect 9305 10102 12591 10104
rect 9305 10099 9371 10102
rect 12525 10099 12591 10102
rect 8385 10026 8451 10029
rect 9489 10026 9555 10029
rect 8385 10024 9555 10026
rect 8385 9968 8390 10024
rect 8446 9968 9494 10024
rect 9550 9968 9555 10024
rect 8385 9966 9555 9968
rect 8385 9963 8451 9966
rect 9489 9963 9555 9966
rect 13997 10028 14063 10029
rect 13997 10024 14044 10028
rect 14108 10026 14114 10028
rect 13997 9968 14002 10024
rect 13997 9964 14044 9968
rect 14108 9966 14154 10026
rect 14108 9964 14114 9966
rect 13997 9963 14063 9964
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 9489 9754 9555 9757
rect 10593 9754 10659 9757
rect 9489 9752 10659 9754
rect 9489 9696 9494 9752
rect 9550 9696 10598 9752
rect 10654 9696 10659 9752
rect 9489 9694 10659 9696
rect 9489 9691 9555 9694
rect 10593 9691 10659 9694
rect 0 9618 400 9648
rect 11145 9618 11211 9621
rect 0 9616 11211 9618
rect 0 9560 11150 9616
rect 11206 9560 11211 9616
rect 0 9558 11211 9560
rect 0 9528 400 9558
rect 11145 9555 11211 9558
rect 28257 9618 28323 9621
rect 31600 9618 32000 9648
rect 28257 9616 32000 9618
rect 28257 9560 28262 9616
rect 28318 9560 32000 9616
rect 28257 9558 32000 9560
rect 28257 9555 28323 9558
rect 31600 9528 32000 9558
rect 10133 9482 10199 9485
rect 10869 9482 10935 9485
rect 10133 9480 10935 9482
rect 10133 9424 10138 9480
rect 10194 9424 10874 9480
rect 10930 9424 10935 9480
rect 10133 9422 10935 9424
rect 10133 9419 10199 9422
rect 10869 9419 10935 9422
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 7925 9074 7991 9077
rect 9029 9074 9095 9077
rect 7925 9072 9095 9074
rect 7925 9016 7930 9072
rect 7986 9016 9034 9072
rect 9090 9016 9095 9072
rect 7925 9014 9095 9016
rect 7925 9011 7991 9014
rect 9029 9011 9095 9014
rect 0 8938 400 8968
rect 8937 8938 9003 8941
rect 0 8936 9003 8938
rect 0 8880 8942 8936
rect 8998 8880 9003 8936
rect 0 8878 9003 8880
rect 0 8848 400 8878
rect 8937 8875 9003 8878
rect 28257 8938 28323 8941
rect 31600 8938 32000 8968
rect 28257 8936 32000 8938
rect 28257 8880 28262 8936
rect 28318 8880 32000 8936
rect 28257 8878 32000 8880
rect 28257 8875 28323 8878
rect 31600 8848 32000 8878
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 17769 8666 17835 8669
rect 17726 8664 17835 8666
rect 17726 8608 17774 8664
rect 17830 8608 17835 8664
rect 17726 8603 17835 8608
rect 8385 8530 8451 8533
rect 12801 8530 12867 8533
rect 8385 8528 12867 8530
rect 8385 8472 8390 8528
rect 8446 8472 12806 8528
rect 12862 8472 12867 8528
rect 8385 8470 12867 8472
rect 8385 8467 8451 8470
rect 12801 8467 12867 8470
rect 13077 8530 13143 8533
rect 16297 8530 16363 8533
rect 13077 8528 16363 8530
rect 13077 8472 13082 8528
rect 13138 8472 16302 8528
rect 16358 8472 16363 8528
rect 13077 8470 16363 8472
rect 13077 8467 13143 8470
rect 16297 8467 16363 8470
rect 13813 8396 13879 8397
rect 13813 8392 13860 8396
rect 13924 8394 13930 8396
rect 13813 8336 13818 8392
rect 13813 8332 13860 8336
rect 13924 8334 13970 8394
rect 13924 8332 13930 8334
rect 15142 8332 15148 8396
rect 15212 8394 15218 8396
rect 15469 8394 15535 8397
rect 15212 8392 15535 8394
rect 15212 8336 15474 8392
rect 15530 8336 15535 8392
rect 15212 8334 15535 8336
rect 15212 8332 15218 8334
rect 13813 8331 13879 8332
rect 15469 8331 15535 8334
rect 17125 8394 17191 8397
rect 17493 8394 17559 8397
rect 17125 8392 17559 8394
rect 17125 8336 17130 8392
rect 17186 8336 17498 8392
rect 17554 8336 17559 8392
rect 17125 8334 17559 8336
rect 17125 8331 17191 8334
rect 17493 8331 17559 8334
rect 17726 8313 17786 8603
rect 18321 8394 18387 8397
rect 20161 8394 20227 8397
rect 18321 8392 20227 8394
rect 18321 8336 18326 8392
rect 18382 8336 20166 8392
rect 20222 8336 20227 8392
rect 18321 8334 20227 8336
rect 18321 8331 18387 8334
rect 20161 8331 20227 8334
rect 17726 8308 17835 8313
rect 0 8258 400 8288
rect 15653 8258 15719 8261
rect 0 8198 2790 8258
rect 0 8168 400 8198
rect 2730 7986 2790 8198
rect 15518 8256 15719 8258
rect 15518 8200 15658 8256
rect 15714 8200 15719 8256
rect 17726 8252 17774 8308
rect 17830 8252 17835 8308
rect 17726 8250 17835 8252
rect 17769 8247 17835 8250
rect 31600 8256 32000 8288
rect 15518 8198 15719 8200
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 14457 8122 14523 8125
rect 15518 8122 15578 8198
rect 15653 8195 15719 8198
rect 31600 8200 31666 8256
rect 31722 8200 32000 8256
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31600 8168 32000 8200
rect 31213 8127 31529 8128
rect 15653 8122 15719 8125
rect 14457 8120 15719 8122
rect 14457 8064 14462 8120
rect 14518 8064 15658 8120
rect 15714 8064 15719 8120
rect 14457 8062 15719 8064
rect 14457 8059 14523 8062
rect 15653 8059 15719 8062
rect 9857 7986 9923 7989
rect 2730 7984 9923 7986
rect 2730 7928 9862 7984
rect 9918 7928 9923 7984
rect 2730 7926 9923 7928
rect 9857 7923 9923 7926
rect 11789 7850 11855 7853
rect 11654 7848 11855 7850
rect 11654 7792 11794 7848
rect 11850 7792 11855 7848
rect 11654 7790 11855 7792
rect 4246 7648 4562 7649
rect 0 7578 400 7608
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 10685 7578 10751 7581
rect 0 7518 2790 7578
rect 0 7488 400 7518
rect 2730 7442 2790 7518
rect 4662 7576 10751 7578
rect 4662 7520 10690 7576
rect 10746 7520 10751 7576
rect 4662 7518 10751 7520
rect 4662 7442 4722 7518
rect 10685 7515 10751 7518
rect 2730 7382 4722 7442
rect 11654 7442 11714 7790
rect 11789 7787 11855 7790
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 12157 7442 12223 7445
rect 11654 7440 12223 7442
rect 11654 7384 12162 7440
rect 12218 7384 12223 7440
rect 11654 7382 12223 7384
rect 12157 7379 12223 7382
rect 20069 7442 20135 7445
rect 21909 7442 21975 7445
rect 20069 7440 21975 7442
rect 20069 7384 20074 7440
rect 20130 7384 21914 7440
rect 21970 7384 21975 7440
rect 20069 7382 21975 7384
rect 20069 7379 20135 7382
rect 21909 7379 21975 7382
rect 19241 7306 19307 7309
rect 20253 7306 20319 7309
rect 19241 7304 20319 7306
rect 19241 7248 19246 7304
rect 19302 7248 20258 7304
rect 20314 7248 20319 7304
rect 19241 7246 20319 7248
rect 19241 7243 19307 7246
rect 20253 7243 20319 7246
rect 19885 7170 19951 7173
rect 22185 7170 22251 7173
rect 19885 7168 22251 7170
rect 19885 7112 19890 7168
rect 19946 7112 22190 7168
rect 22246 7112 22251 7168
rect 19885 7110 22251 7112
rect 19885 7107 19951 7110
rect 22185 7107 22251 7110
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 18689 7034 18755 7037
rect 20345 7034 20411 7037
rect 18689 7032 20411 7034
rect 18689 6976 18694 7032
rect 18750 6976 20350 7032
rect 20406 6976 20411 7032
rect 18689 6974 20411 6976
rect 18689 6971 18755 6974
rect 20345 6971 20411 6974
rect 11421 6898 11487 6901
rect 17677 6898 17743 6901
rect 19701 6898 19767 6901
rect 11421 6896 11714 6898
rect 11421 6840 11426 6896
rect 11482 6840 11714 6896
rect 11421 6838 11714 6840
rect 11421 6835 11487 6838
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11654 6354 11714 6838
rect 17677 6896 19767 6898
rect 17677 6840 17682 6896
rect 17738 6840 19706 6896
rect 19762 6840 19767 6896
rect 17677 6838 19767 6840
rect 17677 6835 17743 6838
rect 19701 6835 19767 6838
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 11881 6354 11947 6357
rect 11654 6352 11947 6354
rect 11654 6296 11886 6352
rect 11942 6296 11947 6352
rect 11654 6294 11947 6296
rect 11881 6291 11947 6294
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 27361 5407 27677 5408
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 10317 3770 10383 3773
rect 14038 3770 14044 3772
rect 10317 3768 14044 3770
rect 10317 3712 10322 3768
rect 10378 3712 14044 3768
rect 10317 3710 14044 3712
rect 10317 3707 10383 3710
rect 14038 3708 14044 3710
rect 14108 3708 14114 3772
rect 9673 3498 9739 3501
rect 13854 3498 13860 3500
rect 9673 3496 13860 3498
rect 9673 3440 9678 3496
rect 9734 3440 13860 3496
rect 9673 3438 13860 3440
rect 9673 3435 9739 3438
rect 13854 3436 13860 3438
rect 13924 3436 13930 3500
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
rect 14089 370 14155 373
rect 15326 370 15332 372
rect 14089 368 15332 370
rect 14089 312 14094 368
rect 14150 312 15332 368
rect 14089 310 15332 312
rect 14089 307 14155 310
rect 15326 308 15332 310
rect 15396 308 15402 372
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 14044 10024 14108 10028
rect 14044 9968 14058 10024
rect 14058 9968 14108 10024
rect 14044 9964 14108 9968
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 13860 8392 13924 8396
rect 13860 8336 13874 8392
rect 13874 8336 13924 8392
rect 13860 8332 13924 8336
rect 15148 8332 15212 8396
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 14044 3708 14108 3772
rect 13860 3436 13924 3500
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
rect 15332 308 15396 372
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11949 12000 12269 13024
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 15801 15808 16121 16832
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 15801 10368 16121 11392
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 14043 10028 14109 10029
rect 14043 9964 14044 10028
rect 14108 9964 14109 10028
rect 14043 9963 14109 9964
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 11949 8736 12269 9760
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 13859 8396 13925 8397
rect 13859 8332 13860 8396
rect 13924 8332 13925 8396
rect 13859 8331 13925 8332
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 11949 6560 12269 7584
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 13862 3501 13922 8331
rect 14046 3773 14106 9963
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15147 8396 15213 8397
rect 15147 8332 15148 8396
rect 15212 8332 15213 8396
rect 15147 8331 15213 8332
rect 15150 5550 15210 8331
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15150 5490 15394 5550
rect 14043 3772 14109 3773
rect 14043 3708 14044 3772
rect 14108 3708 14109 3772
rect 14043 3707 14109 3708
rect 13859 3500 13925 3501
rect 13859 3436 13860 3500
rect 13924 3436 13925 3500
rect 13859 3435 13925 3436
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15334 373 15394 5490
rect 15801 4928 16121 5952
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15801 3840 16121 4864
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19654 12000 19974 13024
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19654 7648 19974 8672
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 19654 4384 19974 5408
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 23506 15808 23826 16832
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
rect 15331 372 15397 373
rect 15331 308 15332 372
rect 15396 308 15397 372
rect 15331 307 15397 308
use sky130_fd_sc_hd__inv_2  _10__5 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16652 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__6
timestamp 1701704242
transform -1 0 15732 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__7
timestamp 1701704242
transform 1 0 13892 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__8
timestamp 1701704242
transform -1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__9
timestamp 1701704242
transform -1 0 8832 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__10
timestamp 1701704242
transform -1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__11
timestamp 1701704242
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__12
timestamp 1701704242
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__13
timestamp 1701704242
transform -1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__14
timestamp 1701704242
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__15
timestamp 1701704242
transform 1 0 17756 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__16
timestamp 1701704242
transform 1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__17
timestamp 1701704242
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__18
timestamp 1701704242
transform -1 0 19780 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__19
timestamp 1701704242
transform 1 0 14536 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__20
timestamp 1701704242
transform -1 0 16192 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10_
timestamp 1701704242
transform -1 0 14260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12880 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _12_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 12420 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _13_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12144 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _14_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12420 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _15_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14168 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _16_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13248 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _17_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16008 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _18_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14628 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _19_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17296 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _20_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17756 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _21_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16928 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1701704242
transform -1 0 17572 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _23_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _24_
timestamp 1701704242
transform 1 0 14904 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _25_
timestamp 1701704242
transform 1 0 17296 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _26_
timestamp 1701704242
transform 1 0 13984 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _27_
timestamp 1701704242
transform 1 0 11868 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _28_
timestamp 1701704242
transform 1 0 9384 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _29_
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _30_
timestamp 1701704242
transform 1 0 9200 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _31_
timestamp 1701704242
transform 1 0 9200 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _32_
timestamp 1701704242
transform 1 0 10672 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _33_
timestamp 1701704242
transform 1 0 12604 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _34_
timestamp 1701704242
transform 1 0 15180 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _35_
timestamp 1701704242
transform 1 0 16928 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _36_
timestamp 1701704242
transform 1 0 18676 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _37_
timestamp 1701704242
transform 1 0 19136 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _38_
timestamp 1701704242
transform 1 0 19228 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _39_
timestamp 1701704242
transform 1 0 19228 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _40_
timestamp 1701704242
transform 1 0 17664 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _41_
timestamp 1701704242
transform 1 0 15824 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _42_
timestamp 1701704242
transform 1 0 17204 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _43_
timestamp 1701704242
transform 1 0 18952 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _44_
timestamp 1701704242
transform 1 0 19136 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _45_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12604 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1701704242
transform -1 0 16468 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _47_
timestamp 1701704242
transform -1 0 16652 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _48_
timestamp 1701704242
transform 1 0 13892 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _49_
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _50_
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _51_
timestamp 1701704242
transform -1 0 9844 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _52_
timestamp 1701704242
transform -1 0 10396 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _53_
timestamp 1701704242
transform 1 0 11040 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _54_
timestamp 1701704242
transform -1 0 13156 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _55_
timestamp 1701704242
transform -1 0 15180 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _56_
timestamp 1701704242
transform -1 0 17296 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _57_
timestamp 1701704242
transform -1 0 18676 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _58_
timestamp 1701704242
transform -1 0 18584 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _59_
timestamp 1701704242
transform -1 0 20240 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _60_
timestamp 1701704242
transform -1 0 20792 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _61_
timestamp 1701704242
transform 1 0 15180 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _62_
timestamp 1701704242
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _63_
timestamp 1701704242
transform 1 0 13432 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _64_
timestamp 1701704242
transform -1 0 19504 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _65_
timestamp 1701704242
transform 1 0 19504 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _66_
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _67_
timestamp 1701704242
transform 1 0 20424 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _68_
timestamp 1701704242
transform 1 0 20608 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _69_
timestamp 1701704242
transform 1 0 15456 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _70_
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _71_
timestamp 1701704242
transform 1 0 10948 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _72_
timestamp 1701704242
transform 1 0 14996 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _73_
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _74_
timestamp 1701704242
transform 1 0 10488 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _75_
timestamp 1701704242
transform 1 0 12144 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _76_
timestamp 1701704242
transform 1 0 13984 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _77_
timestamp 1701704242
transform 1 0 16560 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _78_
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _79_
timestamp 1701704242
transform 1 0 20148 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _80_
timestamp 1701704242
transform 1 0 20608 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _81_
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _82_
timestamp 1701704242
transform 1 0 21252 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _83_
timestamp 1701704242
transform 1 0 19136 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _84_
timestamp 1701704242
transform 1 0 17296 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1701704242
transform -1 0 15916 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1701704242
transform 1 0 12880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_stop pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14168 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net5
timestamp 1701704242
transform 1 0 14812 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_i_stop
timestamp 1701704242
transform -1 0 13432 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net5
timestamp 1701704242
transform -1 0 14076 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_i_stop
timestamp 1701704242
transform 1 0 16744 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net5
timestamp 1701704242
transform 1 0 17388 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__nor2_1  dly_stg1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9936 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg2
timestamp 1701704242
transform 1 0 13064 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  dly_stg5 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13432 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg6_219
timestamp 1701704242
transform 1 0 14444 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_86
timestamp 1701704242
transform 1 0 13616 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_87
timestamp 1701704242
transform -1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_88
timestamp 1701704242
transform -1 0 12236 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_129
timestamp 1701704242
transform -1 0 12236 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_130
timestamp 1701704242
transform 1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_131
timestamp 1701704242
transform -1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_132
timestamp 1701704242
transform 1 0 16376 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_133
timestamp 1701704242
transform -1 0 15088 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_134
timestamp 1701704242
transform 1 0 17756 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_135
timestamp 1701704242
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_136
timestamp 1701704242
transform 1 0 13800 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_137
timestamp 1701704242
transform 1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_182
timestamp 1701704242
transform -1 0 12972 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_183
timestamp 1701704242
transform 1 0 12236 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_184
timestamp 1701704242
transform -1 0 10948 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_89
timestamp 1701704242
transform -1 0 12328 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_90
timestamp 1701704242
transform -1 0 11592 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_91
timestamp 1701704242
transform 1 0 12512 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_92
timestamp 1701704242
transform 1 0 12788 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_93
timestamp 1701704242
transform -1 0 10672 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1701704242
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1701704242
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1701704242
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1701704242
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1701704242
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1701704242
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1701704242
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1701704242
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1701704242
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_329
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1701704242
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1701704242
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1701704242
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1701704242
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1701704242
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1701704242
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1701704242
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1701704242
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1701704242
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1701704242
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1701704242
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1701704242
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1701704242
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1701704242
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1701704242
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1701704242
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1701704242
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1701704242
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1701704242
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1701704242
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1701704242
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1701704242
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1701704242
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1701704242
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1701704242
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1701704242
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1701704242
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1701704242
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1701704242
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1701704242
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1701704242
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1701704242
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1701704242
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1701704242
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1701704242
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1701704242
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1701704242
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1701704242
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1701704242
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1701704242
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1701704242
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_329
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1701704242
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1701704242
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1701704242
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1701704242
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1701704242
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1701704242
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1701704242
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1701704242
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1701704242
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1701704242
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1701704242
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1701704242
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1701704242
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1701704242
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1701704242
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1701704242
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1701704242
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1701704242
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1701704242
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1701704242
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1701704242
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1701704242
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1701704242
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1701704242
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1701704242
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1701704242
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1701704242
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1701704242
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1701704242
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1701704242
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1701704242
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1701704242
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1701704242
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1701704242
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1701704242
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1701704242
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1701704242
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1701704242
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1701704242
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1701704242
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1701704242
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1701704242
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1701704242
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_329
timestamp 1701704242
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1701704242
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1701704242
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1701704242
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1701704242
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1701704242
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1701704242
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1701704242
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1701704242
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1701704242
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1701704242
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1701704242
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1701704242
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1701704242
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1701704242
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1701704242
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1701704242
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1701704242
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1701704242
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1701704242
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1701704242
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1701704242
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_329
timestamp 1701704242
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1701704242
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1701704242
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1701704242
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1701704242
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_121
timestamp 1701704242
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_133
timestamp 1701704242
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1701704242
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1701704242
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1701704242
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1701704242
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1701704242
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1701704242
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1701704242
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1701704242
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1701704242
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1701704242
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1701704242
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1701704242
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1701704242
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1701704242
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1701704242
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1701704242
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1701704242
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1701704242
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 1701704242
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_329
timestamp 1701704242
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1701704242
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1701704242
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1701704242
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1701704242
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1701704242
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1701704242
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_121 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_132
timestamp 1701704242
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_143
timestamp 1701704242
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_148
timestamp 1701704242
transform 1 0 14168 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_160
timestamp 1701704242
transform 1 0 15272 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1701704242
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1701704242
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1701704242
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1701704242
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1701704242
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1701704242
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1701704242
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1701704242
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1701704242
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1701704242
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1701704242
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1701704242
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1701704242
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1701704242
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1701704242
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_329
timestamp 1701704242
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1701704242
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1701704242
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1701704242
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1701704242
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1701704242
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1701704242
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_109
timestamp 1701704242
transform 1 0 10580 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_151
timestamp 1701704242
transform 1 0 14444 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_155
timestamp 1701704242
transform 1 0 14812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_168
timestamp 1701704242
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_174
timestamp 1701704242
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_185
timestamp 1701704242
transform 1 0 17572 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1701704242
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1701704242
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1701704242
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1701704242
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1701704242
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1701704242
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1701704242
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1701704242
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1701704242
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1701704242
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1701704242
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1701704242
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_321
timestamp 1701704242
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 1701704242
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1701704242
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1701704242
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1701704242
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_93
timestamp 1701704242
transform 1 0 9108 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_99
timestamp 1701704242
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_119
timestamp 1701704242
transform 1 0 11500 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_129
timestamp 1701704242
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_147
timestamp 1701704242
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1701704242
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_186
timestamp 1701704242
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_191
timestamp 1701704242
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1701704242
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1701704242
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1701704242
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1701704242
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1701704242
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1701704242
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1701704242
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1701704242
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1701704242
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1701704242
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_329
timestamp 1701704242
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1701704242
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1701704242
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1701704242
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1701704242
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1701704242
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1701704242
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1701704242
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_85
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_94
timestamp 1701704242
transform 1 0 9200 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_126
timestamp 1701704242
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_152
timestamp 1701704242
transform 1 0 14536 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1701704242
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1701704242
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1701704242
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1701704242
transform 1 0 23092 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1701704242
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1701704242
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1701704242
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1701704242
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1701704242
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1701704242
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1701704242
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_321
timestamp 1701704242
transform 1 0 30084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_329
timestamp 1701704242
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1701704242
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1701704242
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1701704242
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1701704242
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1701704242
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 1701704242
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_93
timestamp 1701704242
transform 1 0 9108 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1701704242
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_132
timestamp 1701704242
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_149
timestamp 1701704242
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_169
timestamp 1701704242
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_174
timestamp 1701704242
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1701704242
transform 1 0 20976 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1701704242
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1701704242
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1701704242
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1701704242
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1701704242
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1701704242
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1701704242
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1701704242
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1701704242
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_329
timestamp 1701704242
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1701704242
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_77
timestamp 1701704242
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_94
timestamp 1701704242
transform 1 0 9200 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_107
timestamp 1701704242
transform 1 0 10396 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_114
timestamp 1701704242
transform 1 0 11040 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_124
timestamp 1701704242
transform 1 0 11960 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_170
timestamp 1701704242
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_200
timestamp 1701704242
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_236
timestamp 1701704242
transform 1 0 22264 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_248
timestamp 1701704242
transform 1 0 23368 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1701704242
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1701704242
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1701704242
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1701704242
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1701704242
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1701704242
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_321
timestamp 1701704242
transform 1 0 30084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_329
timestamp 1701704242
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1701704242
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1701704242
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_69
timestamp 1701704242
transform 1 0 6900 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_93
timestamp 1701704242
transform 1 0 9108 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1701704242
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_119
timestamp 1701704242
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_147
timestamp 1701704242
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_173
timestamp 1701704242
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1701704242
transform 1 0 20976 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_240
timestamp 1701704242
transform 1 0 22632 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_252
timestamp 1701704242
transform 1 0 23736 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_264
timestamp 1701704242
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_276
timestamp 1701704242
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1701704242
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1701704242
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1701704242
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1701704242
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_329
timestamp 1701704242
transform 1 0 30820 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1701704242
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1701704242
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1701704242
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_77
timestamp 1701704242
transform 1 0 7636 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_153
timestamp 1701704242
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_175
timestamp 1701704242
transform 1 0 16652 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_200
timestamp 1701704242
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1701704242
transform 1 0 23552 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1701704242
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1701704242
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1701704242
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1701704242
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1701704242
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1701704242
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1701704242
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1701704242
transform 1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_329
timestamp 1701704242
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1701704242
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1701704242
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1701704242
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_81
timestamp 1701704242
transform 1 0 8004 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_119
timestamp 1701704242
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_151
timestamp 1701704242
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_184
timestamp 1701704242
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_202
timestamp 1701704242
transform 1 0 19136 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1701704242
transform 1 0 20976 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1701704242
transform 1 0 22356 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1701704242
transform 1 0 23460 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1701704242
transform 1 0 24564 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1701704242
transform 1 0 25668 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1701704242
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1701704242
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1701704242
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1701704242
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_329
timestamp 1701704242
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1701704242
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1701704242
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1701704242
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1701704242
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1701704242
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1701704242
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_119
timestamp 1701704242
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1701704242
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_147
timestamp 1701704242
transform 1 0 14076 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1701704242
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_230
timestamp 1701704242
transform 1 0 21712 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_242
timestamp 1701704242
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1701704242
transform 1 0 23552 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1701704242
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1701704242
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1701704242
transform 1 0 27140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1701704242
transform 1 0 28244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1701704242
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_321
timestamp 1701704242
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_329
timestamp 1701704242
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1701704242
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1701704242
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1701704242
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1701704242
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1701704242
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1701704242
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_93
timestamp 1701704242
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_138
timestamp 1701704242
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 1701704242
transform 1 0 20976 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1701704242
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1701704242
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1701704242
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1701704242
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1701704242
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1701704242
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1701704242
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1701704242
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1701704242
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1701704242
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_329
timestamp 1701704242
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1701704242
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1701704242
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1701704242
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1701704242
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1701704242
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1701704242
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_97
timestamp 1701704242
transform 1 0 9476 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_105
timestamp 1701704242
transform 1 0 10212 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_135
timestamp 1701704242
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_148
timestamp 1701704242
transform 1 0 14168 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_153
timestamp 1701704242
transform 1 0 14628 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_175
timestamp 1701704242
transform 1 0 16652 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_200
timestamp 1701704242
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_224
timestamp 1701704242
transform 1 0 21160 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_236
timestamp 1701704242
transform 1 0 22264 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_248
timestamp 1701704242
transform 1 0 23368 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1701704242
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1701704242
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1701704242
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1701704242
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1701704242
transform 1 0 28244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1701704242
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1701704242
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_329
timestamp 1701704242
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1701704242
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1701704242
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1701704242
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1701704242
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1701704242
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1701704242
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_154
timestamp 1701704242
transform 1 0 14720 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_158
timestamp 1701704242
transform 1 0 15088 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_169
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_175
timestamp 1701704242
transform 1 0 16652 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_198
timestamp 1701704242
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_212
timestamp 1701704242
transform 1 0 20056 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1701704242
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1701704242
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1701704242
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1701704242
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1701704242
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1701704242
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1701704242
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1701704242
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1701704242
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_329
timestamp 1701704242
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1701704242
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1701704242
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1701704242
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1701704242
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1701704242
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1701704242
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1701704242
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1701704242
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1701704242
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_141
timestamp 1701704242
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_147
timestamp 1701704242
transform 1 0 14076 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_159
timestamp 1701704242
transform 1 0 15180 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1701704242
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_177
timestamp 1701704242
transform 1 0 16836 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_181
timestamp 1701704242
transform 1 0 17204 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_185
timestamp 1701704242
transform 1 0 17572 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1701704242
transform 1 0 18308 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_200
timestamp 1701704242
transform 1 0 18952 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_212
timestamp 1701704242
transform 1 0 20056 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_224
timestamp 1701704242
transform 1 0 21160 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_236
timestamp 1701704242
transform 1 0 22264 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_248
timestamp 1701704242
transform 1 0 23368 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1701704242
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1701704242
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1701704242
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1701704242
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1701704242
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 1701704242
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1701704242
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1701704242
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1701704242
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1701704242
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1701704242
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1701704242
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1701704242
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1701704242
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1701704242
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1701704242
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1701704242
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1701704242
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1701704242
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1701704242
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1701704242
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1701704242
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1701704242
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1701704242
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1701704242
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1701704242
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1701704242
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1701704242
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1701704242
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1701704242
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1701704242
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1701704242
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1701704242
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1701704242
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1701704242
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_329
timestamp 1701704242
transform 1 0 30820 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1701704242
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1701704242
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1701704242
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1701704242
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1701704242
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1701704242
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1701704242
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1701704242
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1701704242
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1701704242
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1701704242
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1701704242
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1701704242
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1701704242
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1701704242
transform 1 0 17940 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1701704242
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1701704242
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1701704242
transform 1 0 20884 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1701704242
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1701704242
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1701704242
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1701704242
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1701704242
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1701704242
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1701704242
transform 1 0 27140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1701704242
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1701704242
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 1701704242
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_329
timestamp 1701704242
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1701704242
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1701704242
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1701704242
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1701704242
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1701704242
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1701704242
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1701704242
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1701704242
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1701704242
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1701704242
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1701704242
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1701704242
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1701704242
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1701704242
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1701704242
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1701704242
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1701704242
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1701704242
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1701704242
transform 1 0 20516 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1701704242
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1701704242
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1701704242
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1701704242
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1701704242
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1701704242
transform 1 0 25668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1701704242
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1701704242
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1701704242
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1701704242
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_329
timestamp 1701704242
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1701704242
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1701704242
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1701704242
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1701704242
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1701704242
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1701704242
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1701704242
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1701704242
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1701704242
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1701704242
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1701704242
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1701704242
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1701704242
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1701704242
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1701704242
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1701704242
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1701704242
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1701704242
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1701704242
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1701704242
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1701704242
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1701704242
transform 1 0 23092 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1701704242
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1701704242
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1701704242
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1701704242
transform 1 0 27140 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1701704242
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1701704242
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1701704242
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1701704242
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1701704242
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1701704242
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1701704242
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1701704242
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1701704242
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1701704242
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1701704242
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1701704242
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1701704242
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1701704242
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1701704242
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1701704242
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1701704242
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1701704242
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1701704242
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1701704242
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1701704242
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1701704242
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1701704242
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1701704242
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1701704242
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1701704242
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1701704242
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_329
timestamp 1701704242
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1701704242
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1701704242
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1701704242
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1701704242
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1701704242
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1701704242
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1701704242
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1701704242
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1701704242
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1701704242
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1701704242
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1701704242
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1701704242
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1701704242
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1701704242
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1701704242
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1701704242
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1701704242
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1701704242
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1701704242
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1701704242
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1701704242
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1701704242
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1701704242
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1701704242
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1701704242
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1701704242
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1701704242
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1701704242
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1701704242
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1701704242
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1701704242
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1701704242
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1701704242
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1701704242
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1701704242
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1701704242
transform 1 0 20516 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1701704242
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1701704242
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1701704242
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1701704242
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1701704242
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1701704242
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1701704242
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1701704242
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1701704242
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1701704242
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1701704242
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1701704242
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1701704242
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1701704242
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1701704242
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1701704242
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1701704242
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1701704242
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1701704242
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1701704242
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1701704242
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1701704242
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1701704242
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1701704242
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1701704242
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1701704242
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1701704242
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1701704242
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1701704242
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1701704242
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1701704242
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1701704242
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1701704242
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1701704242
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1701704242
transform 1 0 20516 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1701704242
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1701704242
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1701704242
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1701704242
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1701704242
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1701704242
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1701704242
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1701704242
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1701704242
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1701704242
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1701704242
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1701704242
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1701704242
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1701704242
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1701704242
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1701704242
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1701704242
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1701704242
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1701704242
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_131
timestamp 1701704242
transform 1 0 12604 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_139
timestamp 1701704242
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_153
timestamp 1701704242
transform 1 0 14628 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1701704242
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 1701704242
transform 1 0 19780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1701704242
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22356 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_249
timestamp 1701704242
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1701704242
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1701704242
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_305
timestamp 1701704242
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_329
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[1\].dly_stg3
timestamp 1701704242
transform 1 0 11040 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_21
timestamp 1701704242
transform -1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_22
timestamp 1701704242
transform 1 0 11592 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_23
timestamp 1701704242
transform -1 0 9108 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_24
timestamp 1701704242
transform -1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_25
timestamp 1701704242
transform -1 0 9016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[2\].dly_stg3
timestamp 1701704242
transform -1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_26
timestamp 1701704242
transform 1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_27
timestamp 1701704242
transform -1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_28
timestamp 1701704242
transform 1 0 8648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_29
timestamp 1701704242
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_30
timestamp 1701704242
transform -1 0 11040 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[3\].dly_stg3
timestamp 1701704242
transform -1 0 12144 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_31
timestamp 1701704242
transform 1 0 12420 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_32
timestamp 1701704242
transform -1 0 8280 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_33
timestamp 1701704242
transform -1 0 9292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_34
timestamp 1701704242
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_35
timestamp 1701704242
transform 1 0 9476 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[4\].dly_stg3
timestamp 1701704242
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_36
timestamp 1701704242
transform -1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_37
timestamp 1701704242
transform -1 0 10856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_38
timestamp 1701704242
transform 1 0 12512 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_39
timestamp 1701704242
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_40
timestamp 1701704242
transform -1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[5\].dly_stg3
timestamp 1701704242
transform -1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_41
timestamp 1701704242
transform -1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_42
timestamp 1701704242
transform -1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_43
timestamp 1701704242
transform 1 0 12144 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_44
timestamp 1701704242
transform -1 0 9844 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_45
timestamp 1701704242
transform 1 0 10672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[6\].dly_stg3
timestamp 1701704242
transform -1 0 12144 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_46
timestamp 1701704242
transform -1 0 12144 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_47
timestamp 1701704242
transform -1 0 8648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_48
timestamp 1701704242
transform -1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_49
timestamp 1701704242
transform 1 0 13432 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_50
timestamp 1701704242
transform 1 0 12880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[7\].dly_stg3
timestamp 1701704242
transform 1 0 13892 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_51
timestamp 1701704242
transform 1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_52
timestamp 1701704242
transform 1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_53
timestamp 1701704242
transform -1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_54
timestamp 1701704242
transform 1 0 15180 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_55
timestamp 1701704242
transform -1 0 14536 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[8\].dly_stg3
timestamp 1701704242
transform 1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_56
timestamp 1701704242
transform 1 0 18584 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_57
timestamp 1701704242
transform -1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_58
timestamp 1701704242
transform -1 0 16560 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_59
timestamp 1701704242
transform 1 0 17296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_60
timestamp 1701704242
transform -1 0 17020 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[9\].dly_stg3
timestamp 1701704242
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_61
timestamp 1701704242
transform -1 0 16560 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_62
timestamp 1701704242
transform -1 0 20332 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_63
timestamp 1701704242
transform 1 0 21436 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_64
timestamp 1701704242
transform 1 0 21712 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_65
timestamp 1701704242
transform 1 0 20608 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[10\].dly_stg3
timestamp 1701704242
transform -1 0 18492 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_66
timestamp 1701704242
transform -1 0 17388 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_67
timestamp 1701704242
transform -1 0 20608 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_68
timestamp 1701704242
transform 1 0 18676 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_69
timestamp 1701704242
transform -1 0 20240 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_70
timestamp 1701704242
transform 1 0 21988 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[11\].dly_stg3
timestamp 1701704242
transform 1 0 20700 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_71
timestamp 1701704242
transform 1 0 20700 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_72
timestamp 1701704242
transform 1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_73
timestamp 1701704242
transform -1 0 18584 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_74
timestamp 1701704242
transform -1 0 20056 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_75
timestamp 1701704242
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[12\].dly_stg3
timestamp 1701704242
transform -1 0 17940 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_76
timestamp 1701704242
transform -1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_77
timestamp 1701704242
transform 1 0 21804 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_78
timestamp 1701704242
transform 1 0 20792 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_79
timestamp 1701704242
transform 1 0 22080 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_80
timestamp 1701704242
transform 1 0 21160 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[13\].dly_stg3
timestamp 1701704242
transform -1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_81
timestamp 1701704242
transform 1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_82
timestamp 1701704242
transform -1 0 17388 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_83
timestamp 1701704242
transform -1 0 15272 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_84
timestamp 1701704242
transform -1 0 14996 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_85
timestamp 1701704242
transform 1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[14\].dly_stg3
timestamp 1701704242
transform -1 0 17204 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg4_218
timestamp 1701704242
transform 1 0 18124 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_138
timestamp 1701704242
transform -1 0 10028 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_139
timestamp 1701704242
transform -1 0 11592 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_140
timestamp 1701704242
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_141
timestamp 1701704242
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_142
timestamp 1701704242
transform -1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_143
timestamp 1701704242
transform -1 0 9936 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_144
timestamp 1701704242
transform -1 0 12144 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg8_185
timestamp 1701704242
transform -1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_94
timestamp 1701704242
transform -1 0 11960 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_95
timestamp 1701704242
transform 1 0 11684 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_96
timestamp 1701704242
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_97
timestamp 1701704242
transform -1 0 10488 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_98
timestamp 1701704242
transform 1 0 9108 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_99
timestamp 1701704242
transform -1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_100
timestamp 1701704242
transform 1 0 8556 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg8_145
timestamp 1701704242
transform 1 0 10488 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_186
timestamp 1701704242
transform 1 0 7728 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_187
timestamp 1701704242
transform -1 0 7452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_188
timestamp 1701704242
transform -1 0 11040 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_189
timestamp 1701704242
transform -1 0 9384 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_190
timestamp 1701704242
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_191
timestamp 1701704242
transform -1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_192
timestamp 1701704242
transform 1 0 8832 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg8_101
timestamp 1701704242
transform -1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_146
timestamp 1701704242
transform -1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_147
timestamp 1701704242
transform 1 0 8924 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_148
timestamp 1701704242
transform 1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_149
timestamp 1701704242
transform -1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_150
timestamp 1701704242
transform 1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_151
timestamp 1701704242
transform -1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_152
timestamp 1701704242
transform -1 0 8832 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg8_193
timestamp 1701704242
transform -1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_102
timestamp 1701704242
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_103
timestamp 1701704242
transform -1 0 10120 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_104
timestamp 1701704242
transform 1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_105
timestamp 1701704242
transform -1 0 11500 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_106
timestamp 1701704242
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_107
timestamp 1701704242
transform -1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_108
timestamp 1701704242
transform -1 0 12512 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg8_153
timestamp 1701704242
transform -1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_194
timestamp 1701704242
transform -1 0 13156 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_195
timestamp 1701704242
transform 1 0 13156 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_196
timestamp 1701704242
transform -1 0 14444 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_197
timestamp 1701704242
transform -1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_198
timestamp 1701704242
transform -1 0 13984 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_199
timestamp 1701704242
transform 1 0 14536 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_200
timestamp 1701704242
transform 1 0 11592 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg8_109
timestamp 1701704242
transform 1 0 12604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_154
timestamp 1701704242
transform 1 0 15732 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_155
timestamp 1701704242
transform 1 0 14904 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_156
timestamp 1701704242
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_157
timestamp 1701704242
transform -1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_158
timestamp 1701704242
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_159
timestamp 1701704242
transform 1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_160
timestamp 1701704242
transform 1 0 13616 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg8_201
timestamp 1701704242
transform -1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_110
timestamp 1701704242
transform 1 0 19688 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_111
timestamp 1701704242
transform 1 0 17020 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_112
timestamp 1701704242
transform -1 0 17204 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_113
timestamp 1701704242
transform -1 0 13156 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_114
timestamp 1701704242
transform 1 0 17388 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_115
timestamp 1701704242
transform 1 0 14352 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_116
timestamp 1701704242
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg8_161
timestamp 1701704242
transform -1 0 13432 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_202
timestamp 1701704242
transform 1 0 20240 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_203
timestamp 1701704242
transform 1 0 20700 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_204
timestamp 1701704242
transform 1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_205
timestamp 1701704242
transform 1 0 22080 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_206
timestamp 1701704242
transform 1 0 16284 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_207
timestamp 1701704242
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_208
timestamp 1701704242
transform -1 0 17572 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg8_117
timestamp 1701704242
transform 1 0 15180 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_162
timestamp 1701704242
transform 1 0 20332 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_163
timestamp 1701704242
transform 1 0 22356 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_164
timestamp 1701704242
transform -1 0 17756 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_165
timestamp 1701704242
transform -1 0 22448 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_166
timestamp 1701704242
transform -1 0 18124 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_167
timestamp 1701704242
transform -1 0 21436 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_168
timestamp 1701704242
transform 1 0 17940 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg8_209
timestamp 1701704242
transform 1 0 16652 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_118
timestamp 1701704242
transform 1 0 23000 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_119
timestamp 1701704242
transform -1 0 23000 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_120
timestamp 1701704242
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_121
timestamp 1701704242
transform 1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_122
timestamp 1701704242
transform 1 0 19780 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_123
timestamp 1701704242
transform 1 0 21804 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_124
timestamp 1701704242
transform -1 0 17848 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg8_169
timestamp 1701704242
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_210
timestamp 1701704242
transform 1 0 20884 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_211
timestamp 1701704242
transform 1 0 21436 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_212
timestamp 1701704242
transform 1 0 19504 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_213
timestamp 1701704242
transform 1 0 20608 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_214
timestamp 1701704242
transform -1 0 18952 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_215
timestamp 1701704242
transform 1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_216
timestamp 1701704242
transform -1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg8_125
timestamp 1701704242
transform 1 0 22448 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_170
timestamp 1701704242
transform 1 0 18676 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_171
timestamp 1701704242
transform -1 0 15548 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_172
timestamp 1701704242
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_173
timestamp 1701704242
transform -1 0 17480 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_174
timestamp 1701704242
transform 1 0 20056 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_175
timestamp 1701704242
transform -1 0 18952 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_176
timestamp 1701704242
transform -1 0 18584 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg8_217
timestamp 1701704242
transform -1 0 18952 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_126
timestamp 1701704242
transform 1 0 17848 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_127
timestamp 1701704242
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  g_dly_chain_interleave\[13\].dly_stg7_128 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16928 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_177
timestamp 1701704242
transform 1 0 16928 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_178
timestamp 1701704242
transform -1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_179
timestamp 1701704242
transform -1 0 13432 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_180
timestamp 1701704242
transform 1 0 14168 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_181
timestamp 1701704242
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[0\].dly_stp_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15180 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[1\].dly_stp_2
timestamp 1701704242
transform 1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[2\].dly_stp_3
timestamp 1701704242
transform -1 0 16928 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[3\].dly_stp_4
timestamp 1701704242
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[0\].inv_chain
timestamp 1701704242
transform -1 0 11868 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[1\].inv_chain
timestamp 1701704242
transform -1 0 11592 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[2\].inv_chain
timestamp 1701704242
transform -1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[3\].inv_chain
timestamp 1701704242
transform 1 0 10488 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1701704242
transform 1 0 12328 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 dbg_delay_stop
port 2 nsew signal tristate
flabel metal2 s 16118 19600 16174 20000 0 FreeSans 224 90 0 0 dbg_dly_sig[0]
port 3 nsew signal tristate
flabel metal2 s 21270 0 21326 400 0 FreeSans 224 90 0 0 dbg_dly_sig[10]
port 4 nsew signal tristate
flabel metal2 s 19982 0 20038 400 0 FreeSans 224 90 0 0 dbg_dly_sig[11]
port 5 nsew signal tristate
flabel metal2 s 19338 0 19394 400 0 FreeSans 224 90 0 0 dbg_dly_sig[12]
port 6 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 dbg_dly_sig[13]
port 7 nsew signal tristate
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 dbg_dly_sig[14]
port 8 nsew signal tristate
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 dbg_dly_sig[15]
port 9 nsew signal tristate
flabel metal2 s 10322 0 10378 400 0 FreeSans 224 90 0 0 dbg_dly_sig[1]
port 10 nsew signal tristate
flabel metal3 s 0 10208 400 10328 0 FreeSans 480 0 0 0 dbg_dly_sig[2]
port 11 nsew signal tristate
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 dbg_dly_sig[3]
port 12 nsew signal tristate
flabel metal3 s 0 8848 400 8968 0 FreeSans 480 0 0 0 dbg_dly_sig[4]
port 13 nsew signal tristate
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 dbg_dly_sig[5]
port 14 nsew signal tristate
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 dbg_dly_sig[6]
port 15 nsew signal tristate
flabel metal2 s 12898 0 12954 400 0 FreeSans 224 90 0 0 dbg_dly_sig[7]
port 16 nsew signal tristate
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 dbg_dly_sig[8]
port 17 nsew signal tristate
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 dbg_dly_sig[9]
port 18 nsew signal tristate
flabel metal2 s 14186 19600 14242 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[0]
port 19 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[1]
port 20 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[2]
port 21 nsew signal tristate
flabel metal3 s 0 11568 400 11688 0 FreeSans 480 0 0 0 dbg_start_pulse
port 22 nsew signal tristate
flabel metal2 s 12254 19600 12310 20000 0 FreeSans 224 90 0 0 i_start
port 23 nsew signal input
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 i_stop
port 24 nsew signal input
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 o_result_ctr[0]
port 25 nsew signal tristate
flabel metal3 s 31600 10888 32000 11008 0 FreeSans 480 0 0 0 o_result_ctr[1]
port 26 nsew signal tristate
flabel metal2 s 20626 19600 20682 20000 0 FreeSans 224 90 0 0 o_result_ctr[2]
port 27 nsew signal tristate
flabel metal2 s 15474 19600 15530 20000 0 FreeSans 224 90 0 0 o_result_ring[0]
port 28 nsew signal tristate
flabel metal2 s 20626 0 20682 400 0 FreeSans 224 90 0 0 o_result_ring[10]
port 29 nsew signal tristate
flabel metal3 s 31600 8168 32000 8288 0 FreeSans 480 0 0 0 o_result_ring[11]
port 30 nsew signal tristate
flabel metal3 s 31600 8848 32000 8968 0 FreeSans 480 0 0 0 o_result_ring[12]
port 31 nsew signal tristate
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 o_result_ring[13]
port 32 nsew signal tristate
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 o_result_ring[14]
port 33 nsew signal tristate
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 o_result_ring[15]
port 34 nsew signal tristate
flabel metal2 s 13542 19600 13598 20000 0 FreeSans 224 90 0 0 o_result_ring[1]
port 35 nsew signal tristate
flabel metal3 s 0 10888 400 11008 0 FreeSans 480 0 0 0 o_result_ring[2]
port 36 nsew signal tristate
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 o_result_ring[3]
port 37 nsew signal tristate
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 o_result_ring[4]
port 38 nsew signal tristate
flabel metal3 s 0 7488 400 7608 0 FreeSans 480 0 0 0 o_result_ring[5]
port 39 nsew signal tristate
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 o_result_ring[6]
port 40 nsew signal tristate
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 o_result_ring[7]
port 41 nsew signal tristate
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 o_result_ring[8]
port 42 nsew signal tristate
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 o_result_ring[9]
port 43 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal1 13370 12342 13370 12342 0 _00_
rlabel metal1 15124 11662 15124 11662 0 _01_
rlabel metal2 17526 12517 17526 12517 0 _02_
rlabel metal1 12466 11288 12466 11288 0 _03_
rlabel metal1 12512 11866 12512 11866 0 _04_
rlabel metal1 13340 11866 13340 11866 0 _05_
rlabel metal1 15180 11594 15180 11594 0 _06_
rlabel metal1 17204 11866 17204 11866 0 _07_
rlabel metal1 17404 11594 17404 11594 0 _08_
rlabel metal2 17342 12308 17342 12308 0 _09_
rlabel metal1 14444 9146 14444 9146 0 clknet_0_i_stop
rlabel metal1 15916 9350 15916 9350 0 clknet_0_net5
rlabel metal1 14260 7990 14260 7990 0 clknet_1_0__leaf_i_stop
rlabel metal1 12604 7310 12604 7310 0 clknet_1_0__leaf_net5
rlabel metal1 16790 7378 16790 7378 0 clknet_1_1__leaf_i_stop
rlabel metal3 15617 8228 15617 8228 0 clknet_1_1__leaf_net5
rlabel metal2 14398 5831 14398 5831 0 dbg_delay_stop
rlabel metal2 16192 19244 16192 19244 0 dbg_dly_sig[0]
rlabel metal1 20884 7786 20884 7786 0 dbg_dly_sig[10]
rlabel metal3 19274 8364 19274 8364 0 dbg_dly_sig[11]
rlabel metal2 19642 9418 19642 9418 0 dbg_dly_sig[12]
rlabel metal1 21942 9656 21942 9656 0 dbg_dly_sig[13]
rlabel metal1 16054 9894 16054 9894 0 dbg_dly_sig[14]
rlabel metal2 14858 5124 14858 5124 0 dbg_dly_sig[15]
rlabel metal4 14076 6868 14076 6868 0 dbg_dly_sig[1]
rlabel metal3 1533 10268 1533 10268 0 dbg_dly_sig[2]
rlabel metal2 12282 619 12282 619 0 dbg_dly_sig[3]
rlabel metal3 4638 8908 4638 8908 0 dbg_dly_sig[4]
rlabel metal3 1533 8228 1533 8228 0 dbg_dly_sig[5]
rlabel metal1 11132 7718 11132 7718 0 dbg_dly_sig[6]
rlabel metal2 12926 1557 12926 1557 0 dbg_dly_sig[7]
rlabel metal1 15180 7174 15180 7174 0 dbg_dly_sig[8]
rlabel metal1 17250 7718 17250 7718 0 dbg_dly_sig[9]
rlabel metal1 14030 11322 14030 11322 0 dbg_ring_ctr[0]
rlabel metal1 18538 12342 18538 12342 0 dbg_ring_ctr[1]
rlabel metal1 19550 12410 19550 12410 0 dbg_ring_ctr[2]
rlabel metal1 11776 11254 11776 11254 0 dbg_start_pulse
rlabel metal1 12328 18802 12328 18802 0 i_start
rlabel metal4 13892 5916 13892 5916 0 i_stop
rlabel metal1 12604 11662 12604 11662 0 net1
rlabel metal1 10994 6188 10994 6188 0 net10
rlabel metal1 10902 10710 10902 10710 0 net100
rlabel metal2 8694 10676 8694 10676 0 net101
rlabel metal2 8142 9894 8142 9894 0 net102
rlabel metal1 10442 6222 10442 6222 0 net103
rlabel viali 9798 7311 9798 7311 0 net104
rlabel metal3 11753 7820 11753 7820 0 net105
rlabel metal1 11178 6426 11178 6426 0 net106
rlabel metal1 13110 6188 13110 6188 0 net107
rlabel metal1 12604 6222 12604 6222 0 net108
rlabel metal1 11730 5338 11730 5338 0 net109
rlabel metal1 9614 11050 9614 11050 0 net11
rlabel metal2 12742 6817 12742 6817 0 net110
rlabel metal1 16974 6290 16974 6290 0 net111
rlabel metal1 17250 6222 17250 6222 0 net112
rlabel metal1 16514 7956 16514 7956 0 net113
rlabel metal1 12788 8058 12788 8058 0 net114
rlabel metal1 18630 6766 18630 6766 0 net115
rlabel metal1 15226 7854 15226 7854 0 net116
rlabel metal1 15088 6630 15088 6630 0 net117
rlabel metal1 16330 6154 16330 6154 0 net118
rlabel metal1 23230 9486 23230 9486 0 net119
rlabel metal1 10810 5746 10810 5746 0 net12
rlabel metal2 22126 9367 22126 9367 0 net120
rlabel metal2 21482 10574 21482 10574 0 net121
rlabel metal2 18998 7140 18998 7140 0 net122
rlabel metal1 20332 10098 20332 10098 0 net123
rlabel metal1 22494 9520 22494 9520 0 net124
rlabel metal1 19274 8058 19274 8058 0 net125
rlabel metal2 22586 9248 22586 9248 0 net126
rlabel metal1 18078 10574 18078 10574 0 net127
rlabel metal2 16698 9520 16698 9520 0 net128
rlabel metal1 12190 9044 12190 9044 0 net129
rlabel metal2 8970 10370 8970 10370 0 net13
rlabel metal1 11362 9452 11362 9452 0 net130
rlabel via2 10166 9469 10166 9469 0 net132
rlabel metal1 16514 11254 16514 11254 0 net133
rlabel metal1 14623 11254 14623 11254 0 net134
rlabel metal1 16974 11696 16974 11696 0 net135
rlabel metal1 15640 12206 15640 12206 0 net136
rlabel metal1 13892 11798 13892 11798 0 net137
rlabel metal1 12190 11696 12190 11696 0 net138
rlabel metal2 9706 10880 9706 10880 0 net139
rlabel via1 11270 11185 11270 11185 0 net14
rlabel metal1 10534 11220 10534 11220 0 net140
rlabel metal1 10580 12138 10580 12138 0 net141
rlabel metal1 11546 9554 11546 9554 0 net142
rlabel metal1 8510 8942 8510 8942 0 net143
rlabel metal2 10534 9316 10534 9316 0 net144
rlabel metal1 11408 11322 11408 11322 0 net145
rlabel metal2 10626 9537 10626 9537 0 net146
rlabel metal1 8464 8058 8464 8058 0 net147
rlabel metal1 10074 6868 10074 6868 0 net148
rlabel metal1 12466 7378 12466 7378 0 net149
rlabel metal2 16974 9622 16974 9622 0 net15
rlabel metal1 11546 6426 11546 6426 0 net150
rlabel metal1 12282 6256 12282 6256 0 net151
rlabel metal1 9614 7446 9614 7446 0 net152
rlabel metal2 7958 9520 7958 9520 0 net153
rlabel metal1 8602 6834 8602 6834 0 net154
rlabel metal1 15180 6086 15180 6086 0 net155
rlabel metal1 15134 6222 15134 6222 0 net156
rlabel metal1 16054 6698 16054 6698 0 net157
rlabel metal1 11638 6800 11638 6800 0 net158
rlabel metal1 14490 8806 14490 8806 0 net159
rlabel metal2 17894 7582 17894 7582 0 net16
rlabel metal1 13340 7514 13340 7514 0 net160
rlabel metal2 14122 6018 14122 6018 0 net161
rlabel metal1 13018 7990 13018 7990 0 net162
rlabel metal1 21252 7514 21252 7514 0 net163
rlabel metal1 20194 6766 20194 6766 0 net164
rlabel metal1 18722 8466 18722 8466 0 net165
rlabel metal1 20562 10540 20562 10540 0 net166
rlabel metal1 17342 6800 17342 6800 0 net167
rlabel metal1 19366 6800 19366 6800 0 net168
rlabel metal1 18170 6086 18170 6086 0 net169
rlabel metal1 17710 6188 17710 6188 0 net17
rlabel metal1 19320 6970 19320 6970 0 net170
rlabel metal1 19090 10574 19090 10574 0 net171
rlabel metal1 14950 10608 14950 10608 0 net172
rlabel metal1 15226 10540 15226 10540 0 net173
rlabel metal2 17342 9452 17342 9452 0 net174
rlabel metal1 21850 9486 21850 9486 0 net175
rlabel metal1 16974 11220 16974 11220 0 net176
rlabel metal1 18216 6630 18216 6630 0 net177
rlabel metal1 13478 7854 13478 7854 0 net179
rlabel metal1 21068 9010 21068 9010 0 net18
rlabel metal1 12282 10064 12282 10064 0 net180
rlabel metal1 14536 10166 14536 10166 0 net181
rlabel metal1 16054 10166 16054 10166 0 net182
rlabel metal2 12926 11424 12926 11424 0 net183
rlabel metal1 13110 10132 13110 10132 0 net184
rlabel metal1 10396 9690 10396 9690 0 net185
rlabel metal2 11730 10880 11730 10880 0 net186
rlabel metal1 8234 9622 8234 9622 0 net187
rlabel metal1 8694 6902 8694 6902 0 net188
rlabel metal1 9246 10608 9246 10608 0 net189
rlabel metal1 18262 6256 18262 6256 0 net19
rlabel metal1 8556 9962 8556 9962 0 net190
rlabel metal1 12374 5746 12374 5746 0 net191
rlabel metal1 10948 6630 10948 6630 0 net192
rlabel metal1 10856 5882 10856 5882 0 net193
rlabel metal1 10074 6630 10074 6630 0 net194
rlabel metal1 12972 5134 12972 5134 0 net195
rlabel metal1 13386 5746 13386 5746 0 net196
rlabel metal1 13800 6358 13800 6358 0 net197
rlabel metal1 8602 8364 8602 8364 0 net198
rlabel metal1 13524 7446 13524 7446 0 net199
rlabel metal1 14605 8058 14605 8058 0 net2
rlabel metal1 14260 6970 14260 6970 0 net20
rlabel metal1 14628 6426 14628 6426 0 net200
rlabel metal1 11822 6970 11822 6970 0 net201
rlabel metal1 11638 6698 11638 6698 0 net202
rlabel metal1 20516 6970 20516 6970 0 net203
rlabel metal1 21298 7854 21298 7854 0 net204
rlabel metal1 20516 6630 20516 6630 0 net205
rlabel metal3 21068 7140 21068 7140 0 net206
rlabel metal1 16468 6222 16468 6222 0 net207
rlabel metal2 16698 7548 16698 7548 0 net208
rlabel metal1 16560 8058 16560 8058 0 net209
rlabel metal1 15962 8398 15962 8398 0 net21
rlabel metal1 17158 6970 17158 6970 0 net210
rlabel metal1 21114 10574 21114 10574 0 net211
rlabel metal1 21574 10200 21574 10200 0 net212
rlabel metal1 20792 9486 20792 9486 0 net213
rlabel metal1 21850 9044 21850 9044 0 net214
rlabel metal1 17434 8500 17434 8500 0 net215
rlabel metal1 20102 12750 20102 12750 0 net216
rlabel metal2 17802 7353 17802 7353 0 net217
rlabel metal1 20424 12614 20424 12614 0 net218
rlabel metal2 18262 11050 18262 11050 0 net219
rlabel metal1 11178 6732 11178 6732 0 net22
rlabel metal1 14536 9690 14536 9690 0 net220
rlabel metal1 9062 9622 9062 9622 0 net24
rlabel metal1 11132 10098 11132 10098 0 net25
rlabel metal1 9092 10166 9092 10166 0 net26
rlabel metal1 10166 10506 10166 10506 0 net27
rlabel metal1 12098 5780 12098 5780 0 net29
rlabel metal1 15226 8500 15226 8500 0 net3
rlabel metal1 13110 8602 13110 8602 0 net30
rlabel metal1 13744 8398 13744 8398 0 net31
rlabel metal1 9338 7344 9338 7344 0 net32
rlabel metal1 7820 9010 7820 9010 0 net34
rlabel metal1 9936 6834 9936 6834 0 net35
rlabel metal1 9563 9010 9563 9010 0 net36
rlabel metal1 10442 8466 10442 8466 0 net37
rlabel metal2 12650 5848 12650 5848 0 net39
rlabel metal1 15525 8602 15525 8602 0 net4
rlabel metal1 10212 6834 10212 6834 0 net40
rlabel metal1 9046 7990 9046 7990 0 net41
rlabel metal1 13064 7310 13064 7310 0 net42
rlabel metal1 12098 6868 12098 6868 0 net44
rlabel metal1 10074 7514 10074 7514 0 net45
rlabel metal2 10810 6834 10810 6834 0 net46
rlabel metal1 17572 6834 17572 6834 0 net47
rlabel metal2 12558 8772 12558 8772 0 net49
rlabel metal1 14559 9418 14559 9418 0 net5
rlabel metal1 13294 5882 13294 5882 0 net50
rlabel metal1 12972 5338 12972 5338 0 net51
rlabel metal1 21528 8806 21528 8806 0 net52
rlabel metal1 14766 6834 14766 6834 0 net54
rlabel metal2 15318 6800 15318 6800 0 net55
rlabel metal1 14950 6698 14950 6698 0 net56
rlabel metal1 18078 6222 18078 6222 0 net57
rlabel metal1 15502 7820 15502 7820 0 net59
rlabel metal1 15686 7956 15686 7956 0 net6
rlabel metal1 17296 6426 17296 6426 0 net60
rlabel metal1 16928 6426 16928 6426 0 net61
rlabel metal1 17802 7956 17802 7956 0 net63
rlabel metal1 20010 6222 20010 6222 0 net64
rlabel metal1 20194 7990 20194 7990 0 net65
rlabel metal1 20102 7446 20102 7446 0 net66
rlabel metal1 18676 11186 18676 11186 0 net68
rlabel metal2 18814 8772 18814 8772 0 net69
rlabel metal1 15318 6426 15318 6426 0 net7
rlabel metal1 18538 8330 18538 8330 0 net70
rlabel metal1 20470 8500 20470 8500 0 net71
rlabel metal1 18722 9486 18722 9486 0 net72
rlabel metal1 17894 6256 17894 6256 0 net74
rlabel metal1 20010 7514 20010 7514 0 net75
rlabel metal1 20051 9010 20051 9010 0 net76
rlabel metal1 16836 10098 16836 10098 0 net77
rlabel metal1 18216 6834 18216 6834 0 net79
rlabel metal1 14076 5746 14076 5746 0 net8
rlabel metal1 21344 9418 21344 9418 0 net80
rlabel metal1 20419 10166 20419 10166 0 net81
rlabel metal1 17204 9146 17204 9146 0 net83
rlabel metal1 14030 7922 14030 7922 0 net84
rlabel metal1 15318 10200 15318 10200 0 net85
rlabel metal1 18487 10098 18487 10098 0 net86
rlabel metal2 13754 10370 13754 10370 0 net87
rlabel metal1 13754 8058 13754 8058 0 net88
rlabel metal1 12328 8398 12328 8398 0 net89
rlabel metal2 12282 6970 12282 6970 0 net9
rlabel metal2 11868 7684 11868 7684 0 net90
rlabel metal1 11086 11254 11086 11254 0 net91
rlabel metal1 12926 9962 12926 9962 0 net92
rlabel metal1 13938 10166 13938 10166 0 net93
rlabel metal1 11760 10506 11760 10506 0 net94
rlabel metal1 11408 9146 11408 9146 0 net95
rlabel metal1 12696 8398 12696 8398 0 net96
rlabel metal1 8694 8466 8694 8466 0 net97
rlabel metal1 9614 9452 9614 9452 0 net98
rlabel metal1 9338 9622 9338 9622 0 net99
rlabel metal1 18814 10778 18814 10778 0 o_result_ctr[0]
rlabel metal1 24564 11050 24564 11050 0 o_result_ctr[1]
rlabel metal1 20746 11866 20746 11866 0 o_result_ctr[2]
rlabel metal2 15502 18099 15502 18099 0 o_result_ring[0]
rlabel metal2 20562 6619 20562 6619 0 o_result_ring[10]
rlabel metal1 21666 8364 21666 8364 0 o_result_ring[11]
rlabel via2 28290 8891 28290 8891 0 o_result_ring[12]
rlabel via2 31694 10251 31694 10251 0 o_result_ring[13]
rlabel metal2 19734 19652 19734 19652 0 o_result_ring[14]
rlabel metal2 17480 11492 17480 11492 0 o_result_ring[15]
rlabel metal2 13570 18099 13570 18099 0 o_result_ring[1]
rlabel metal3 1533 10948 1533 10948 0 o_result_ring[2]
rlabel metal3 15341 8364 15341 8364 0 o_result_ring[3]
rlabel metal2 11178 9197 11178 9197 0 o_result_ring[4]
rlabel metal3 1533 7548 1533 7548 0 o_result_ring[5]
rlabel metal1 12006 7786 12006 7786 0 o_result_ring[6]
rlabel metal1 13754 7242 13754 7242 0 o_result_ring[7]
rlabel metal2 16882 6109 16882 6109 0 o_result_ring[8]
rlabel metal2 18906 6347 18906 6347 0 o_result_ring[9]
rlabel metal1 18722 10574 18722 10574 0 r_dly_store_ctr\[0\]
rlabel metal1 20562 11288 20562 11288 0 r_dly_store_ctr\[1\]
rlabel metal1 20654 11594 20654 11594 0 r_dly_store_ctr\[2\]
rlabel metal1 15502 11254 15502 11254 0 r_dly_store_ring\[0\]
rlabel metal1 20194 7922 20194 7922 0 r_dly_store_ring\[10\]
rlabel metal1 20654 8398 20654 8398 0 r_dly_store_ring\[11\]
rlabel metal1 21390 8976 21390 8976 0 r_dly_store_ring\[12\]
rlabel metal1 21390 10200 21390 10200 0 r_dly_store_ring\[13\]
rlabel metal1 19182 9486 19182 9486 0 r_dly_store_ring\[14\]
rlabel metal1 17434 10472 17434 10472 0 r_dly_store_ring\[15\]
rlabel metal1 13662 10472 13662 10472 0 r_dly_store_ring\[1\]
rlabel metal1 10948 10234 10948 10234 0 r_dly_store_ring\[2\]
rlabel metal1 15042 8398 15042 8398 0 r_dly_store_ring\[3\]
rlabel metal1 10856 9078 10856 9078 0 r_dly_store_ring\[4\]
rlabel metal2 10626 8194 10626 8194 0 r_dly_store_ring\[5\]
rlabel metal1 12236 7446 12236 7446 0 r_dly_store_ring\[6\]
rlabel metal1 14076 6698 14076 6698 0 r_dly_store_ring\[7\]
rlabel metal1 16652 6902 16652 6902 0 r_dly_store_ring\[8\]
rlabel metal1 18814 7208 18814 7208 0 r_dly_store_ring\[9\]
rlabel metal1 13846 11594 13846 11594 0 r_ring_ctr\[0\]
rlabel via1 19269 11254 19269 11254 0 r_ring_ctr\[1\]
rlabel metal1 17710 11730 17710 11730 0 r_ring_ctr\[2\]
rlabel metal1 11597 12274 11597 12274 0 w_dly_strt_ana_\[1\]
rlabel metal1 10838 11186 10838 11186 0 w_dly_strt_ana_\[2\]
rlabel via1 10649 11322 10649 11322 0 w_dly_strt_ana_\[3\]
rlabel metal2 12834 11458 12834 11458 0 w_dly_strt_ana_\[4\]
rlabel metal1 14904 11662 14904 11662 0 w_ring_ctr_clk
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
