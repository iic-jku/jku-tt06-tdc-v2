* PEX produced on Fri Mar 29 11:41:37 PM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tt_um_hpretl_tt06_tdc_v2.ext - technology: sky130A

.subckt tt_um_hpretl_tt06_tdc_v2 clk ena rst_n ui_in[3] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[7] uio_out[3] uo_out[0] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] ui_in[0] ui_in[2] uio_oe[0] ui_in[4] uio_out[2] uo_out[1] uio_out[0] uio_oe[5]
+ uio_oe[4] uio_out[7] uio_out[1] uio_out[6] uio_oe[1] uio_oe[6] uio_out[5] uio_oe[2]
+ uio_oe[3] uio_out[4] ui_in[1] VPWR VGND
X0 VGND a_7902_8725# a_7860_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1 a_12150_10749# a_11877_10383# a_12065_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3 VGND _078_ _079_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.172 ps=1.83 w=0.65 l=0.15
X4 _150_ a_9167_14763# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X6 a_17751_3829# a_17576_3855# a_17930_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7 a_26969_9839# tdc1.w_ring_buf[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND a_3439_14191# _003_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X11 tdc1.r_dly_store_ring[21] a_15871_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_9577_10933# a_9411_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_14421_15823# a_14377_16065# a_14255_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X14 a_16477_15823# a_16311_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_9008_15279# _148_ a_8543_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X16 a_23834_14191# a_23395_14197# a_23749_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X18 VPWR net32 a_21647_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X19 a_12813_3311# _175_ a_12731_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_7223_9813# a_7139_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X22 VPWR a_2932_14165# net27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X23 a_29035_7663# a_28253_7669# a_28951_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X25 a_15703_7485# a_15005_7119# a_15446_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X26 VPWR a_17895_5461# a_17811_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 VGND a_9447_5309# a_9615_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 tdc1.g_ring3[25].stg01_70.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X28 a_27065_6575# net40 tdc1.w_ring_int_norsz[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X30 VGND tdc0.w_ring_buf[0] a_18059_16375# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X31 a_6357_12559# a_6191_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X33 VGND net26 a_3247_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X34 a_4595_6005# a_4420_6031# a_4774_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X36 a_11115_4007# tdc1.r_ring_ctr[6] a_11349_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X37 VPWR a_19805_3285# a_19695_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X38 a_21997_5493# a_21831_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X40 a_19237_6281# tdc1.w_ring_norsz[13] a_19153_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X42 a_21361_7369# _075_ a_21445_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X43 VGND a_28951_9839# a_29119_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R1 net51 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X44 a_26479_11159# a_26575_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X45 VPWR a_17475_13621# a_17482_13921# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X46 a_28331_12233# net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X47 a_24420_12393# a_24021_12021# a_24294_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X48 VPWR _072_ a_11233_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X49 VPWR tdc1.r_ring_ctr[4] a_12139_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 VPWR a_14342_10901# a_14269_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X51 VGND _095_ a_25973_9301# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X52 VGND tdc0.w_ring_norsz[24] a_9135_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X54 VPWR a_19692_4777# a_19867_4703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X56 VGND _138_ a_10946_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X57 a_22163_14735# a_21647_14735# a_22068_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X59 a_17100_4765# _017_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X60 VPWR net30 a_11619_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X61 VPWR tdc1.r_ring_ctr[12] a_6373_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X62 a_22649_4399# _167_ _025_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X64 net15 a_9103_4659# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X65 VGND a_22903_14709# a_22837_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X66 a_20533_6575# _077_ a_20617_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X67 VPWR a_5951_7485# a_6119_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
R2 VGND uio_out[7] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X68 VGND net7 a_10975_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X70 _066_ a_15335_8181# a_15283_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 net11 a_5271_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X74 VGND tdc0.w_dly_stop[1] a_2603_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X75 VPWR a_12594_7637# a_12521_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X78 a_8270_7637# a_8102_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
R3 VGND net61 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X80 a_17221_6575# net67 tdc1.w_ring_int_norsz[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X81 a_9785_15645# _143_ a_9713_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X82 a_11693_7663# tdc1.w_ring_norsz[23] a_11609_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X83 VPWR a_24151_9813# a_24067_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X84 VPWR a_20810_13621# a_20739_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X85 VPWR net5 a_16771_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X86 tdc1.w_ring_norsz[25] net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X87 a_30101_8751# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X88 VGND a_8159_8751# a_8327_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X89 a_19345_4373# a_19127_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X90 VPWR net9 a_11619_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X91 VPWR a_25071_6549# a_24987_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X92 a_24294_15101# a_23855_14735# a_24209_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X93 tdc1.w_dly_stop[1] a_26615_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X94 VGND tdc0.w_ring_norsz[16] a_4627_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X95 VPWR net10 a_21831_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X96 net21 a_3484_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X97 a_23565_13103# tdc0.w_ring_buf[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X98 a_11809_15279# _146_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X99 a_14008_9545# _193_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X100 a_12729_11721# tdc0.w_ring_norsz[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X102 tdc1.w_ring_norsz[5] tdc1.w_ring_norsz[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 a_10291_4373# _179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X105 VPWR a_29035_9447# _096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X106 tdc1.r_ring_ctr[10] a_17935_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X107 VPWR a_20152_3689# a_20327_3615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X108 a_11792_12015# _130_ a_11623_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X110 VGND net39 tdc0.w_ring_int_norsz[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R4 VPWR tdc1.g_ring3[23].stg01_68.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X111 VPWR _066_ a_11987_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X112 VGND net13 a_7571_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X113 VGND net28 a_6191_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X114 VGND _196_ _049_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X115 a_25511_10927# _083_ a_25689_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X117 a_17417_11721# tdc0.w_ring_int_norsz[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X118 VPWR a_7364_14569# a_7539_14495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 a_5560_13647# a_5161_13647# a_5434_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X120 a_19142_10749# a_18703_10383# a_19057_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X121 a_7274_6397# a_6835_6031# a_7189_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X122 tdc0.w_ring_norsz[20] net24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X125 a_3115_9813# net28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X126 tdc0.r_dly_store_ring[16] a_5935_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X127 VGND a_22254_13759# a_22212_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X128 a_22833_11721# net22 tdc0.w_ring_norsz[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X131 tdc0.r_dly_store_ctr[9] a_19735_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X132 tdc1.w_ring_norsz[28] net18 a_26149_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X133 VGND tdc1.w_ring_int_norsz[20] tdc1.w_ring_norsz[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X134 a_17746_15823# _041_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X136 VPWR net32 a_19623_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X137 a_29035_9447# tdc1.r_dly_store_ring[10] a_29181_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X138 VPWR tdc0.w_ring_int_norsz[5] a_16385_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X139 uo_out[4] a_21912_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X140 a_26513_13423# tdc0.r_dly_store_ring[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X141 VGND _070_ _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X142 VGND net16 tdc1.w_ring_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X143 a_7783_6397# a_7001_6031# a_7699_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X144 VPWR a_17746_8319# a_17673_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X145 VGND net36 a_29007_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X148 _023_ a_20735_3017# a_20985_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X149 a_12521_7663# a_11987_7669# a_12426_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X150 tdc0.w_ring_buf[25] a_17875_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X151 a_2894_10927# a_2768_11043# a_2490_11059# VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X152 tdc0.w_ring_int_norsz[7] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X153 a_27491_5108# tdc1.w_dly_stop[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X156 tdc1.r_dly_store_ctr[4] a_25899_4123# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X157 a_15256_10535# _116_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X160 tdc0.w_ring_int_norsz[17] net44 a_4725_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X161 VGND net30 a_10055_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X162 VPWR net7 a_10975_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X164 a_15539_13647# a_15023_13647# a_15444_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X165 a_14431_4373# tdc1.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X166 VGND net28 a_8399_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X167 VGND a_11792_12015# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X169 VGND _044_ a_4577_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X170 VGND net33 a_21739_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X171 VGND a_8235_13077# a_8193_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X172 VPWR tdc0.w_ring_norsz[3] a_23201_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X173 VPWR a_11950_14165# a_11877_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X174 VGND tdc0.w_ring_norsz[26] a_19255_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X176 VGND a_30039_7387# a_29997_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X177 a_14090_9295# _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X178 VPWR tdc0.w_ring_norsz[10] a_24775_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X179 VGND net8 a_16495_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X180 VGND net41 tdc0.w_ring_int_norsz[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X181 a_2840_12533# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X182 a_20985_3017# tdc1.r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R5 VPWR tdc0.g_ring3[25].stg01_52.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X184 VPWR _150_ a_9647_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X185 a_3484_13077# net24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X186 VPWR tdc1.w_ring_norsz[4] a_18785_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X187 tdc1.w_ring_buf[17] a_23855_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X188 VGND tdc1.w_ring_norsz[12] tdc1.w_ring_norsz[28] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X189 a_18605_8029# a_18335_7663# a_18501_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X190 a_15701_8457# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X191 VGND _070_ a_18243_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X192 a_19315_15823# a_18869_15823# a_19219_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X193 a_21095_12559# _088_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X195 VPWR _195_ _037_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X196 a_28885_12393# a_28338_12137# a_28538_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X197 VPWR tdc0.w_ring_int_norsz[12] a_19881_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X198 VGND _075_ a_12793_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X199 a_25864_8457# _100_ a_25609_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X200 tdc1.r_dly_store_ring[0] a_4279_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X201 VGND net7 a_19071_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X203 a_7649_8751# tdc1.w_ring_buf[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X205 VPWR a_8527_7663# a_8695_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X206 VGND a_5507_6005# _184_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X207 VGND _126_ a_11713_6691# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X208 a_21729_12015# net24 tdc0.w_ring_norsz[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X209 a_19805_3285# a_19587_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X210 VGND net34 a_23487_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X211 VPWR a_28538_12292# a_28467_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X212 VGND tdc0.w_ring_norsz[11] tdc0.w_ring_int_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X213 a_7400_6031# a_7001_6031# a_7274_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X214 net7 a_6980_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X215 a_16826_9813# a_16658_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X216 VPWR _038_ a_8451_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X218 a_23021_8457# tdc1.w_ring_norsz[17] a_22937_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R6 tt_um_hpretl_tt06_tdc_v2_78.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X220 _080_ a_19631_8867# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X221 tdc0.r_dly_store_ring[2] a_24887_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X222 _039_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X225 a_17673_8573# a_17139_8207# a_17578_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X226 VPWR a_25071_10901# a_24987_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X227 a_19805_15279# tdc0.r_ring_ctr[1] a_19723_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X228 a_26701_8751# tdc1.w_ring_norsz[9] a_26617_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X229 a_19034_10901# a_18866_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X230 tdc0.r_dly_store_ring[2] a_24887_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X232 a_7275_15279# _039_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X233 a_15703_7485# a_14839_7119# a_15446_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X234 a_8573_6575# net38 tdc1.w_ring_int_norsz[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X235 VGND a_11655_6397# a_11823_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X236 net17 a_27036_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X238 a_12077_16341# a_11859_16745# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X239 VGND a_24887_11989# a_24845_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X240 _099_ a_18501_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X241 a_10309_5807# tdc1.r_dly_store_ring[30] a_9963_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X242 a_15333_9545# _121_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X243 VPWR net20 _046_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X244 a_3871_12925# _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X245 tdc1.w_ring_norsz[16] net15 a_6813_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X248 a_23074_15279# a_21997_15285# a_22912_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X249 VPWR a_22926_10357# a_22855_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X250 a_15627_14709# tdc0.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X251 VPWR tdc1.r_ring_ctr[1] a_21279_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X253 tdc0.r_dly_store_ctr[3] a_24887_15003# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X254 VPWR tdc1.w_ring_norsz[20] a_22741_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X255 a_4582_6397# a_3505_6031# a_4420_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X256 VPWR net23 a_19255_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X257 tdc0.w_ring_int_norsz[16] tdc0.w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X260 VGND net61 tdc1.w_ring_int_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X261 VPWR a_17323_8759# net31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X265 a_11509_16373# a_11343_16373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X266 _090_ a_21095_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.26 ps=1.45 w=0.65 l=0.15
X269 a_14442_9295# _193_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X270 a_22070_15823# _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X273 VGND a_28694_7637# a_28652_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X274 a_9240_13481# a_8841_13109# a_9114_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X275 VGND a_17923_12234# tdc0.w_ring_buf[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X276 a_12337_4405# a_12171_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X277 a_17627_9661# a_16845_9295# a_17543_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X278 a_9103_4659# net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X279 a_19715_14985# tdc0.r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X280 VGND a_17682_13621# a_17611_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X281 a_8193_13481# a_7203_13109# a_8067_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X283 a_29614_7231# a_29446_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X286 VPWR a_15627_14709# _155_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X287 _103_ a_23947_12809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X288 VPWR net8 a_16495_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X289 a_4073_6273# a_3855_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X290 a_8527_7663# a_7663_7669# a_8270_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X291 VGND net32 a_21647_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X292 a_7810_13077# a_7642_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X293 VPWR tdc1.w_ring_norsz[19] a_23855_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X294 tdc0.r_dly_store_ring[28] a_19459_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X295 a_29614_7231# a_29446_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X296 _065_ a_16771_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X297 _187_ a_12815_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X298 VPWR net9 a_18703_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X299 uo_out[2] a_26420_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X300 VPWR a_10443_11989# a_10359_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X301 VGND net22 a_18703_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X302 a_6357_12559# a_6191_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X303 VGND _039_ a_7429_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X304 a_25765_5865# a_24775_5493# a_25639_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X305 VPWR a_25899_13077# a_25815_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X307 a_12231_14735# a_11785_14735# a_12135_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X308 a_7642_13103# a_7369_13109# a_7557_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X309 VPWR a_19291_10927# a_19459_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X310 VGND _040_ a_14421_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X311 VPWR _092_ a_26506_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X312 a_20152_3689# a_19071_3317# a_19805_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X313 a_9298_8573# a_9025_8207# a_9213_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X314 a_26597_12021# a_26431_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 net24 a_3799_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X317 a_23166_4221# a_22089_3855# a_23004_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X318 VGND a_25347_7637# a_25305_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R7 tdc0.g_ring3[17].stg01_44.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X319 VPWR a_27066_11204# a_26995_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X320 a_10229_13103# tdc0.r_dly_store_ring[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X321 VGND a_17475_13621# a_17482_13921# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X322 VGND a_18003_8573# a_18171_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X323 a_12318_10495# a_12150_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X326 a_22438_5461# a_22270_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X327 a_19567_14013# a_18703_13647# a_19310_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X329 VGND tdc0.r_ring_ctr[14] _162_ VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.106 ps=0.975 w=0.65 l=0.15
X330 a_4025_7119# a_3981_7361# a_3859_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X332 a_20319_13621# a_20603_13621# a_20538_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X333 VGND tdc1.w_ring_norsz[31] tdc1.w_ring_int_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X334 tdc0.w_ring_int_norsz[16] net38 a_6749_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X335 a_20847_11837# a_20065_11471# a_20763_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X336 a_20487_12925# a_19789_12559# a_20230_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X337 a_5161_13647# a_4995_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X338 VPWR net10 a_17415_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X340 tdc0.w_ring_norsz[10] net22 a_19065_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X341 a_19237_14013# a_18703_13647# a_19142_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X342 a_26593_6031# tdc1.r_dly_store_ring[20] a_26247_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X343 a_24477_6031# tdc1.r_dly_store_ctr[1] a_24131_6281# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X344 a_25348_10633# _105_ a_25616_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X346 VPWR tdc1.r_dly_store_ring[25] a_30101_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X347 a_11517_12809# _123_ a_11435_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X349 a_18243_8751# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X350 net25 a_15719_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X351 VGND a_9924_14165# net29 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X352 a_29997_8207# a_29007_8207# a_29871_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X353 a_5043_8372# tdc1.w_ring_norsz[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X354 tdc1.w_ring_buf[4] a_20083_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
R8 VGND uio_out[0] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X356 a_22273_10927# tdc0.w_ring_norsz[20] a_22189_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X357 VGND a_5951_7485# a_6119_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X358 a_25847_8751# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X359 a_4295_10749# a_3597_10383# a_4038_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X361 tdc0.w_ring_buf[30] a_8583_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X363 _136_ a_10147_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X364 VGND a_15399_4399# _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X366 a_10781_10633# tdc0.r_dly_store_ring[16] a_10699_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X367 VGND _065_ a_19163_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X368 VPWR a_21923_4399# _166_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X369 a_24276_9269# net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X370 a_24481_7669# a_24315_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X371 VGND a_17100_14165# net32 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X372 a_10291_4373# _166_ a_10689_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X375 a_26329_6281# tdc1.r_dly_store_ctr[4] a_26247_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X376 VGND tdc0.w_ring_norsz[28] a_18151_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X377 a_5629_12809# net59 tdc0.w_ring_int_norsz[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X378 a_9551_15511# tdc0.r_ring_ctr[6] a_9785_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X379 _036_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X380 a_14155_4917# tdc1.r_ring_ctr[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X381 tdc1.w_ring_buf[29] a_15023_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X382 a_23009_6575# tdc1.w_ring_norsz[20] a_22925_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X384 a_5871_11146# tdc0.w_ring_norsz[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X385 a_21449_4765# tdc1.r_ring_ctr[1] a_21361_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X386 a_13551_7119# _076_ a_13729_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X387 a_24765_9839# _090_ a_24849_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X388 a_14351_10633# _191_ a_14279_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X389 net30 a_11763_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X390 VGND net33 a_21279_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X391 VPWR a_17095_13799# tdc0.r_dly_store_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X393 a_8569_14191# tdc0.r_ring_ctr[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X394 a_10405_14013# a_9871_13647# a_10310_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X395 a_9740_3855# a_9514_3901# a_9371_4007# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X396 VPWR a_17413_3009# a_17303_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X397 VGND net40 tdc1.w_ring_int_norsz[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X399 a_21633_9839# tdc0.w_ring_buf[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X400 a_16385_9845# a_16219_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X401 a_25041_7369# _099_ a_24959_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X402 a_3859_12559# a_3413_12559# a_3763_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X403 VGND ui_in[1] a_855_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X404 a_10478_13759# a_10310_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X405 VGND a_6503_10749# a_6671_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X406 tdc1.r_dly_store_ring[8] a_13019_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X407 a_18751_8359# _084_ a_19220_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X408 VGND net32 a_19623_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X409 a_7369_6397# a_6835_6031# a_7274_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X410 VPWR _166_ a_10607_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X412 a_7009_7369# net38 tdc1.w_ring_int_norsz[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X413 _048_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X414 tdc0.w_ring_buf[8] a_11435_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X415 a_2490_11059# a_2807_11169# a_2765_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X416 a_7539_4777# a_7093_4405# a_7443_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X417 _106_ a_26247_6281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X418 _078_ a_24131_6281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X419 VPWR a_29871_7485# a_30039_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X420 a_12875_14709# _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X421 tdc0.w_ring_norsz[11] net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X422 tdc1.r_dly_store_ring[14] a_19459_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X423 VPWR a_15543_7895# _118_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X424 VPWR a_15871_7387# a_15787_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X427 _057_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X428 VPWR a_9204_3689# a_9379_3615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X429 a_15738_6397# a_15299_6031# a_15653_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X430 a_15391_10633# _114_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X431 VGND tdc0.w_ring_norsz[11] a_21739_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X432 VPWR a_22811_3615# tdc1.r_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X433 VGND tdc0.w_ring_norsz[20] a_22843_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X435 a_5015_9295# a_4761_9622# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X436 VGND net24 tdc0.w_ring_norsz[19] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X437 tdc0.w_ring_buf[11] a_21739_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X439 a_5257_11471# tdc0.w_ring_buf[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X440 VGND tdc1.r_ring_ctr[15] a_2519_7369# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X441 a_22695_5487# a_21997_5493# a_22438_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X444 a_23033_7663# tdc1.w_ring_norsz[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X445 a_16003_4917# a_15828_4943# a_16182_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X446 a_6813_8457# net60 a_6559_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X447 uo_out[1] a_24849_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X448 a_3855_4943# a_3339_4943# a_3760_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X449 _066_ _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X450 VGND a_27066_11204# a_26995_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X452 a_21545_10633# _072_ a_21399_10535# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X453 a_9493_9839# _071_ a_9577_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X454 VPWR tdc0.w_ring_norsz[12] a_19245_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X456 VGND _173_ a_10761_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X458 a_15278_7485# a_14839_7119# a_15193_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X459 tdc0.w_ring_norsz[16] tdc0.w_ring_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X460 a_18029_13647# a_17482_13921# a_17682_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X462 VGND _175_ a_15657_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X464 VPWR a_20083_8751# _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X466 a_20613_13423# tdc0.r_dly_store_ctr[1] a_20175_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X469 VGND a_19567_5309# a_19735_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X470 VPWR a_22657_4097# a_22547_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X471 VGND a_10569_7093# _131_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X472 a_17100_14165# net33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X473 a_21445_9845# a_21279_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X474 VPWR a_10478_13759# a_10405_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X475 VPWR a_8695_7637# a_8611_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X478 a_20062_12925# a_19789_12559# a_19977_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X479 a_28441_7663# tdc1.w_ring_buf[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X480 tdc0.r_dly_store_ring[5] a_17251_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X482 a_27705_5487# tdc1.w_ring_buf[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X484 VGND a_16771_7663# _070_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X485 tdc1.r_ring_ctr[1] a_22811_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X486 a_10662_5055# a_10494_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X487 VGND tdc1.r_ring_ctr[3] _167_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 VGND tdc1.r_ring_ctr[0] _016_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X489 VGND net16 tdc1.w_ring_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X490 a_20065_9661# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X491 _050_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X492 a_12353_14977# a_12135_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X493 a_23021_8751# tdc1.w_ring_norsz[1] a_22937_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 VPWR a_21891_15797# a_21878_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X495 VPWR a_9466_8319# a_9393_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X496 a_18869_10383# a_18703_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X499 VPWR a_12667_5309# a_12835_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X500 tdc0.w_ring_norsz[7] tdc0.w_ring_norsz[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X501 VGND _086_ a_13814_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X502 VPWR tdc0.r_ring_ctr[0] _000_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X503 a_21633_8751# tdc1.w_ring_buf[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X504 a_7539_14495# _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X505 a_16163_6397# a_15299_6031# a_15906_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X506 VPWR tdc1.r_ring_ctr[0] a_20635_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X509 net6 a_15575_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X510 a_8493_10927# tdc0.w_ring_int_norsz[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X511 a_9976_11305# a_9577_10933# a_9850_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X512 VGND tdc1.w_ring_norsz[6] tdc1.w_ring_norsz[22] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X513 a_8546_11989# a_8378_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X514 a_8544_3677# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X515 VGND _064_ a_19605_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X516 tdc1.w_ring_norsz[8] net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X517 VPWR a_24519_4373# a_24435_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X518 tdc1.r_ring_ctr[14] a_4595_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X519 tdc1.w_ring_buf[26] a_27443_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X520 tdc0.r_dly_store_ring[21] a_14767_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X522 a_11245_11471# tdc0.r_dly_store_ring[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X523 tdc1.r_ring_ctr[0] a_20327_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X524 a_15864_6031# a_15465_6031# a_15738_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X525 VPWR a_12743_10651# a_12659_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X526 a_25221_13103# tdc0.w_ring_buf[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X527 tdc1.r_ring_ctr[7] a_7723_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X529 a_11299_6794# tdc1.w_ring_norsz[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X531 tdc1.w_ring_buf[30] a_8491_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X533 a_6983_3855# a_6633_3855# a_6888_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X534 VPWR _080_ a_21637_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X535 tdc0.r_dly_store_ctr[8] a_14583_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R9 VPWR tdc1.g_ring3[21].stg01_66.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X536 a_7001_6031# a_6835_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X538 VGND a_27038_11989# a_26996_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X539 _015_ a_15687_15823# a_15925_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X542 a_30254_7895# a_30350_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X545 VGND a_13243_5705# a_13250_5609# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X546 a_16217_3311# _166_ a_16135_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X547 VPWR ui_in[4] a_16219_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X548 a_10594_9295# _139_ a_10124_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X550 a_18501_7663# a_18335_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X553 a_14610_3311# a_13533_3317# a_14448_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X554 a_22511_14013# a_21647_13647# a_22254_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X556 tdc0.r_ring_ctr[1] a_21891_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X557 a_20717_4765# tdc1.r_ring_ctr[0] a_20635_4512# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X558 VPWR _067_ a_25125_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X561 a_22535_3855# a_22089_3855# a_22439_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X563 a_15404_7119# a_15005_7119# a_15278_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X564 a_20617_6575# tdc1.r_dly_store_ring[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X565 a_18087_8573# a_17305_8207# a_18003_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X567 a_4503_7093# _063_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X568 a_28047_12247# a_28331_12233# a_28266_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X569 a_23473_9839# tdc1.w_ring_buf[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X570 tdc0.r_ring_ctr[14] a_4503_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X571 a_27517_5493# a_27351_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X572 tdc1.r_dly_store_ctr[6] a_11087_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X574 _065_ a_16771_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X575 a_22181_14013# a_21647_13647# a_22086_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X576 VPWR tdc1.w_ring_norsz[3] a_23661_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X577 VPWR _064_ a_19066_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X578 a_27479_9839# a_26781_9845# a_27222_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X579 VGND net26 a_4259_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X580 a_27054_9839# a_26615_9845# a_26969_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X581 a_3337_11721# _161_ a_3255_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X583 VGND tdc0.w_ring_norsz[30] a_8583_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X584 a_9393_8573# a_8859_8207# a_9298_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X585 a_22254_13759# a_22086_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X586 VPWR net31 a_18427_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X587 a_8527_7663# a_7829_7669# a_8270_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X588 VPWR a_22771_13077# a_22687_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X589 a_7055_12925# a_6191_12559# a_6798_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X590 a_8686_15395# _152_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X591 VGND tdc0.r_ring_ctr[8] a_12823_16073# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X592 a_24669_7663# tdc1.w_ring_buf[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X593 VGND tdc0.w_ring_norsz[18] tdc0.w_ring_int_norsz[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X594 a_10401_12393# a_9411_12021# a_10275_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X595 VGND a_10443_10901# a_10401_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X596 a_7167_15657# a_6817_15285# a_7072_15645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X598 a_6035_7485# a_5253_7119# a_5951_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X599 VPWR a_3399_12275# net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X600 VGND a_20223_13799# tdc0.r_dly_store_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X601 VPWR _150_ a_10239_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
R10 uio_out[4] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X603 VGND a_9103_4659# net15 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X604 a_5161_13647# a_4995_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X605 VGND a_15256_10535# _117_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X607 _001_ a_16595_14985# a_16845_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X609 VPWR _161_ a_3505_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X610 a_16104_13647# a_15023_13647# a_15757_13889# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X611 _108_ a_20451_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X612 a_8451_15797# a_8654_16075# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X613 a_17865_6575# net19 tdc1.w_ring_norsz[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X614 a_22565_15253# a_22347_15657# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X615 a_29361_7119# tdc1.w_ring_buf[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X616 a_24922_7637# a_24754_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X618 a_19310_13759# a_19142_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X619 a_26334_11721# _092_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X620 a_10797_8457# tdc1.w_ring_norsz[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X621 VPWR a_24719_12015# a_24887_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X622 VPWR net37 a_13551_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X623 a_19959_15797# a_19784_15823# a_20138_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X624 a_24294_15101# a_24021_14735# a_24209_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X626 a_25129_5487# tdc1.w_ring_buf[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X627 VGND a_15906_6143# a_15864_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X628 VGND _062_ a_4117_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X629 _049_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X630 VPWR net30 a_14839_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X631 VGND a_24719_12015# a_24887_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X632 VGND net21 tdc0.w_ring_norsz[23] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X633 VGND a_8399_3855# _196_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X634 VGND tdc0.w_ring_norsz[19] tdc0.w_ring_int_norsz[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X635 _190_ a_13814_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X636 a_8887_12015# a_8105_12021# a_8803_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X638 a_3981_12801# a_3763_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X639 VGND a_3399_12275# net20 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X641 a_14059_8983# a_14332_8983# a_14290_9111# VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X643 VPWR a_24719_15101# a_24887_15003# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X645 VGND net29 a_9411_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X648 VGND net10 a_16311_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X649 VPWR _143_ a_9551_15511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X650 _018_ a_14644_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.327 ps=1.65 w=1 l=0.15
X652 VPWR a_22254_13759# a_22181_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X653 VGND a_15446_7231# a_15404_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X654 _043_ net23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X655 tdc1.w_ring_norsz[11] net17 a_27529_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X656 VGND net29 a_14103_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X658 VPWR a_3981_12801# a_3871_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X660 a_5449_4719# _180_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X661 a_9631_6397# a_8767_6031# a_9374_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X662 tdc1.w_ring_norsz[25] tdc1.w_ring_int_norsz[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X663 VGND a_29062_8725# a_29020_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X664 VPWR net27 a_4903_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X665 a_9897_4737# tdc1.r_ring_ctr[6] a_9811_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X666 a_19651_10749# a_18869_10383# a_19567_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 VGND net8 a_16679_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X670 VGND a_21115_6299# a_21073_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X671 a_19439_9111# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X672 uo_out[2] a_26420_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X673 a_14008_9545# _189_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X674 a_15919_14735# tdc0.r_ring_ctr[10] a_15823_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X675 a_7539_14495# a_7364_14569# a_7718_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X676 VGND _069_ a_27329_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X677 a_20525_4943# a_20359_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X679 a_26781_9845# a_26615_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X680 VPWR tdc1.w_ring_norsz[27] a_26145_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X681 a_21361_7369# _094_ a_21279_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X682 a_21056_15823# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
R11 tt_um_hpretl_tt06_tdc_v2_79.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X683 VPWR a_17740_10071# _122_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X686 a_19849_3677# a_19805_3285# a_19683_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X687 a_11950_14165# a_11782_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X688 tdc0.w_ring_buf[12] a_19899_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X689 VPWR net34 a_23303_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X690 VGND tdc1.r_dly_store_ring[11] a_30021_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X691 a_8929_15823# a_8451_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X692 VPWR a_16104_13647# a_16279_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X693 tdc0.w_ring_buf[28] a_18151_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X695 VPWR tdc0.w_ring_int_norsz[8] a_8197_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X696 a_7061_14557# a_7017_14165# a_6895_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X698 a_10124_9269# _134_ a_10946_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X699 a_26420_11721# _093_ a_26334_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X700 a_19329_9839# a_19163_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X702 VGND a_24462_11989# a_24420_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X703 VPWR _173_ a_10291_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X704 VGND tdc1.w_ring_norsz[0] a_5547_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X705 VGND net7 a_21555_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X707 VGND a_29871_7485# a_30039_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X711 a_9117_5309# a_8583_4943# a_9022_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X712 a_15481_4399# _177_ a_15399_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X713 a_9836_4105# _171_ a_9371_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X714 VPWR a_16331_6299# a_16247_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X715 tdc1.r_dly_store_ring[10] a_27647_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X716 net38 a_16463_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X718 a_6105_5807# tdc1.r_ring_ctr[13] a_6002_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X719 tdc0.r_ring_ctr[13] a_7539_14495# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X720 VGND a_7223_9813# a_7181_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X721 a_26065_6575# tdc1.w_ring_int_norsz[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X722 a_25815_14191# a_25033_14197# a_25731_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X723 VGND net17 tdc1.w_ring_norsz[20] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X725 a_11655_6397# a_10791_6031# a_11398_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X727 VGND tdc1.w_ring_norsz[27] tdc1.w_ring_norsz[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X729 net33 a_17283_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X730 a_12291_14191# a_11509_14197# a_12207_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X731 VPWR tdc0.r_dly_store_ring[1] a_21270_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X733 VPWR net27 a_4995_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X734 a_23937_8457# net17 tdc1.w_ring_norsz[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X735 VPWR tdc0.r_ring_ctr[14] a_4219_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X736 tdc1.w_ring_int_norsz[19] net64 a_24137_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X737 _124_ a_11435_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X739 a_25616_10633# _104_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X741 VPWR tdc1.r_dly_store_ring[27] a_29733_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X742 a_16155_7895# tdc1.r_dly_store_ring[29] a_16301_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X743 a_14158_13077# a_13990_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X745 a_14644_5487# _180_ a_14471_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X746 a_10787_7369# _084_ a_10569_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X749 VGND a_21912_6575# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X750 a_22189_10927# net22 tdc0.w_ring_norsz[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X751 a_17831_13647# a_17611_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X752 VGND net8 a_21923_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X753 a_22269_10217# a_21279_9845# a_22143_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X754 a_22179_3311# a_21555_3317# a_22071_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X755 VPWR tdc0.r_ring_ctr[1] a_21157_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X758 VPWR a_19034_6549# a_18961_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X759 a_24205_10933# a_24039_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X760 a_20617_6397# a_20083_6031# a_20522_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X761 a_6633_3855# a_6467_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X762 _115_ a_15207_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X764 VGND tdc0.w_ring_norsz[18] tdc0.w_ring_norsz[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X765 a_20817_3017# tdc1.r_ring_ctr[1] a_20735_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X766 VGND a_22339_10535# tdc0.r_dly_store_ring[20] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X767 a_21707_7881# net33 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X769 a_2769_7369# tdc1.r_ring_ctr[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X770 a_25765_12335# tdc0.r_dly_store_ring[2] a_25327_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X771 a_19977_12559# tdc0.w_ring_buf[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X774 VPWR a_16771_7663# _070_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X775 a_21912_6575# _113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X776 a_30856_7895# ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X777 VGND net17 tdc1.w_ring_norsz[19] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X778 a_18243_8751# _065_ a_18243_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X779 VPWR net8 a_16679_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X780 a_9953_7119# tdc1.r_dly_store_ctr[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X781 _130_ a_11713_6691# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X782 a_23358_3855# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X783 VGND a_22771_13077# a_22729_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X784 VGND a_4219_13621# _161_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X785 a_5234_14735# _044_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X786 a_17433_14013# a_17095_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X787 a_25221_3855# tdc1.r_ring_ctr[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X788 a_29035_9447# tdc1.r_dly_store_ring[26] a_29181_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X792 VPWR a_17739_8970# tdc1.w_ring_buf[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X793 VGND _129_ a_11713_6691# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R12 net50 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X794 VPWR a_4503_7093# a_4490_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X795 VPWR a_9799_6299# a_9715_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X796 VPWR _195_ _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X797 VPWR a_14899_15797# tdc0.r_ring_ctr[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X799 a_15701_8457# _065_ a_15283_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X800 a_12594_7637# a_12426_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X803 a_22269_9129# a_21279_8757# a_22143_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X804 a_7348_4765# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X805 a_7829_7669# a_7663_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X806 a_8285_9129# a_7295_8757# a_8159_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X807 VPWR _006_ a_3526_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X809 VPWR net1 a_26983_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X810 VGND tdc0.w_ring_norsz[27] tdc0.w_ring_norsz[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X811 a_15333_9545# _117_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X812 a_13882_6549# a_13714_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X813 a_14351_4943# tdc1.r_ring_ctr[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X814 VGND tdc1.w_ring_int_norsz[13] tdc1.w_ring_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X815 _134_ a_10241_7779# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X816 a_8753_7119# tdc1.w_ring_buf[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X817 a_25029_6953# a_24039_6581# a_24903_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X820 VPWR _066_ a_21445_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X821 _087_ a_19329_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X822 VGND _006_ a_3526_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X823 _014_ _152_ a_13073_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X824 a_15653_6031# tdc1.w_ring_buf[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X827 a_27054_9839# a_26781_9845# a_26969_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X828 a_14553_4943# tdc1.r_ring_ctr[9] a_14447_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X830 tdc0.w_ring_buf[23] a_7755_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X831 net22 a_19255_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X832 _133_ a_9595_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X833 VPWR net8 a_21923_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X834 VGND a_25071_6549# a_25029_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X836 a_21886_9813# a_21718_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X837 a_27958_5461# a_27790_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X838 a_21914_7940# a_21707_7881# a_22090_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X839 VGND a_13735_12559# net23 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X840 a_11839_13103# a_10975_13109# a_11582_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X841 a_18149_14165# a_17931_14569# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X842 a_6633_3855# a_6467_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X843 a_22289_3285# a_22071_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X844 VPWR a_14800_6549# net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X845 _061_ net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X846 net12 a_19255_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X847 a_11621_8457# tdc1.w_ring_int_norsz[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X848 a_16845_9295# a_16679_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X849 VPWR net36 a_26615_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X850 a_15193_7119# tdc1.w_ring_buf[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X851 VGND a_8527_7663# a_8695_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X852 a_28441_9839# tdc1.w_ring_buf[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X854 VPWR _107_ a_21998_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X855 a_9029_13103# tdc0.w_ring_buf[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X857 VGND _151_ a_10699_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X860 a_22252_15645# _009_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X861 VPWR a_8822_14165# a_8749_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X862 a_15649_4719# tdc1.r_ring_ctr[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X863 _175_ a_11067_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X864 VGND tdc1.w_ring_norsz[19] a_23855_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X865 a_16826_9813# a_16658_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X867 a_4237_8207# a_3247_8207# a_4111_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X868 tdc0.w_ring_norsz[18] tdc0.w_ring_int_norsz[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X869 a_13989_7119# tdc1.r_dly_store_ctr[5] a_13551_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X870 tdc1.w_ring_norsz[16] net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X871 _059_ net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X872 VPWR a_7897_7284# net13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X874 a_12793_13423# tdc0.r_dly_store_ctr[4] a_12447_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X875 a_22270_5487# a_21831_5493# a_22185_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X876 a_6273_14985# _157_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X878 a_24674_9295# _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X879 a_3413_9295# a_3247_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X880 VPWR a_22143_9839# a_22311_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X881 VGND net30 a_14839_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X883 a_21878_16189# a_20801_15823# a_21716_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X885 a_20241_9295# _064_ a_20169_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X886 _083_ a_20083_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X887 a_11414_13103# a_11141_13109# a_11329_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X888 a_13887_8359# net25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X889 a_11059_9955# _137_ a_10977_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X890 VGND net20 tdc0.w_ring_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X891 VGND net75 tdc1.w_ring_int_norsz[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X892 VPWR a_10124_9269# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X893 VPWR net30 a_15299_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X894 tdc0.r_dly_store_ring[21] a_14767_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X895 a_20314_3311# a_19237_3317# a_20152_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X896 a_15333_9545# _122_ a_15504_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X897 VPWR a_11823_6299# a_11739_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X898 VGND tdc1.w_ring_norsz[31] a_7295_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X899 a_17303_4399# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X901 a_21886_8725# a_21718_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X902 tdc0.w_ring_buf[19] a_23303_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X903 tdc0.r_ring_ctr[3] a_23087_15583# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X904 VPWR tdc0.w_ring_int_norsz[29] a_13809_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X905 a_11398_6143# a_11230_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X906 VPWR a_6503_10749# a_6671_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X908 VPWR tdc1.r_ring_ctr[7] a_9811_4737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X909 VGND net37 a_2511_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X910 a_17493_12559# tdc0.w_ring_buf[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X911 a_17581_14197# a_17415_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X913 VPWR a_5510_11583# a_5437_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X914 a_22090_7663# a_21843_8041# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X915 a_10436_13647# a_10037_13647# a_10310_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X917 a_24305_8457# net63 tdc1.w_ring_int_norsz[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X918 VPWR a_25163_8725# a_25079_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X919 a_8008_4777# a_6927_4405# a_7661_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X920 tdc0.r_dly_store_ctr[15] a_4463_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X921 a_11978_3631# _166_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X922 tdc0.w_ring_norsz[25] net23 a_17869_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X923 a_2932_14165# net28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X924 a_20046_5461# a_19878_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X925 a_12959_5719# a_13250_5609# a_13201_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X926 a_26995_11305# a_26866_11049# a_26575_11159# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X928 tdc1.w_ring_norsz[27] net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X929 a_14265_14569# a_13275_14197# a_14139_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X930 a_8749_4943# a_8583_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X931 a_29319_8751# a_28621_8757# a_29062_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X934 a_28253_9845# a_28087_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X935 a_19142_5309# a_18869_4943# a_19057_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X937 a_18781_6575# tdc1.w_ring_buf[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X938 a_7348_4765# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X941 a_9677_7663# tdc1.r_dly_store_ring[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X942 a_16468_9111# net4 a_16396_9111# VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X943 a_23021_12015# tdc0.w_ring_norsz[2] a_22937_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 a_24922_7637# a_24754_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X945 VGND _196_ _048_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X946 a_9577_9839# tdc0.r_dly_store_ctr[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X947 a_17305_8207# a_17139_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X948 tdc0.w_ring_int_norsz[6] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X951 a_12897_6575# net16 tdc1.w_ring_norsz[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X952 VPWR _083_ a_25609_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X954 a_17935_4703# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X955 VGND _068_ a_10173_10411# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X956 tdc1.w_ring_int_norsz[10] tdc1.w_ring_norsz[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X957 a_12613_12809# tdc0.w_ring_norsz[14] a_12529_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X959 a_11981_11721# tdc0.w_ring_norsz[22] a_11897_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X960 VPWR _118_ a_15179_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X961 VGND a_4503_7093# a_4437_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X962 a_11697_14191# tdc0.r_ring_ctr[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X963 a_9389_7119# a_8399_7119# a_9263_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X964 a_24765_9839# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X966 a_22903_14709# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X967 _021_ _184_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X969 a_15635_13647# a_15189_13647# a_15539_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X971 VGND a_14059_8983# _076_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X972 a_24903_10927# a_24205_10933# a_24646_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X973 tdc1.w_ring_buf[29] a_15023_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X974 a_12667_5309# a_11969_4943# a_12410_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X975 VPWR net3 _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X976 a_5635_5193# _181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X977 VGND tdc1.w_ring_norsz[3] a_24223_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X978 tdc0.r_ring_ctr[12] a_5055_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X980 tdc0.w_ring_norsz[17] net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X981 VPWR a_28215_5487# a_28383_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X984 a_11973_9295# tdc1.w_ring_buf[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X985 VPWR tdc0.w_ring_int_norsz[28] a_19697_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X986 VPWR a_3399_12275# net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X988 net16 a_14800_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X989 a_19032_4765# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X990 a_22396_5865# a_21997_5493# a_22270_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X992 a_26859_11145# net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X993 tdc0.w_ring_int_norsz[19] net46 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X994 VPWR tdc0.r_ring_ctr[8] _153_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X995 VGND net20 tdc0.w_ring_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X996 VGND _045_ a_7061_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X997 a_5253_7119# a_5087_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X998 VGND a_22311_9813# a_22269_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1000 VGND net27 a_4995_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1001 tdc1.w_ring_buf[12] a_27167_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1003 a_20801_15823# a_20635_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1005 tdc1.w_ring_norsz[26] tdc1.w_ring_norsz[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1006 VPWR a_22143_8751# a_22311_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1007 VPWR tdc1.w_ring_norsz[17] a_23855_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1008 a_14967_12015# a_14269_12021# a_14710_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1010 VPWR net22 _042_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1012 tdc1.w_ring_norsz[0] net16 a_6997_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1013 VGND _058_ a_17457_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1014 a_14833_15823# a_13643_15823# a_14724_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1015 VGND a_20506_11583# a_20464_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1016 VPWR a_20655_12827# a_20571_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1018 a_15189_13647# a_15023_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1019 a_10494_5309# a_10055_4943# a_10409_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1020 a_12863_5719# a_12959_5719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1021 a_24719_12015# a_24021_12021# a_24462_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1022 a_7017_14165# a_6799_14569# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1023 VPWR a_14583_13915# a_14499_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1024 a_21997_5493# a_21831_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1025 VPWR _070_ a_19991_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1027 VPWR a_8183_4703# tdc1.r_ring_ctr[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1028 VGND a_3399_12275# net20 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1029 VGND tdc1.w_ring_int_norsz[29] tdc1.w_ring_norsz[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1030 tdc0.w_ring_int_norsz[20] net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1032 VPWR a_27222_9813# a_27149_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1033 a_19492_3677# _016_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1034 a_9493_9839# net3 a_9411_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1035 tdc1.w_ring_norsz[2] net17 a_23389_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1036 a_20223_13799# a_20319_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1037 VGND a_20046_5461# a_20004_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1038 VPWR net19 _058_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1039 tdc1.w_ring_norsz[9] net18 a_27069_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1040 VGND tdc0.w_ring_int_norsz[14] tdc0.w_ring_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1041 VPWR net29 a_11343_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1042 a_12701_10383# a_11711_10383# a_12575_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1043 VGND a_9371_4007# _029_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1045 _074_ a_14794_9922# a_15057_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X1046 a_21743_6895# _107_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
X1048 VPWR a_12207_14191# a_12375_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1051 tdc0.w_dly_stop[3] a_2787_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1052 a_26870_12015# a_26431_12021# a_26785_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1054 a_19567_10749# a_18703_10383# a_19310_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1055 VPWR a_20327_3615# tdc1.r_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1056 a_7369_13109# a_7203_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1057 tdc1.r_dly_store_ring[8] a_13019_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1058 VGND _141_ _144_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1059 VGND a_14431_4373# _178_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1060 a_15717_8001# _071_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X1061 VPWR tdc0.r_dly_store_ring[20] a_21545_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X1063 VGND net36 a_26615_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1064 a_12851_7663# a_11987_7669# a_12594_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1065 a_19237_10749# a_18703_10383# a_19142_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1066 a_17413_4373# a_17195_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1068 VGND _068_ a_13161_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1069 a_13441_14197# a_13275_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1070 VPWR a_4420_4943# a_4595_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1071 tdc1.r_dly_store_ring[14] a_19459_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1072 VPWR a_25179_7663# a_25347_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1073 a_9585_11721# net50 tdc0.w_ring_int_norsz[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1074 a_7734_8751# a_7461_8757# a_7649_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1075 a_12897_12809# net57 tdc0.w_ring_int_norsz[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1077 VGND net10 a_21831_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1078 a_16279_13621# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1079 VGND a_19723_15279# _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X1080 a_8197_10927# tdc0.w_ring_norsz[24] a_8113_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1081 VPWR a_18149_14165# a_18039_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1082 VPWR net33 a_19899_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1083 a_17935_2741# a_17760_2767# a_18114_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1085 tdc0.r_dly_store_ctr[5] a_14307_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1086 net38 a_16463_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1087 VPWR _134_ a_10512_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1088 a_25071_9813# _085_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1090 a_14448_3689# a_13533_3317# a_14101_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1091 VPWR _081_ a_19655_8235# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1092 VPWR a_18751_8359# _129_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X1093 a_12525_4399# tdc1.r_ring_ctr[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1095 VPWR tdc1.w_ring_norsz[11] a_27065_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1097 tdc1.r_ring_ctr[0] a_20327_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1098 net6 a_15575_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1100 VPWR a_17392_15823# a_17567_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1102 VPWR net30 a_10791_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1103 tdc1.w_ring_buf[26] a_27443_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1104 a_15481_5185# a_15263_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
R13 VPWR tdc0.g_ring3[19].stg01_46.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1105 a_28687_12381# a_28467_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1106 VGND _049_ a_22333_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1107 tdc0.r_dly_store_ring[7] a_5291_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1108 a_12207_14191# a_11343_14197# a_11950_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1109 a_13882_14165# a_13714_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1110 a_10620_4943# a_10221_4943# a_10494_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1111 VGND net34 a_28087_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1116 a_20046_5461# a_19878_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1117 tdc1.w_ring_buf[30] a_8491_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1118 a_13714_6575# a_13275_6581# a_13629_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1119 a_26847_9460# tdc1.w_ring_norsz[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1120 a_10594_9295# _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X1121 a_6078_10749# a_5805_10383# a_5993_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1123 tdc1.r_ring_ctr[3] a_23179_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1124 a_28813_6575# _072_ a_28897_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1125 VPWR tdc1.w_ring_int_norsz[12] a_26781_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1126 VPWR _065_ a_19425_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X1127 VGND a_15159_8725# _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1129 a_3871_12925# a_3247_12559# a_3763_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1131 a_24803_12015# a_24021_12021# a_24719_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1132 a_22779_5487# a_21997_5493# a_22695_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1133 VGND ui_in[4] a_16219_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1134 a_11299_6794# tdc1.w_ring_norsz[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1135 VGND a_8543_15253# _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1136 VPWR a_19310_5055# a_19237_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1137 net34 a_24276_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1138 VPWR a_14899_15797# a_14886_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1139 VPWR net31 a_19439_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1140 VPWR net27 a_3431_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1141 VGND tdc0.w_ring_norsz[19] a_23303_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1142 VPWR a_9459_8970# tdc1.w_ring_buf[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1144 a_6545_9839# tdc0.w_ring_buf[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1145 a_10037_13647# a_9871_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1146 a_21031_6397# a_20249_6031# a_20947_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1147 VGND a_14899_15797# a_14833_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1149 a_13882_6549# a_13714_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1150 a_16658_9839# a_16219_9845# a_16573_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1152 VGND a_17727_5487# a_17895_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1153 VPWR a_24887_15003# a_24803_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1154 VGND a_4279_8475# a_4237_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1155 VGND a_25899_13077# a_25857_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1157 a_19310_10495# a_19142_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1158 tdc0.w_ring_norsz[2] tdc0.w_ring_int_norsz[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1160 VPWR tdc1.w_ring_norsz[21] a_17221_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1161 a_15335_8181# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1162 a_10229_9839# tdc0.r_dly_store_ctr[15] a_10147_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1163 a_16385_12015# tdc0.w_ring_norsz[17] a_16301_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1164 a_29169_6895# tdc1.r_dly_store_ring[28] a_28731_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1167 a_21151_15823# a_20635_15823# a_21056_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1168 a_4425_9845# a_4259_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1169 a_15757_13889# a_15539_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1170 VGND _066_ a_11987_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1171 VGND a_12575_10749# a_12743_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R14 VGND uio_oe[0] sky130_fd_pr__res_generic_po w=0.48 l=0.045
R15 tt_um_hpretl_tt06_tdc_v2_91.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1172 a_12437_6281# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1173 a_21914_7940# a_21714_7785# a_22063_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
R16 net72 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1175 a_17045_16065# a_16827_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1176 a_6824_13647# tdc0.r_ring_ctr[12] a_6521_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1177 VPWR a_17010_13077# a_16937_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1179 a_11623_12335# _125_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1180 a_6027_9295# a_5773_9622# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1181 a_17760_4777# a_16679_4405# a_17413_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1182 a_20739_13647# a_20610_13921# a_20319_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1183 a_11878_12015# _125_ a_11792_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1184 VGND tdc1.r_dly_store_ctr[6] a_12725_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1187 a_17195_4777# a_16679_4405# a_17100_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1188 a_9573_4943# a_8583_4943# a_9447_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1190 VGND a_14307_14165# a_14265_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1191 a_4529_6031# a_3339_6031# a_4420_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1192 a_8102_9839# a_7829_9845# a_8017_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1193 _047_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1195 VPWR tdc0.w_ring_norsz[2] a_23855_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1196 a_29446_7485# a_29173_7119# a_29361_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1197 a_13620_9269# _194_ a_14008_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1199 VGND a_20947_6397# a_21115_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1200 VPWR tdc0.w_ring_int_norsz[13] a_13441_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1201 tdc0.r_ring_ctr[8] a_14899_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X1202 a_19219_15823# a_18869_15823# a_19124_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1204 a_11599_3133# _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1205 a_25033_13109# a_24867_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1207 net15 a_9103_4659# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1208 VPWR a_18169_10137# a_18199_9878# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1209 _136_ a_10147_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1210 VGND a_5043_11146# tdc0.w_ring_buf[16] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1211 a_23650_13103# a_23211_13109# a_23565_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1212 a_6077_8457# net15 tdc1.w_ring_norsz[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1213 a_9205_14569# a_8215_14197# a_9079_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1214 a_21327_7895# a_21423_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1216 a_25723_5487# a_24941_5493# a_25639_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1217 tdc0.w_ring_norsz[9] net23 a_17501_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1218 a_6364_14985# _160_ a_6191_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1219 VGND a_27411_7093# net19 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1220 a_23473_9839# tdc1.w_ring_buf[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1221 a_15828_4943# a_14913_4943# a_15481_5185# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1223 a_25815_4221# a_25033_3855# a_25731_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1224 a_13553_8867# _187_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1225 a_24393_6575# tdc1.w_ring_buf[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1226 _067_ a_11987_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1227 a_6177_6575# tdc1.r_ring_ctr[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1228 a_10946_9295# _138_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X1229 a_6357_9845# a_6191_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1231 a_13840_6953# a_13441_6581# a_13714_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1232 VGND a_3115_9813# net26 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1233 tdc1.r_dly_store_ring[7] a_5291_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1234 a_17029_5493# a_16863_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1236 a_16589_7983# _066_ a_16155_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1238 a_17305_8207# a_17139_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1239 tdc0.w_dly_stop[3] a_2787_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1240 VGND a_21399_10535# _109_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1243 a_25973_9301# _096_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1244 a_17286_9407# a_17118_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1245 a_9366_3311# a_8289_3317# a_9204_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1246 a_13265_6281# net39 tdc1.w_ring_int_norsz[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1247 VGND a_9431_7387# a_9389_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1249 VGND net15 _063_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1250 a_17286_9407# a_17118_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1252 a_20261_3689# a_19071_3317# a_20152_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1253 VGND net53 tdc0.w_ring_int_norsz[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1254 a_26053_6281# net74 tdc1.w_ring_int_norsz[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1259 VGND a_11067_4399# _175_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R17 VGND net44 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1260 VPWR a_27958_5461# a_27885_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1261 VGND tdc1.w_ring_int_norsz[21] tdc1.w_ring_norsz[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1262 a_22351_9545# _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1263 a_5257_11471# tdc0.w_ring_buf[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1264 VGND _066_ a_9941_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1265 a_24297_8757# a_24131_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1266 _037_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1267 a_12483_9661# a_11785_9295# a_12226_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1268 a_5253_7119# a_5087_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1269 VGND a_15135_11989# a_15093_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1270 VGND a_7723_3829# a_7657_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1271 a_22677_10749# a_22339_10535# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1272 a_22261_8041# a_21707_7881# a_21914_7940# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1273 a_22653_10927# tdc0.w_ring_norsz[4] a_22569_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1274 VPWR _196_ _057_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1275 a_13814_11471# tdc0.r_dly_store_ctr[8] a_13728_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1276 a_18677_8029# _064_ a_18605_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
R18 tt_um_hpretl_tt06_tdc_v2_80.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1279 tdc0.w_ring_int_norsz[12] net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1280 _081_ _065_ a_18690_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X1281 VGND tdc0.w_ring_norsz[13] tdc0.w_ring_int_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1283 a_29587_7895# tdc1.r_dly_store_ring[27] a_29733_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X1284 VPWR a_24094_4373# a_24021_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1285 a_8289_3317# a_8123_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1287 VPWR a_7902_8725# a_7829_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1288 a_29469_9295# _072_ a_29035_9447# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1289 VGND tdc1.w_ring_int_norsz[0] tdc1.w_ring_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1290 VPWR a_14583_13077# a_14499_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1291 tdc1.w_ring_int_norsz[25] net70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1293 a_7245_3855# a_7201_4097# a_7079_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1294 a_6733_7369# net77 tdc1.w_ring_int_norsz[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1295 a_16669_12015# net38 tdc0.w_ring_int_norsz[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1296 VPWR a_14139_6575# a_14307_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1297 a_14139_6575# a_13441_6581# a_13882_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1298 a_13717_7369# tdc1.r_dly_store_ctr[13] a_13633_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1299 a_22071_3689# a_21555_3317# a_21976_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1303 a_23285_9845# a_23119_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1304 a_22339_10535# a_22435_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1305 VPWR _156_ _157_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1306 VPWR net34 a_24775_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1307 VGND a_11987_9839# _067_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1309 a_24205_6581# a_24039_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1310 a_9723_8573# a_9025_8207# a_9466_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1312 a_15189_13647# a_15023_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1313 tdc1.r_ring_ctr[15] a_4503_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1314 tdc1.w_ring_int_norsz[5] net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1315 a_7829_8751# a_7295_8757# a_7734_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1316 VGND a_14623_3615# tdc1.r_ring_ctr[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1317 a_8841_13109# a_8675_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1318 _105_ a_25511_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1319 VGND tdc1.r_ring_ctr[0] a_20735_3017# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1320 a_24754_7663# a_24315_7669# a_24669_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1321 a_28526_7663# a_28253_7669# a_28441_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1323 tdc1.w_ring_norsz[23] tdc1.w_ring_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1324 a_20065_9661# a_19899_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X1325 VPWR tdc0.w_ring_int_norsz[27] a_21813_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1326 a_12056_2767# a_11141_2767# a_11709_3009# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1327 a_5069_11471# a_4903_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1328 VPWR tdc1.w_ring_norsz[14] a_8573_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1329 a_30537_7895# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1330 VPWR net27 a_7939_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1331 a_4111_8573# a_3247_8207# a_3854_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1332 _156_ a_16127_14557# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1333 a_3951_6031# a_3505_6031# a_3855_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1334 a_9190_5055# a_9022_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1335 VPWR a_27295_12015# a_27463_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1336 a_13809_12015# tdc0.w_ring_norsz[13] a_13725_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1337 a_8067_13103# a_7369_13109# a_7810_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1338 a_14064_15823# _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1339 a_6503_10749# a_5805_10383# a_6246_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1340 a_4328_12559# a_3413_12559# a_3981_12801# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1341 _159_ tdc0.r_ring_ctr[12] a_6093_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1342 VGND a_27295_12015# a_27463_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1343 a_19973_15279# tdc0.r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1344 VGND net10 a_17415_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1345 _023_ tdc1.r_ring_ctr[1] a_20985_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X1346 a_11895_3311# tdc1.r_ring_ctr[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X1347 tdc1.w_ring_norsz[16] tdc1.w_ring_int_norsz[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X1349 a_17229_4097# a_17011_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1352 a_23910_5461# a_23742_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1353 a_17869_11721# tdc0.w_ring_norsz[9] a_17785_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1354 a_24002_14165# a_23834_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1356 tdc1.r_dly_store_ctr[14] a_7867_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1357 tdc0.w_ring_buf[17] a_15483_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1358 VGND a_17739_8970# tdc1.w_ring_buf[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1359 a_27885_5487# a_27351_5493# a_27790_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1360 VPWR a_21914_7940# a_21843_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1362 a_25474_14165# a_25306_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1363 a_5015_9622# tdc0.r_dly_store_ring[0] a_5015_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1364 uo_out[4] a_21912_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1365 VPWR net27 a_4259_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1366 VGND a_14703_12724# tdc0.w_ring_buf[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1367 a_13990_14013# a_13717_13647# a_13905_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1369 a_9365_15823# _038_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X1370 a_22855_10383# a_22726_10657# a_22435_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1371 a_4315_14735# a_3965_14735# a_4220_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1372 a_8381_14197# a_8215_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1373 VPWR a_25731_4221# a_25899_4123# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1374 a_7825_6031# a_6835_6031# a_7699_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1375 VGND _195_ _039_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1376 VGND a_28331_12233# a_28338_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1377 a_19693_13647# a_18703_13647# a_19567_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1378 a_23259_7882# tdc1.w_ring_norsz[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1379 tdc0.r_dly_store_ctr[7] a_9247_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1380 _098_ a_25973_9301# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1381 a_12529_12809# net21 tdc0.w_ring_norsz[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1383 a_11897_11721# tdc0.w_ring_int_norsz[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1385 a_20503_15253# _142_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X1386 a_24393_10927# tdc0.w_ring_buf[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1387 a_21223_5309# a_20359_4943# a_20966_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1389 VPWR a_14415_14013# a_14583_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1390 a_18877_13423# tdc0.r_dly_store_ring[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1392 a_12243_15101# _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1393 VGND net2 a_3247_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1394 VPWR _181_ a_6541_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1395 VGND a_14342_10901# a_14300_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
R19 net67 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1396 VGND a_10903_13915# a_10861_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1397 _075_ a_14011_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1398 VGND tdc1.w_ring_norsz[10] tdc1.w_ring_int_norsz[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1399 VPWR a_8270_9813# a_8197_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1400 a_27295_12015# a_26431_12021# a_27038_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1401 VGND _146_ _149_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1402 a_29077_8041# a_28087_7669# a_28951_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1403 a_25264_10633# _084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X1404 a_19697_11721# tdc0.w_ring_norsz[12] a_19613_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1405 VGND a_6798_12671# a_6756_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1406 tdc1.w_ring_int_norsz[24] tdc1.w_ring_norsz[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1407 a_9643_12724# tdc0.w_ring_norsz[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1408 VPWR a_14101_3285# a_13991_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1409 a_29955_8573# a_29173_8207# a_29871_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1410 VPWR tdc0.w_ring_norsz[22] a_9585_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1411 a_9514_3901# _175_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X1412 VPWR tdc0.w_ring_norsz[29] a_12897_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1413 VGND a_24002_14165# a_23960_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
R20 VPWR tdc0.stg01_59.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1414 _089_ a_18795_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1415 a_12157_4943# tdc1.r_ring_ctr[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1416 VPWR a_29614_7231# a_29541_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1417 a_22179_3311# _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1419 _166_ a_21923_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X1420 a_18869_4943# a_18703_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1421 a_10229_13423# tdc0.r_dly_store_ctr[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1422 VGND a_18703_14735# _195_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1423 a_12410_2767# _053_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1424 a_3399_12275# net21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1425 VPWR net10 a_20635_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1426 a_20303_5487# a_19439_5493# a_20046_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1428 a_8838_7485# a_8565_7119# a_8753_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1429 a_24880_8041# a_24481_7669# a_24754_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1431 VGND a_13620_9269# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1432 a_18249_11721# tdc0.w_ring_norsz[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1433 VGND net19 tdc1.w_ring_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1435 VPWR a_8857_3285# a_8747_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1436 VGND net41 tdc1.w_ring_int_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1437 a_8017_9839# tdc0.w_ring_buf[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1438 a_17100_2767# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1439 a_21545_10633# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1440 a_15371_5309# _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1441 _042_ net22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1442 a_22937_8457# tdc1.w_ring_int_norsz[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1443 VGND tdc0.r_ring_ctr[5] _147_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1444 a_12353_14977# a_12135_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1445 a_6798_9813# a_6630_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1446 VPWR _084_ a_25264_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1447 a_12242_5309# a_11803_4943# a_12157_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1449 a_10037_13647# a_9871_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1450 a_28467_12393# a_28338_12137# a_28047_12247# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1451 a_17751_3829# _057_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1452 a_9163_14191# a_8381_14197# a_9079_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1453 VPWR net28 a_7295_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1454 tdc0.r_dly_store_ring[1] a_20655_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1455 a_20966_5055# a_20798_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1457 a_17576_3855# a_16661_3855# a_17229_4097# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1458 net19 a_27411_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1459 a_11517_12809# _075_ a_11601_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1460 a_19535_7637# _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X1461 tdc0.w_ring_buf[23] a_7755_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1462 a_17578_12925# a_17139_12559# a_17493_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1465 a_3521_14191# _158_ a_3439_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1466 a_14683_10927# a_13901_10933# a_14599_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1467 net32 a_17100_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1468 VPWR a_20223_13799# tdc0.r_dly_store_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1469 a_24849_7663# a_24315_7669# a_24754_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1470 a_2490_11059# a_2768_11043# a_2724_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1472 tdc0.w_ring_norsz[14] tdc0.w_ring_norsz[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1473 VGND a_12007_13077# a_11965_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1474 a_6246_10495# a_6078_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1475 VGND a_26983_8207# net41 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1478 tdc0.r_dly_store_ctr[15] a_4463_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1479 VPWR net35 a_23211_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1480 a_26251_11471# _098_ a_26420_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1481 VGND a_9247_14165# a_9205_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1482 _031_ a_14951_3855# a_15189_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X1483 net9 a_18059_16375# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1485 a_15289_10927# tdc0.r_dly_store_ring[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1486 _111_ a_20065_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X1487 VPWR a_24075_13103# a_24243_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1488 a_21178_12809# _089_ a_21095_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
X1490 a_25179_7663# a_24481_7669# a_24922_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1491 _003_ a_3439_14191# a_3689_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1492 VGND a_24075_13103# a_24243_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1493 a_29541_7485# a_29007_7119# a_29446_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1495 a_5529_14013# a_4995_13647# a_5434_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1497 _196_ a_8399_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1498 a_24209_14735# tdc0.r_ring_ctr[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1499 a_25309_5487# a_24775_5493# a_25214_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1500 VPWR net37 a_23671_15287# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1501 _030_ _175_ a_12981_3631# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X1502 a_17233_7369# tdc1.w_ring_int_norsz[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1503 VGND a_19567_14013# a_19735_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1504 a_14541_13647# a_13551_13647# a_14415_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1505 a_11785_14735# a_11619_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1506 VPWR a_27038_11989# a_26965_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1507 VPWR net29 a_13275_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1508 a_7442_6143# a_7274_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1509 VGND tdc1.w_ring_norsz[25] tdc1.w_ring_norsz[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1511 a_5602_13759# a_5434_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1512 VGND a_10291_4373# _181_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1515 VGND a_16826_9813# a_16784_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1516 a_8654_16075# a_8971_15965# a_8929_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1518 a_3024_8725# net26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1519 VPWR a_14139_14191# a_14307_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1520 VGND a_16771_8751# _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1521 _056_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1522 a_23742_5487# a_23303_5493# a_23657_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1524 VPWR a_28694_7637# a_28621_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1527 a_17567_15797# _041_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1528 _163_ tdc1.r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1529 a_13533_3317# a_13367_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1530 VPWR _081_ a_22351_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X1531 a_21157_13647# a_20610_13921# a_20810_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1532 a_13637_7983# _071_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X1534 a_4866_9813# a_4698_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1536 a_19291_10927# a_18593_10933# a_19034_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1538 tdc1.w_ring_norsz[27] tdc1.w_ring_int_norsz[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1539 a_12368_4943# a_11969_4943# a_12242_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1541 tdc1.r_dly_store_ring[12] a_28291_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1542 VPWR _064_ a_15159_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1543 a_16003_4917# _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1544 VGND tdc0.w_ring_int_norsz[22] tdc0.w_ring_norsz[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1545 _064_ a_16587_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1546 a_24075_13103# a_23211_13109# a_23818_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1549 a_12291_6183# tdc1.r_dly_store_ring[22] a_12437_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X1550 _192_ a_13551_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1551 a_12897_8751# tdc1.r_dly_store_ring[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1552 VPWR a_4880_14735# a_5055_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1553 _623_.X a_4588_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1554 VGND net32 a_18703_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1555 VGND net35 a_23855_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1558 a_21976_3677# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1559 VGND a_19959_15797# tdc0.r_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1560 a_8170_4399# a_7093_4405# a_8008_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1561 VGND a_17935_2741# tdc1.r_ring_ctr[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1562 tdc1.r_dly_store_ring[26] a_29119_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1563 a_27222_9813# a_27054_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1564 a_4774_6031# _062_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1565 a_24719_12015# a_23855_12021# a_24462_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1566 a_12207_14191# a_11509_14197# a_11950_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1567 VGND a_11035_3543# _169_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1568 VPWR net7 a_3339_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1569 a_14886_16189# a_13809_15823# a_14724_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1570 a_20253_14735# tdc0.r_ring_ctr[1] a_20165_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1571 a_16757_13103# tdc0.w_ring_buf[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1572 VGND net7 a_3339_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1573 a_15107_7779# _120_ a_15025_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1575 tdc0.w_ring_int_norsz[31] tdc0.w_ring_norsz[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1577 a_21743_6895# _113_ a_21912_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1578 VPWR tdc1.w_ring_norsz[27] a_28179_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1579 a_24389_12015# a_23855_12021# a_24294_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1580 a_7732_15657# a_6651_15285# a_7385_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1582 a_20629_6895# tdc1.r_dly_store_ctr[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1583 VGND a_22679_13915# a_22637_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1585 VPWR _067_ a_11601_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1586 VGND tdc1.w_ring_norsz[17] a_23855_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
R21 VGND net48 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1587 a_14139_14191# a_13275_14197# a_13882_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1588 a_27517_5493# a_27351_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1589 a_28289_12015# a_27951_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1592 VPWR a_21391_5211# a_21307_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1593 VGND tdc0.w_ring_norsz[17] a_15483_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1594 VGND _083_ a_25765_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1595 a_26055_9545# _097_ a_25973_9301# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1596 a_18039_14191# a_17415_14197# a_17931_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1597 a_10494_5309# a_10221_4943# a_10409_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1599 VPWR a_22719_10357# a_22726_10657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1600 a_9945_10927# a_9411_10933# a_9850_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1601 a_11277_3855# _168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1602 a_11706_12015# _124_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X1604 _000_ tdc0.r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1605 VPWR _064_ a_18501_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X1608 a_10087_10411# tdc0.r_dly_store_ring[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1609 a_28621_7663# a_28087_7669# a_28526_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1610 a_3789_13897# tdc0.r_ring_ctr[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.153 ps=1.3 w=1 l=0.15
X1611 VGND net31 a_18427_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1612 VGND net7 a_8123_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1613 a_23960_14569# a_23561_14197# a_23834_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1614 a_14431_4373# _175_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X1615 VPWR tdc1.w_ring_int_norsz[3] a_23469_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1617 a_11785_14735# a_11619_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1618 VPWR net25 a_14011_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1619 tdc0.r_ring_ctr[10] a_18671_14495# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1620 a_21997_15285# a_21831_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1621 VPWR a_3484_13077# net21 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1622 a_14442_9295# _189_ a_13620_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1623 tdc1.w_ring_buf[12] a_27167_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1624 VGND a_15809_12234# tdc0.w_ring_buf[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1625 a_23868_5865# a_23469_5493# a_23742_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1626 VPWR a_20471_5461# a_20387_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1627 a_17578_12925# a_17305_12559# a_17493_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1628 a_27215_11293# a_26995_11305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
R22 net73 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1630 tdc0.w_ring_norsz[18] net24 a_23021_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1631 a_13990_13103# a_13717_13109# a_13905_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1632 a_13707_8867# _187_ a_13635_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1633 a_6357_9845# a_6191_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1634 _097_ a_22257_9545# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.172 ps=1.35 w=1 l=0.15
X1635 _067_ a_11987_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
R23 VGND uio_oe[4] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1637 a_29955_8983# tdc1.r_dly_store_ring[9] a_30101_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1638 VPWR a_8183_4703# tdc1.r_ring_ctr[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1639 a_24845_14735# a_23855_14735# a_24719_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1640 tdc0.w_ring_norsz[6] net21 a_11981_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1641 a_16935_16189# _041_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1642 a_8017_7663# tdc1.w_ring_buf[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1643 VGND a_9643_12724# tdc0.w_ring_buf[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1645 tdc0.w_ring_norsz[24] net21 a_8577_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1647 VGND a_12410_5055# a_12368_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1649 VPWR a_15504_9295# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1650 a_23305_8457# tdc1.w_ring_int_norsz[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1652 VGND net15 _062_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1653 a_4866_8725# a_4698_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1654 a_12447_13103# _077_ a_12529_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1655 a_6739_13897# _158_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1656 VGND net28 a_8767_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1657 VGND a_7867_6299# a_7825_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1658 tdc1.r_dly_store_ring[9] a_29487_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1659 VGND tdc0.r_ring_ctr[15] a_3255_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1660 tdc1.w_dly_stop[2] a_26891_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1661 tdc0.r_ring_ctr[4] a_12599_16671# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1662 a_16213_13647# a_15023_13647# a_16104_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1663 a_10275_12015# a_9577_12021# a_10018_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1664 a_9447_5309# a_8583_4943# a_9190_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1666 VPWR tdc1.w_ring_norsz[1] a_23119_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1668 VPWR a_18243_8751# _081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1669 a_19789_12559# a_19623_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1671 a_20789_4765# tdc1.r_ring_ctr[1] a_20717_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1672 a_19693_4943# a_18703_4943# a_19567_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1674 VGND net3 a_9503_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1675 VGND net35 a_23119_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1677 VPWR a_7055_9839# a_7223_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1680 VPWR net19 a_26615_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1681 a_3621_5487# _184_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1682 VGND a_5291_8725# a_5249_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1683 tdc0.w_ring_int_norsz[18] net45 a_16961_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1684 a_9437_15823# a_9058_16189# a_9365_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1685 VGND a_2807_11169# a_2768_11043# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1686 a_8735_3689# a_8289_3317# a_8639_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1687 a_21891_15797# _033_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1689 tdc1.r_dly_store_ring[29] a_16331_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1690 VGND tdc1.w_ring_norsz[6] tdc1.w_ring_int_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1691 VGND tdc0.w_ring_norsz[6] tdc0.w_ring_int_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1692 a_13633_10383# tdc0.r_dly_store_ring[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1693 a_26329_6281# tdc1.r_dly_store_ring[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1694 VPWR a_19867_4703# a_19854_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1695 a_25593_10927# _086_ a_25511_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1696 a_24420_14735# a_24021_14735# a_24294_15101# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1697 VGND _164_ _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1698 a_16209_8751# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1699 a_23004_3855# a_21923_3855# a_22657_4097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1700 a_22569_10927# tdc0.w_ring_int_norsz[20] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1701 a_8569_14191# tdc0.r_ring_ctr[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1704 a_17739_7882# tdc1.w_ring_norsz[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1705 VGND a_27036_7637# net17 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1706 a_21905_13109# a_21739_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1707 a_3763_7119# a_3413_7119# a_3668_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1708 a_28299_5487# a_27517_5493# a_28215_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1709 a_25071_9813# _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X1710 a_8933_7485# a_8399_7119# a_8838_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1711 _066_ a_15335_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1712 VGND _093_ a_26251_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X1714 a_20947_6397# a_20083_6031# a_20690_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1715 VPWR _145_ a_10363_15617# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1717 tdc1.r_dly_store_ring[21] a_15871_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1719 VGND net34 a_23303_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1720 VPWR net31 a_20359_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1721 a_12073_8457# tdc1.w_ring_norsz[8] a_11989_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1722 a_19268_10383# a_18869_10383# a_19142_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1723 _107_ a_28731_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1724 VGND tdc1.w_ring_int_norsz[31] tdc1.w_ring_norsz[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1725 VPWR a_12575_10749# a_12743_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1726 VPWR a_26420_11721# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1727 a_7907_15583# a_7732_15657# a_8086_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1728 VPWR a_7385_15253# a_7275_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1730 tdc0.r_dly_store_ring[25] a_19735_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1731 a_22937_8751# tdc1.w_ring_int_norsz[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1732 VPWR a_4279_9563# a_4195_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1733 tdc1.w_ring_norsz[16] tdc1.w_ring_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1734 a_15829_7119# a_14839_7119# a_15703_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1735 VGND a_9459_8970# tdc1.w_ring_buf[23] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1736 a_8243_8751# a_7461_8757# a_8159_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1738 a_14899_15797# a_14724_15823# a_15078_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1739 VPWR a_7661_4373# a_7551_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1740 VPWR net28 a_8675_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1741 VPWR tdc1.w_ring_buf[18] a_22261_8041# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1742 tdc1.w_ring_int_norsz[24] net69 a_10797_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1745 VGND net5 a_16468_9111# VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
X1746 VPWR _070_ a_14332_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1747 a_25689_11247# tdc0.r_dly_store_ring[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1748 _068_ a_16309_8867# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1749 a_12058_9661# a_11619_9295# a_11973_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1750 VPWR _098_ a_26420_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X1751 VPWR a_23983_9839# a_24151_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1752 VPWR a_9539_13103# a_9707_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1753 a_17740_10071# tdc0.r_dly_store_ring[5] a_17882_9878# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1754 VPWR tdc0.w_ring_norsz[8] a_11435_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1755 VGND tdc0.w_ring_norsz[14] tdc0.w_ring_int_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1756 VPWR a_24903_6575# a_25071_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1757 VPWR a_6687_6575# a_6855_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1758 a_4220_14735# _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1759 VPWR a_16913_756# net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1760 a_28813_6575# _106_ a_28731_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1761 a_26697_6575# net18 tdc1.w_ring_norsz[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1763 VGND a_9539_13103# a_9707_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1764 VGND a_22511_14013# a_22679_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1766 a_9253_14763# tdc0.r_ring_ctr[6] a_9167_14763# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1767 VGND a_10018_10901# a_9976_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1768 a_26847_9460# tdc1.w_ring_norsz[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1770 VPWR tdc0.r_ring_ctr[9] a_15687_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X1771 a_18869_6281# tdc1.w_ring_norsz[29] a_18785_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1772 VPWR tdc0.r_ring_ctr[0] a_19805_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 tdc1.w_ring_norsz[18] tdc1.w_ring_norsz[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1775 net11 a_5271_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1778 a_5123_9839# a_4425_9845# a_4866_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1779 VPWR net32 a_17139_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1780 _045_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1783 VGND _067_ a_19141_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1784 tdc0.w_dly_stop[4] a_2879_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1785 a_5349_13647# tdc0.r_ring_ctr[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1787 a_12135_14735# a_11785_14735# a_12040_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1788 a_16853_7369# net19 tdc1.w_ring_norsz[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1789 VGND net5 a_16771_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1790 _066_ _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1791 a_8857_3285# a_8639_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1792 a_11764_16733# _010_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1793 VPWR net34 a_27259_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1794 VPWR a_23087_15583# a_23074_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1795 VPWR _196_ _051_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1796 VGND a_25179_7663# a_25347_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1797 VPWR net27 a_8215_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1799 _135_ a_10087_10411# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1800 a_24481_7669# a_24315_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1801 tdc1.r_dly_store_ring[23] a_9891_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1803 VPWR a_16003_4917# a_15990_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1806 VPWR a_9079_14191# a_9247_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1807 _141_ a_20727_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1808 VPWR a_10662_5055# a_10589_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1809 VPWR net13 a_7571_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1811 VGND a_9263_7485# a_9431_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1812 _127_ a_9963_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1813 VGND a_20763_11837# a_20931_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1814 _063_ net15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1816 _075_ a_14011_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1818 a_19310_5055# a_19142_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1819 a_3871_7485# a_3247_7119# a_3763_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1820 a_3785_10383# tdc0.r_ring_ctr[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1821 a_5342_11837# a_4903_11471# a_5257_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1822 VPWR a_16771_8751# _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1823 a_9539_13103# a_8675_13109# a_9282_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1825 a_5799_6031# tdc1.r_ring_ctr[14] a_5703_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X1826 VPWR a_14599_10927# a_14767_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1827 VPWR a_19959_15797# a_19946_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1828 a_25731_14191# a_24867_14197# a_25474_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1829 _120_ a_13551_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X1830 tdc0.w_ring_int_norsz[2] net40 a_22389_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1832 a_17581_6575# tdc1.w_ring_norsz[5] a_17497_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1833 VPWR _160_ a_6364_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.195 ps=1.39 w=1 l=0.15
X1834 VPWR tdc0.r_dly_store_ring[25] a_19329_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X1835 tdc1.w_ring_int_norsz[27] net72 a_26529_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1836 VGND tdc0.w_ring_norsz[2] a_23855_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1837 VPWR net8 a_13367_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1838 VGND net25 a_13989_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1839 a_7718_14557# _045_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1840 VGND _181_ a_6105_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1841 a_23558_9839# a_23285_9845# a_23473_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1842 a_18869_15823# a_18703_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1843 a_17882_9878# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1844 a_15543_7895# _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X1845 a_9765_12015# tdc0.w_ring_buf[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1846 _195_ a_18703_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1848 a_24478_6575# a_24205_6581# a_24393_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1849 a_25472_8181# tdc1.r_dly_store_ring[3] a_25692_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
R24 VGND net42 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1850 a_24167_5487# a_23303_5493# a_23910_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1851 a_14457_12015# tdc0.w_ring_buf[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1852 a_6771_6575# a_5989_6581# a_6687_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1853 tdc0.w_ring_buf[26] a_27535_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1854 VGND a_9103_4659# net15 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1855 a_12184_9295# a_11785_9295# a_12058_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1856 VPWR _130_ a_11792_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X1857 uo_out[0] a_13620_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1859 a_25474_3967# a_25306_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1861 a_11343_15279# tdc0.r_ring_ctr[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X1862 a_12424_16745# a_11343_16373# a_12077_16341# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1865 VGND a_8527_9839# a_8695_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1866 a_11149_11721# _083_ a_11233_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1867 tdc0.r_dly_store_ring[8] a_12743_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1868 VPWR tdc0.w_dly_stop[4] a_3155_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1869 VPWR tdc0.w_ring_int_norsz[23] a_7829_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1870 tdc1.r_ring_ctr[8] a_14623_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X1871 a_17413_3009# a_17195_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1872 a_19801_4777# a_18611_4405# a_19692_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1873 a_9079_14191# a_8215_14197# a_8822_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1874 VPWR a_9615_5211# a_9531_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1876 a_9114_13103# a_8841_13109# a_9029_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1877 VGND a_12539_9839# _072_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1878 a_12157_4943# tdc1.r_ring_ctr[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1879 a_6799_14569# a_6449_14197# a_6704_14557# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1880 a_15772_9295# _122_ a_15504_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1881 a_25616_10633# _105_ a_25348_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1882 a_10337_16073# tdc0.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1883 a_20561_14013# a_20223_13799# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1884 VGND a_27866_6549# a_27824_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1885 VGND a_20503_15253# _143_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1886 a_16403_14557# tdc0.r_ring_ctr[10] a_16297_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1887 VPWR net20 _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1889 a_15653_6031# tdc1.w_ring_buf[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1890 tdc1.r_dly_store_ring[11] a_29119_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1891 a_25029_11305# a_24039_10933# a_24903_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1892 a_7853_11721# tdc0.w_ring_norsz[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1894 VGND a_7539_14495# a_7473_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1895 a_14599_10927# a_13735_10933# a_14342_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1896 tdc1.w_dly_stop[2] a_26891_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1897 a_8912_15599# a_8686_15395# a_8543_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1898 VGND net19 tdc1.w_ring_norsz[21] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1899 VPWR tdc0.w_ring_int_norsz[4] a_22273_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1901 VGND _075_ a_25121_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1903 a_24765_13897# _103_ a_24683_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1904 _070_ a_16771_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1905 a_8008_4777# a_7093_4405# a_7661_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1907 tdc0.w_ring_int_norsz[29] net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1908 VGND tdc0.w_ring_norsz[21] a_13459_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1909 a_8689_15823# a_8654_16075# a_8451_15797# VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X1911 a_14269_10927# a_13735_10933# a_14174_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1912 _040_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1914 VGND a_22695_5487# a_22863_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1916 VPWR _070_ a_18690_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1919 VGND net30 a_11803_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1920 a_14431_4373# tdc1.r_ring_ctr[8] a_14829_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X1921 a_10699_10633# _066_ a_10781_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1922 a_15105_13103# tdc0.r_dly_store_ctr[13] a_15023_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1924 a_23653_4405# a_23487_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1925 VGND tdc1.r_ring_ctr[12] a_6291_5193# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1926 VPWR a_12778_4373# a_12705_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1927 _104_ a_24683_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1928 VPWR a_13019_7637# a_12935_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1929 VPWR a_19345_4373# a_19235_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1931 a_10819_14013# a_10037_13647# a_10735_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1932 a_7091_4221# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1934 a_20690_6143# a_20522_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1936 VPWR a_12424_16745# a_12599_16671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1937 VPWR a_24427_14165# a_24343_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1939 a_5526_7485# a_5253_7119# a_5441_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1941 _132_ a_9871_7369# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1942 VPWR a_19459_6549# a_19375_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1943 a_24029_12809# tdc0.r_dly_store_ring[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1946 a_21445_9845# a_21279_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1947 a_16104_13647# a_15189_13647# a_15757_13889# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1948 a_17107_3855# a_16661_3855# a_17011_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1949 a_22657_4097# a_22439_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1951 a_7429_15645# a_7385_15253# a_7263_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1952 VGND _084_ _085_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1953 VPWR net26 a_3247_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1954 a_5043_10548# tdc0.w_ring_norsz[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1956 VGND a_12226_9407# a_12184_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1957 VPWR a_11299_6794# tdc1.w_ring_buf[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1958 VPWR net28 a_8859_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1960 tdc0.r_dly_store_ring[31] a_6671_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1961 VGND a_22346_13077# a_22304_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1962 a_3505_4943# a_3339_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1964 a_19789_12559# a_19623_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1965 VPWR a_11655_6397# a_11823_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1966 VPWR a_5231_4631# _020_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X1967 a_25373_10159# _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1968 uo_out[2] a_26420_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1970 a_27866_6549# a_27698_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1971 VPWR a_12700_14735# a_12875_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1972 a_17760_2767# a_16845_2767# a_17413_3009# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1973 a_10787_7369# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1974 net18 a_26615_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1976 a_4698_9839# a_4259_9845# a_4613_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1977 net3 a_855_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1978 tdc0.w_ring_norsz[22] tdc0.w_ring_norsz[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1979 a_22603_13103# a_21905_13109# a_22346_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
R25 VPWR tdc1.g_ring3[22].stg01_67.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1980 VPWR tdc1.r_dly_store_ctr[11] a_18501_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X1981 VPWR _195_ _040_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1982 VPWR tdc1.w_ring_norsz[0] a_5547_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1984 _170_ tdc1.r_ring_ctr[5] a_11895_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1985 VGND a_24094_4373# a_24052_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1988 VPWR a_7548_3855# a_7723_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1989 a_22346_13077# a_22178_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1990 a_25382_5461# a_25214_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1991 tdc0.w_ring_norsz[19] tdc0.w_ring_norsz[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1993 tdc0.r_dly_store_ring[30] a_9707_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1995 VGND _069_ a_15369_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1996 tdc0.r_dly_store_ring[30] a_9707_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1997 VGND net71 tdc1.w_ring_int_norsz[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1998 VGND a_14139_6575# a_14307_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1999 VGND _079_ a_25373_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2000 a_22178_13103# a_21905_13109# a_22093_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2001 VGND a_8399_3855# _196_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2002 a_19878_5487# a_19439_5493# a_19793_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2003 VGND a_21886_8725# a_21844_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2004 a_12705_4399# a_12171_4405# a_12610_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2005 a_24959_7119# _075_ a_25137_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X2006 VPWR a_29062_8725# a_28989_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2007 VGND tdc0.w_ring_norsz[0] a_5271_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2009 a_7473_14569# a_6283_14197# a_7364_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2010 a_21399_10535# tdc0.r_dly_store_ring[12] a_21545_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2012 a_11859_16745# a_11343_16373# a_11764_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2013 a_6791_11636# tdc0.w_ring_norsz[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2014 a_8105_12021# a_7939_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2016 _621_.X a_3024_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2017 a_16182_4943# _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2019 _125_ a_11067_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2020 a_9924_14165# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2021 a_9941_7983# tdc1.r_dly_store_ring[23] a_9595_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2023 a_10583_4765# _173_ a_10487_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X2024 a_22381_14977# a_22163_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2026 VGND net41 a_27351_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2027 VGND a_27411_7093# net19 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2028 VGND a_15871_7387# a_15829_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2029 a_12751_5309# a_11969_4943# a_12667_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2030 a_26575_11159# a_26859_11145# a_26794_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2032 VGND a_19255_14735# net22 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2033 a_14139_14191# a_13441_14197# a_13882_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2035 a_19437_16065# a_19219_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2036 VPWR a_20931_11739# a_20847_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2037 a_27479_9839# a_26615_9845# a_27222_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2038 tdc0.w_ring_buf[18] a_26063_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2040 a_14921_14735# _152_ _157_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2042 VPWR a_23726_9813# a_23653_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2043 a_23926_4399# a_23487_4405# a_23841_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2044 a_13178_5853# a_12863_5719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2046 a_14279_10633# _192_ a_14197_10389# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2047 a_11877_14191# a_11343_14197# a_11782_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2048 VPWR a_24646_6549# a_24573_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2049 a_23983_9839# a_23285_9845# a_23726_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2051 VGND tdc1.r_ring_ctr[4] a_16135_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2052 VPWR a_18003_8573# a_18171_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2053 a_21009_12015# tdc0.w_ring_norsz[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2054 VGND tdc0.w_dly_stop[4] a_3155_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2055 a_5823_8457# tdc1.w_ring_int_norsz[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2056 VPWR a_24335_5461# a_24251_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2057 a_23004_3855# a_22089_3855# a_22657_4097# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2058 tdc1.w_ring_int_norsz[31] net76 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2059 a_5905_12015# net20 tdc0.w_ring_norsz[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2060 VPWR a_14951_3855# _031_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X2061 _164_ a_20635_4512# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2062 a_24109_10217# a_23119_9845# a_23983_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2063 a_19124_15823# _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2064 VPWR tdc1.w_ring_norsz[28] a_27075_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2065 net38 a_16463_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2066 a_7645_6575# tdc1.w_ring_norsz[31] a_7561_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2067 VGND net32 a_17139_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2069 a_7181_12559# a_6191_12559# a_7055_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2070 _053_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2071 VGND tdc0.w_ring_int_norsz[7] tdc0.w_ring_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2072 a_7093_4405# a_6927_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2074 a_9347_7485# a_8565_7119# a_9263_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2075 a_24094_4373# a_23926_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2076 _034_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2077 VPWR tdc1.w_ring_norsz[17] a_24305_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2078 a_8577_10927# tdc0.w_ring_norsz[8] a_8493_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R26 VGND net43 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2080 VGND a_14623_3615# a_14557_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2081 a_12529_13103# tdc0.r_dly_store_ctr[12] a_12447_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2082 tdc1.w_ring_norsz[30] net16 a_14649_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2084 a_22990_3677# _049_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2085 VPWR a_29587_7895# _101_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X2086 VPWR _069_ a_25677_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X2088 a_21813_14735# a_21647_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2089 VGND a_24922_7637# a_24880_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2092 VPWR net10 a_13643_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2093 a_14145_3677# a_14101_3285# a_13979_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2094 _195_ a_18703_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2096 VGND a_29487_8725# a_29445_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2097 VGND net29 a_11343_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2098 a_15647_14013# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2099 VGND a_22143_8751# a_22311_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2100 VPWR tdc0.w_ring_norsz[11] a_20441_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2101 VGND a_25382_5461# a_25340_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2102 VGND tdc1.w_ring_norsz[19] tdc1.w_ring_int_norsz[20] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2103 a_27613_6575# tdc1.w_ring_buf[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2104 a_21327_7895# a_21423_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2105 net30 a_11763_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2106 VPWR ui_in[1] a_855_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2107 a_20004_5865# a_19605_5493# a_19878_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2108 VGND net23 tdc0.w_ring_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2109 tdc0.w_dly_stop[1] a_2327_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2110 _196_ a_8399_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2111 net35 a_23080_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2112 a_22595_14013# a_21813_13647# a_22511_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2113 a_29035_9839# a_28253_9845# a_28951_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2115 tdc1.w_ring_int_norsz[13] net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2116 VGND a_24276_9269# net34 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2119 a_24485_8751# tdc1.w_ring_buf[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2120 _165_ a_21279_4765# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X2121 a_23653_9839# a_23119_9845# a_23558_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2122 VGND a_20303_5487# a_20471_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2125 a_24573_6575# a_24039_6581# a_24478_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2126 a_6357_6575# a_5823_6581# a_6262_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2127 VPWR _064_ a_19329_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X2128 VPWR tdc1.w_ring_norsz[24] a_12345_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2130 a_9693_16367# _148_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2131 a_17195_4777# a_16845_4405# a_17100_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2132 a_12700_14735# a_11785_14735# a_12353_14977# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2133 VPWR a_9447_5309# a_9615_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2134 VGND net13 tdc1.w_ring_int_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2135 a_14158_13077# a_13990_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2136 VPWR a_5694_7231# a_5621_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2137 a_10363_15617# _143_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2138 a_3413_7119# a_3247_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2139 a_13441_14197# a_13275_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2140 VPWR a_17935_2741# a_17922_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2141 a_12437_6281# _075_ a_12291_6183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X2142 VGND a_16135_3311# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X2143 a_6027_9622# tdc0.r_dly_store_ring[7] a_6027_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2145 a_11885_7369# net68 tdc1.w_ring_int_norsz[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2146 a_25677_10927# tdc0.r_dly_store_ring[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2147 a_19567_5309# a_18703_4943# a_19310_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2148 a_12575_10749# a_11877_10383# a_12318_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2149 a_7139_12925# a_6357_12559# a_7055_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2150 net27 a_2932_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2151 a_21279_4765# tdc1.r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X2152 a_15189_3855# tdc1.r_ring_ctr[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2154 VGND a_21511_9447# _112_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X2155 a_17302_5487# a_16863_5493# a_17217_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2156 a_17045_16065# a_16827_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2157 VPWR tdc0.w_ring_norsz[11] a_21739_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2158 a_20223_13799# a_20319_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2160 a_7274_6397# a_7001_6031# a_7189_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2162 tdc0.w_ring_buf[11] a_21739_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2163 a_12040_14735# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2165 VPWR _179_ _180_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2168 a_20531_3855# tdc1.r_ring_ctr[0] _163_ VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2169 VGND _083_ a_14090_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2170 a_20249_6031# a_20083_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2171 a_8270_9813# a_8102_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2173 VPWR net27 a_5639_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2175 VGND a_3392_8725# _620_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2176 VPWR a_10275_10927# a_10443_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2177 a_12403_8970# tdc1.w_ring_norsz[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2178 a_15687_15823# _153_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2179 VGND net20 tdc0.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2180 a_6798_12671# a_6630_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2181 VPWR tdc1.w_dly_stop[3] a_27167_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2182 VGND a_7055_12925# a_7223_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2183 VGND _131_ a_10241_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2184 _070_ a_16771_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2186 VGND a_19735_10651# a_19693_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2187 a_21813_14735# a_21647_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2188 _622_.X a_2840_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2190 VGND net31 a_19439_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2192 VPWR a_9127_16060# a_9058_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X2193 a_3760_4943# _020_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
R27 VPWR tdc1.g_ring3[28].stg01_73.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2194 VPWR a_24351_4399# a_24519_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2196 VGND net30 a_11619_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2197 a_5507_6005# tdc1.r_ring_ctr[12] a_5905_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X2198 a_18593_10933# a_18427_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2200 VGND _195_ _033_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2201 a_9577_12021# a_9411_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2202 VGND a_12731_3311# _030_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X2203 a_27180_10217# a_26781_9845# a_27054_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2204 a_12121_16733# a_12077_16341# a_11955_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2205 a_16477_15823# a_16311_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2206 a_9551_15511# tdc0.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2207 _054_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2208 a_21833_10383# _072_ a_21399_10535# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2209 VGND net9 a_3799_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2210 VGND a_7810_13077# a_7768_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2212 VPWR net23 _043_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2213 net15 a_9103_4659# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2214 a_5621_7485# a_5087_7119# a_5526_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2215 a_12815_8751# _067_ a_12897_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2216 VGND a_14599_10927# a_14767_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2217 a_14269_12021# a_14103_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2219 a_23385_7369# net17 tdc1.w_ring_norsz[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2220 VPWR tdc1.w_ring_norsz[16] a_6743_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2221 a_21633_8751# tdc1.w_ring_buf[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2223 a_7275_15279# a_6651_15285# a_7167_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2225 a_12567_9661# a_11785_9295# a_12483_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2226 a_19683_3689# a_19237_3317# a_19587_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2227 a_17303_4399# a_16679_4405# a_17195_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2228 VPWR a_27647_9813# a_27563_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2229 VPWR a_9503_9295# _086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2232 _007_ tdc0.r_ring_ctr[1] a_19973_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2233 a_25474_3967# a_25306_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2235 VGND net28 a_8859_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2236 a_8544_3677# _028_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2237 net40 a_27351_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2238 a_6629_10383# a_5639_10383# a_6503_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2239 a_10275_10927# a_9411_10933# a_10018_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2240 tdc1.r_dly_store_ring[12] a_28291_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2241 VPWR tdc1.r_ring_ctr[10] a_14431_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X2242 a_21644_9295# _081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2243 tdc0.r_dly_store_ctr[6] a_10903_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2244 a_17428_5865# a_17029_5493# a_17302_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2245 a_13839_7663# tdc1.r_dly_store_ctr[8] a_13637_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2246 VPWR _077_ a_13645_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2247 _150_ a_9167_14763# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X2248 a_28441_9839# tdc1.w_ring_buf[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
R28 VGND uio_oe[3] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2249 a_25731_14191# a_25033_14197# a_25474_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2250 a_13905_13647# tdc0.r_ring_ctr[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2251 a_8293_12015# tdc0.w_ring_buf[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2252 a_21637_9545# _081_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X2253 VPWR a_15504_9295# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2254 a_16961_12015# tdc0.w_ring_norsz[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2256 a_29173_7119# a_29007_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2257 _113_ a_20729_9955# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X2258 VGND net25 a_13897_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2259 a_23834_14191# a_23561_14197# a_23749_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2260 VPWR a_12539_9839# _072_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2261 a_3668_12559# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2262 a_5277_7663# net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2263 a_11989_8457# tdc1.w_ring_int_norsz[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2264 a_14655_8751# _065_ a_14909_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2267 _055_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2268 a_17555_7284# tdc1.w_ring_norsz[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2269 VGND _070_ a_19631_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2270 VGND a_12539_9839# _072_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2271 _052_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2272 a_25125_7369# tdc1.r_dly_store_ring[19] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2274 a_7364_14569# a_6449_14197# a_7017_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2275 a_22439_3855# a_21923_3855# a_22344_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2276 a_7829_10927# tdc0.w_ring_norsz[7] a_7745_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2277 VPWR a_17283_14709# net33 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2278 VPWR a_5602_13759# a_5529_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R29 VGND uio_oe[2] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2280 a_11969_4943# a_11803_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2281 a_17029_5493# a_16863_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2282 tdc1.w_ring_norsz[29] tdc1.w_ring_norsz[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2283 VPWR _135_ a_11131_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2284 VGND a_19066_7895# _128_ VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X2285 VGND tdc1.w_ring_norsz[1] a_23119_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2286 VPWR a_10124_9269# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2287 a_20062_12925# a_19623_12559# a_19977_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2288 tdc1.w_ring_buf[27] a_28179_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2289 a_21279_7119# _075_ a_21457_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X2290 a_9871_7369# _076_ a_9953_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2291 VPWR net6 a_16771_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2292 a_15333_9545# _083_ a_15504_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2293 a_23080_14165# net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2294 a_28694_7637# a_28526_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2295 VGND net27 a_4259_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2297 a_17118_9661# a_16845_9295# a_17033_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2298 a_11582_13077# a_11414_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2300 a_12337_5309# a_11803_4943# a_12242_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2301 VGND _108_ a_21743_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2302 _083_ a_20083_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2304 VGND _086_ a_25327_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2305 VPWR tdc0.w_ring_int_norsz[16] a_5989_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2306 VPWR tdc0.w_ring_norsz[30] a_8583_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2307 a_8822_14165# a_8654_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2308 a_9079_14191# a_8381_14197# a_8822_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2312 VGND a_24151_9813# a_24109_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2313 net37 a_3247_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2314 VPWR a_8527_9839# a_8695_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2315 a_28266_12381# a_27951_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2318 a_8117_4777# a_6927_4405# a_8008_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2319 a_24669_7663# tdc1.w_ring_buf[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2320 a_26965_12015# a_26431_12021# a_26870_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2321 VGND a_4866_9813# a_4824_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2323 _066_ a_15335_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2324 a_16845_4405# a_16679_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2325 a_22798_3311# a_21721_3317# a_22636_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2326 _620_.X a_3392_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2328 tdc0.w_ring_norsz[2] net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2329 a_13441_12015# tdc0.w_ring_norsz[29] a_13357_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2330 VPWR net9 a_3799_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2332 _123_ a_10147_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2333 a_22339_10535# a_22435_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2334 _028_ _172_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2336 _194_ a_5015_9622# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
R30 tt_um_hpretl_tt06_tdc_v2_85.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2337 tdc1.r_dly_store_ring[7] a_5291_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2339 tdc1.r_dly_store_ctr[2] a_21391_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2340 VGND a_5871_11146# tdc0.w_ring_buf[31] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2341 tdc1.r_ring_ctr[2] a_19867_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2342 VPWR a_19735_5211# a_19651_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2343 a_26789_8457# net40 tdc1.w_ring_int_norsz[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2344 tdc1.w_ring_norsz[10] tdc1.w_ring_int_norsz[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2346 a_12599_16671# _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2347 VPWR net15 _060_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2348 a_14471_5807# _178_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X2349 VPWR a_20763_11837# a_20931_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2350 VPWR a_10018_10901# a_9945_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2352 a_4698_8751# a_4259_8757# a_4613_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2353 VPWR a_8971_11989# a_8887_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2354 VGND a_25474_13077# a_25432_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2355 a_24351_4399# a_23487_4405# a_24094_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2356 VGND net34 a_24775_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2357 a_22163_14735# a_21813_14735# a_22068_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2358 a_13119_4399# a_12337_4405# a_13035_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2359 net26 a_3115_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2360 VPWR a_14710_11989# a_14637_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2361 a_24205_6581# a_24039_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2362 VPWR a_7442_6143# a_7369_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2363 a_14913_4943# a_14747_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2366 a_25731_13103# a_25033_13109# a_25474_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2367 VGND tdc0.w_ring_norsz[8] a_11435_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2368 a_23845_7663# net40 tdc1.w_ring_int_norsz[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2369 a_3854_8319# a_3686_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2370 VGND a_16913_756# net4 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2372 a_4490_12925# a_3413_12559# a_4328_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2374 VPWR a_17727_5487# a_17895_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2376 VGND a_15023_5487# net8 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2377 a_25474_13077# a_25306_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2379 a_15420_9295# _121_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2380 a_17682_13621# a_17482_13921# a_17831_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2381 VPWR tdc1.w_ring_norsz[13] a_13265_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2382 VPWR tdc0.w_ring_norsz[19] a_22557_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2383 VGND a_30039_8475# a_29997_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2384 a_8527_9839# a_7663_9845# a_8270_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2386 tdc0.w_dly_stop[4] a_2879_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2387 a_5851_11837# a_5069_11471# a_5767_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2388 VPWR tdc1.w_dly_stop[1] a_26891_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2389 a_18690_8751# _065_ _081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X2390 VPWR _064_ a_20065_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X2391 a_7139_9839# a_6357_9845# a_7055_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2392 tdc0.r_dly_store_ring[8] a_12743_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2393 a_2840_12533# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2394 a_15719_10357# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2395 VGND tdc1.w_dly_stop[3] a_27167_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2397 VPWR tdc1.r_ring_ctr[12] a_5635_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2398 a_24213_6281# tdc1.r_dly_store_ctr[9] a_24131_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2399 a_11141_13109# a_10975_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2400 tdc1.r_dly_store_ring[28] a_28383_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R31 tdc1.g_ring3[31].stg01_76.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2401 _087_ a_19329_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X2403 a_8381_14197# a_8215_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2404 a_25033_14197# a_24867_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2406 tdc0.r_dly_store_ring[0] a_4279_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2407 a_21373_12015# tdc0.w_ring_int_norsz[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2409 a_3413_7119# a_3247_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2410 a_6630_9839# a_6191_9845# a_6545_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2411 VGND a_20471_5461# a_20429_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2412 a_21073_6031# a_20083_6031# a_20947_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2413 _072_ a_12539_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2414 a_17493_12559# tdc0.w_ring_buf[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2415 VPWR a_13511_7895# _188_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X2418 VGND tdc1.r_ring_ctr[3] a_21555_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X2419 VGND tdc0.w_ring_int_norsz[16] tdc0.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2421 tdc0.r_ring_ctr[1] a_21891_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2422 a_13717_13109# a_13551_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2423 VGND a_12587_8372# tdc1.w_ring_buf[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2424 _012_ _149_ a_9693_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2426 VPWR a_25472_8181# _102_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X2427 a_11073_8457# tdc1.w_ring_norsz[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2429 VGND a_24903_6575# a_25071_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2430 VGND a_6687_6575# a_6855_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2431 a_20083_14735# tdc0.r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2432 VGND a_20327_3615# a_20261_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2434 a_19417_11305# a_18427_10933# a_19291_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
R32 tt_um_hpretl_tt06_tdc_v2_83.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
R33 VPWR tdc1.g_ring3[27].stg01_72.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2436 a_17291_2767# a_16845_2767# a_17195_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2437 VGND a_5043_8372# tdc1.w_ring_buf[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2438 a_4824_9129# a_4425_8757# a_4698_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2441 VGND a_14307_6549# a_14265_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2442 _066_ _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X2443 a_11967_16367# _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2445 a_11393_14763# tdc0.r_ring_ctr[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2446 a_22435_10357# a_22719_10357# a_22654_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2447 _077_ a_9963_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2448 net38 a_16463_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2450 a_23113_3855# a_21923_3855# a_23004_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2452 VGND _195_ _037_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2453 a_23745_13103# a_23211_13109# a_23650_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2454 a_19567_14013# a_18869_13647# a_19310_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2458 tdc0.w_ring_buf[26] a_27535_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2459 a_8723_11636# tdc0.w_ring_norsz[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2460 VGND _100_ a_25472_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2461 VPWR a_27769_5108# tdc1.w_dly_stop[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2462 VPWR tdc1.w_ring_norsz[30] a_8849_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2463 a_24067_9839# a_23285_9845# a_23983_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2464 a_25639_5487# a_24775_5493# a_25382_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2466 tdc1.w_ring_norsz[14] tdc1.w_ring_norsz[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2467 a_20359_14735# tdc0.r_ring_ctr[2] a_20253_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X2468 VGND net17 tdc1.w_ring_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2469 uo_out[7] a_10124_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2470 a_19605_10205# _070_ a_19505_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X2472 a_15539_13647# a_15189_13647# a_15444_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2473 a_8565_7119# a_8399_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2474 a_15772_9295# _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2475 a_15738_6397# a_15465_6031# a_15653_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2476 VGND tdc1.w_ring_norsz[17] tdc1.w_ring_norsz[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2477 _039_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2479 a_19141_13423# tdc0.r_dly_store_ring[17] a_18795_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2480 tdc0.r_dly_store_ring[31] a_6671_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2481 VPWR tdc0.w_ring_norsz[18] a_23569_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2483 a_29614_8319# a_29446_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2484 VPWR a_17286_9407# a_17213_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2485 a_24646_10901# a_24478_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2486 a_12594_7637# a_12426_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2487 VGND net10 a_21647_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2489 a_29614_8319# a_29446_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2490 a_18777_4405# a_18611_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2491 tdc1.w_ring_norsz[16] net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2492 a_10229_9839# tdc0.r_dly_store_ring[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2493 VGND net9 a_18703_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2495 a_20522_6397# a_20249_6031# a_20437_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2496 a_24478_10927# a_24205_10933# a_24393_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2497 VGND net35 a_24039_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2498 uo_out[3] a_25348_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2499 a_11209_3649# _168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2500 uo_out[0] a_13620_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2501 VGND net35 a_24867_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2502 VGND _036_ a_12121_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2503 a_12913_10927# tdc0.w_ring_norsz[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2505 a_11599_3133# a_10975_2767# a_11491_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2506 VGND tdc0.w_ring_norsz[5] tdc0.w_ring_int_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2508 VGND a_9551_15511# _148_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2509 tdc0.w_ring_int_norsz[8] tdc0.w_ring_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2510 VGND a_24167_5487# a_24335_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2511 a_13714_14191# a_13441_14197# a_13629_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2512 VPWR tdc1.w_ring_int_norsz[19] a_24021_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2513 VPWR tdc0.w_ring_int_norsz[30] a_12613_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2515 tdc1.r_ring_ctr[9] a_17751_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X2517 VPWR a_22728_14735# a_22903_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2518 a_15925_15823# tdc0.r_ring_ctr[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2519 _140_ tdc0.r_ring_ctr[0] a_19798_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X2520 a_29173_7119# a_29007_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2521 _084_ net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2524 VGND a_15627_14709# _155_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X2525 VPWR a_23818_13077# a_23745_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2526 VGND net29 a_13275_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2527 VPWR _166_ a_16385_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2529 a_25264_10633# _102_ a_25348_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2530 a_17501_15823# a_16311_15823# a_17392_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2531 tdc1.w_ring_buf[16] a_7111_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2532 a_17746_12671# a_17578_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2533 tdc0.r_dly_store_ring[0] a_4279_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2534 tdc0.w_ring_norsz[0] tdc0.w_ring_norsz[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2535 net10 a_14983_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2536 a_5043_10548# tdc0.w_ring_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2538 a_21445_7369# tdc1.r_dly_store_ring[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2541 a_17869_4777# a_16679_4405# a_17760_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2544 tdc1.r_dly_store_ring[11] a_29119_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2545 a_8857_3285# a_8639_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2548 a_11753_2767# a_11709_3009# a_11587_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2549 VGND a_10275_10927# a_10443_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2550 VGND net52 tdc0.w_ring_int_norsz[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2551 a_28951_7663# a_28087_7669# a_28694_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2552 VGND a_10478_13759# a_10436_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2553 a_5123_8751# a_4425_8757# a_4866_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2554 a_17213_9661# a_16679_9295# a_17118_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2556 VGND a_11299_6794# tdc1.w_ring_buf[22] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2557 net3 a_855_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2558 a_26817_10927# a_26479_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2559 a_14415_14013# a_13717_13647# a_14158_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2560 VPWR net30 a_12171_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2561 a_22185_5487# tdc1.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2562 VPWR a_8695_9813# a_8611_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2563 tdc0.r_dly_store_ring[17] a_17435_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2564 VGND a_12778_4373# a_12736_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2565 a_10229_10159# tdc0.r_dly_store_ctr[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2566 VPWR tdc1.r_ring_ctr[8] a_12813_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2567 VPWR tdc0.w_ring_norsz[5] a_16219_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2568 VPWR a_19567_5309# a_19735_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2569 a_4595_6005# _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2570 VPWR _069_ a_28897_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X2571 VPWR net10 a_21647_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2572 VPWR net7 a_6927_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2574 tdc0.w_ring_buf[5] a_16219_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2576 tdc1.r_dly_store_ring[20] a_25807_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2577 a_10045_5807# tdc1.r_dly_store_ctr[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2578 _044_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2579 tdc0.w_ring_int_norsz[21] net48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2580 VGND tdc1.w_dly_stop[1] a_26891_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2581 VPWR net32 a_18427_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2582 a_11509_14197# a_11343_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2583 _033_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2584 a_16577_7369# net39 tdc1.w_ring_int_norsz[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2585 a_16163_6397# a_15465_6031# a_15906_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2586 a_6791_11636# tdc0.w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2588 tdc0.r_dly_store_ctr[4] a_12375_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2590 VPWR a_24995_8751# a_25163_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2591 VGND net8 a_16679_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2592 tdc1.w_ring_buf[2] a_21003_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2593 VPWR tdc0.w_ring_int_norsz[0] a_5437_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2594 VPWR net15 _061_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2595 a_11396_2767# _027_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2598 a_15479_11721# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2599 VPWR a_29871_8573# a_30039_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2600 uo_out[6] a_11792_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2601 VPWR _174_ a_11067_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2602 a_11785_9295# a_11619_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2603 a_16301_7983# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X2604 a_26329_6031# tdc1.r_dly_store_ctr[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2605 VPWR tdc1.w_ring_norsz[31] a_7295_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2606 net19 a_27411_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2609 VPWR tdc0.w_dly_stop[3] a_2879_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2610 a_15283_8457# a_15335_8181# _066_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2611 a_17351_13103# a_16569_13109# a_17267_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
R34 net54 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2616 VPWR a_9190_5055# a_9117_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2617 VPWR _165_ a_21923_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2618 a_19066_7895# tdc1.r_dly_store_ring[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X2619 a_15479_11721# _086_ a_15261_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2620 a_21997_15285# a_21831_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2622 VPWR net26 a_7663_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2623 VPWR _086_ a_5229_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2624 a_5249_10217# a_4259_9845# a_5123_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2625 a_23179_3829# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2627 a_3785_10383# tdc0.r_ring_ctr[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2628 a_5055_14709# _044_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2630 a_25221_3855# tdc1.r_ring_ctr[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2631 VPWR tdc1.w_ring_int_norsz[7] a_11693_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2632 VGND _099_ a_24959_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2633 VPWR a_25807_5461# a_25723_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2635 a_22745_3689# a_21555_3317# a_22636_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2636 a_12897_9071# tdc1.r_dly_store_ring[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2637 a_12313_3883# tdc1.r_ring_ctr[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2638 a_9204_3689# a_8123_3317# a_8857_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2639 VPWR tdc1.w_ring_int_norsz[5] a_17949_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2640 _092_ a_26891_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X2641 a_7364_14569# a_6283_14197# a_7017_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2642 a_18751_8359# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X2644 a_18114_2767# _052_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2645 a_14565_6281# tdc1.w_ring_int_norsz[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2646 VGND a_14158_13077# a_14116_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2647 VGND tdc1.w_ring_norsz[28] a_27075_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2648 tdc1.w_ring_int_norsz[16] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2651 VGND _069_ a_10493_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2652 VPWR a_15906_6143# a_15833_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2653 a_5229_9622# tdc0.r_dly_store_ring[0] a_5015_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X2654 VGND a_18171_12827# a_18129_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2656 VPWR net32 a_16219_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2658 _106_ a_26247_6281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2659 _078_ a_24131_6281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2660 _137_ a_9411_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2661 a_2963_10901# a_2807_11169# a_3108_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X2662 VGND a_14899_15797# tdc0.r_ring_ctr[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2663 a_22071_3689# a_21721_3317# a_21976_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2664 VGND a_27769_5108# tdc1.w_dly_stop[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2665 a_17931_14569# a_17415_14197# a_17836_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2668 a_23259_7882# tdc1.w_ring_norsz[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2669 tdc1.r_dly_store_ctr[6] a_11087_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2671 a_13883_3689# a_13367_3317# a_13788_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2672 VPWR _068_ a_10781_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2673 a_29181_9295# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X2674 a_28909_6895# tdc1.r_dly_store_ring[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X2675 a_15179_7779# _119_ a_15107_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2676 a_4437_7119# a_3247_7119# a_4328_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2678 _009_ _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2679 _007_ a_19723_15279# a_19973_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X2680 a_15369_13423# tdc0.r_dly_store_ring[29] a_15023_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2681 VPWR a_20690_6143# a_20617_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2682 a_26996_12393# a_26597_12021# a_26870_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2683 a_15263_4943# a_14913_4943# a_15168_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2684 VPWR _177_ a_15649_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2685 VGND a_16771_8751# _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
R35 VPWR tdc0.g_ring3[31].stg01_58.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2687 VPWR tdc1.w_ring_norsz[3] a_24223_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2688 a_21718_9839# a_21279_9845# a_21633_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2689 a_3597_10383# a_3431_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2690 a_3601_8207# net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2692 tdc0.w_dly_stop[1] a_2327_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2693 VPWR a_7055_12925# a_7223_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2694 tdc1.w_ring_norsz[16] net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2695 a_24719_15101# a_24021_14735# a_24462_14847# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2696 VGND a_12375_14165# a_12333_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2697 a_21511_9447# tdc0.r_dly_store_ring[4] a_21751_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X2698 a_25755_8751# _078_ _079_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
R36 net52 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2699 a_11349_3855# _166_ a_11277_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2700 _071_ _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2701 VPWR _047_ a_3108_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X2702 tdc0.w_ring_norsz[31] tdc0.w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2704 a_16842_13103# a_16403_13109# a_16757_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2705 VGND a_2287_10901# tdc0.r_ring_ctr[15] VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2706 a_12065_10383# tdc0.w_ring_buf[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2707 a_13357_12015# net23 tdc0.w_ring_norsz[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2709 VPWR tdc0.w_ring_int_norsz[1] a_16385_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2710 tdc1.r_dly_store_ring[9] a_29487_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2711 net31 a_17323_8759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2712 _077_ a_9963_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2713 VGND tdc0.w_ring_int_norsz[3] tdc0.w_ring_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2715 a_12403_8970# tdc1.w_ring_norsz[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2716 a_4533_14977# a_4315_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2717 a_17923_12234# tdc0.w_ring_norsz[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2718 a_16916_3855# _031_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2722 a_8565_7119# a_8399_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2723 VPWR tdc0.r_dly_store_ring[28] a_20065_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X2724 VGND a_26859_11145# a_26866_11049# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2725 a_28894_8751# a_28455_8757# a_28809_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2726 tdc0.r_ring_ctr[0] a_19959_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X2727 VGND _070_ a_19991_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2728 a_15833_6397# a_15299_6031# a_15738_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2731 VGND a_6798_9813# a_6756_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2732 a_13629_6575# tdc1.w_ring_buf[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2733 a_13620_9269# _194_ a_14090_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2734 a_4866_9813# a_4698_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2735 a_8749_14191# a_8215_14197# a_8654_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2736 VPWR tdc0.r_ring_ctr[13] a_3789_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X2737 a_4073_5185# a_3855_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2738 VGND _196_ _055_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2741 a_20713_4943# tdc1.r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2742 a_3859_7119# a_3413_7119# a_3763_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2743 _022_ a_2519_7369# a_2769_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X2744 VPWR a_11115_4007# _171_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2745 a_12700_14735# a_11619_14735# a_12353_14977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2749 a_19492_3677# _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2750 a_9631_6397# a_8933_6031# a_9374_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2751 a_10919_5309# a_10055_4943# a_10662_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2753 VPWR _166_ a_11035_3543# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2754 a_13990_14013# a_13551_13647# a_13905_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2756 a_14800_6549# tdc1.w_dly_stop[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
R37 VGND net64 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2757 VGND _133_ a_10241_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2758 tdc0.w_ring_buf[3] a_23763_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2759 VPWR a_19784_15823# a_19959_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2761 a_22093_13103# tdc0.w_ring_buf[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2762 VGND tdc1.w_ring_norsz[16] a_6743_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2763 tdc0.w_ring_norsz[10] tdc0.w_ring_int_norsz[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2764 a_19237_3317# a_19071_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2765 a_17413_4373# a_17195_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2767 VGND a_13620_9269# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X2768 a_19245_11721# net41 tdc0.w_ring_int_norsz[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2769 a_28341_5865# a_27351_5493# a_28215_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2771 VGND a_13019_7637# a_12977_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2772 _021_ _185_ a_3621_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2774 a_20798_5309# a_20359_4943# a_20713_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2775 VPWR a_11219_14887# _145_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X2776 a_20157_7663# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X2777 a_29062_8725# a_28894_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2778 a_5767_11837# a_4903_11471# a_5510_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2779 a_16784_10217# a_16385_9845# a_16658_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2781 a_15371_5309# a_14747_4943# a_15263_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2782 VGND a_2932_14165# net27 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2783 a_15283_8457# _065_ a_15701_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2784 a_7929_6575# net15 tdc1.w_ring_norsz[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2786 tdc1.w_ring_norsz[25] net18 a_26701_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2787 VGND a_10443_11989# a_10401_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2788 VGND net29 a_10975_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2789 a_20445_4105# tdc1.r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2790 _100_ a_24959_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2791 VGND net34 a_27259_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2792 a_15787_7485# a_15005_7119# a_15703_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2793 a_5437_11837# a_4903_11471# a_5342_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2794 tdc1.r_dly_store_ring[22] a_11823_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2795 a_5993_10383# tdc0.w_ring_buf[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2796 VGND net27 a_8215_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2798 a_17392_15823# a_16477_15823# a_17045_16065# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2799 VGND a_7699_6397# a_7867_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2800 VGND _067_ a_25397_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X2801 tdc1.w_ring_int_norsz[19] tdc1.w_ring_norsz[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2802 a_18027_14569# a_17581_14197# a_17931_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2803 a_22259_14735# a_21813_14735# a_22163_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2804 tdc0.w_ring_int_norsz[9] net39 a_12913_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2806 VGND a_24335_5461# a_24293_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2808 VGND _196_ _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2809 VPWR a_25731_14191# a_25899_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2810 a_11655_6397# a_10957_6031# a_11398_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2812 a_22254_13759# a_22086_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2813 a_11955_16745# a_11509_16373# a_11859_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2814 a_25593_10927# _083_ a_25677_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2815 a_18781_10927# tdc0.w_ring_buf[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2816 a_29361_8207# tdc1.w_ring_buf[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2817 a_27038_11989# a_26870_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2819 VPWR a_4595_6005# a_4582_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2820 tdc0.w_ring_norsz[16] net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2821 tdc0.w_ring_norsz[20] net24 a_22653_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2822 _027_ _170_ a_11533_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2823 a_19327_16189# a_18703_15823# a_19219_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2824 a_15444_13647# _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2825 _025_ _167_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2826 tdc0.w_ring_int_norsz[15] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2827 _086_ a_9503_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2828 tdc0.r_dly_store_ring[13] a_15135_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2829 a_23776_13481# a_23377_13109# a_23650_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2830 a_29020_9129# a_28621_8757# a_28894_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2831 a_10881_16073# _143_ a_10799_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2833 a_22729_13481# a_21739_13109# a_22603_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2834 a_6813_6953# a_5823_6581# a_6687_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2836 net23 a_13735_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2837 a_7705_4765# a_7661_4373# a_7539_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2838 a_4420_4943# a_3505_4943# a_4073_5185# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2839 a_12153_7669# a_11987_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2840 VPWR tdc0.r_ring_ctr[9] a_16127_14557# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X2841 VGND _181_ a_5720_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2842 VGND _065_ a_19425_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X2843 a_14655_8751# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2844 tdc1.w_ring_norsz[22] net19 a_17317_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2846 a_5907_5487# tdc1.r_ring_ctr[14] _185_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.27 ps=2.54 w=1 l=0.15
X2848 tdc0.w_ring_buf[27] a_25971_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2849 VGND net28 a_7295_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2850 VPWR tdc0.w_ring_norsz[19] a_23303_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2851 a_8086_15645# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
R38 net47 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2854 VGND a_27222_9813# a_27180_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2855 uo_out[6] a_11792_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2856 a_15078_15823# _040_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2859 tdc0.r_dly_store_ring[18] a_27463_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2860 a_19784_15823# a_18703_15823# a_19437_16065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2861 a_5510_11583# a_5342_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2862 tdc0.w_ring_int_norsz[16] tdc0.w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2863 tdc1.r_dly_store_ring[6] a_18171_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2864 tdc0.r_dly_store_ring[18] a_27463_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2865 a_20924_4943# a_20525_4943# a_20798_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2867 a_16827_15823# a_16477_15823# a_16732_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2868 a_25401_13103# a_24867_13109# a_25306_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2869 a_22373_4399# _164_ _167_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2870 a_13441_6581# a_13275_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2871 a_13714_14191# a_13275_14197# a_13629_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2872 a_21665_7663# a_21327_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2873 VPWR a_24738_8725# a_24665_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2874 a_15051_12015# a_14269_12021# a_14967_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2875 a_14623_3615# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2876 a_11491_2767# a_10975_2767# a_11396_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2877 VPWR a_12353_14977# a_12243_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2878 a_18003_8573# a_17305_8207# a_17746_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2879 VGND a_5291_9813# a_5249_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2880 _172_ _169_ a_10245_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2884 VPWR _196_ _053_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2885 VPWR _070_ a_18243_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2886 VGND a_29871_8573# a_30039_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2887 a_4249_13103# _162_ _005_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2889 a_28331_12233# net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2892 tdc1.r_dly_store_ctr[15] a_6119_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2893 VGND net19 _058_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2894 a_27413_11305# a_26866_11049# a_27066_11204# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2895 _154_ a_15115_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2900 a_11873_12559# tdc0.r_dly_store_ring[22] a_11435_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2901 VGND _091_ a_26891_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2902 a_16297_14557# tdc0.r_ring_ctr[9] a_16209_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2903 tdc0.r_dly_store_ctr[8] a_14583_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2904 VGND _094_ a_21279_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2905 VPWR a_20947_6397# a_21115_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2906 a_5951_7485# a_5253_7119# a_5694_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2909 _080_ a_19631_8867# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2910 a_21718_9839# a_21445_9845# a_21633_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2911 a_24478_10927# a_24039_10933# a_24393_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2912 VPWR _180_ a_14644_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.195 ps=1.39 w=1 l=0.15
X2913 VPWR net29 a_9411_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2914 VPWR net29 a_11711_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2915 a_11233_11721# tdc0.r_dly_store_ring[6] a_11149_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2916 a_27379_12015# a_26597_12021# a_27295_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2917 a_25348_10633# _102_ a_25264_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2919 VPWR _095_ a_26127_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
R39 VPWR tdc0.g_ring3[26].stg01_53.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2920 VPWR tdc1.r_dly_store_ring[8] a_13637_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
R40 VGND net76 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2922 tdc1.w_ring_int_norsz[2] tdc1.w_ring_norsz[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2923 tdc1.w_ring_buf[25] a_28271_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2924 a_13897_10383# tdc0.r_dly_store_ctr[0] a_13551_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2925 a_9953_7369# tdc1.r_dly_store_ctr[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2926 VPWR tdc0.w_ring_norsz[25] a_17875_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2928 a_29319_8751# a_28455_8757# a_29062_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2929 VPWR tdc0.w_ring_norsz[27] a_20349_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2930 _143_ a_20503_15253# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2931 a_3392_8725# net26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2933 net39 a_17375_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2934 VPWR net33 a_17323_8759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2935 VPWR a_11763_8725# net30 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2936 a_9850_12015# a_9411_12021# a_9765_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2937 VPWR net32 a_16403_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2938 VGND a_23671_15287# net36 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2939 tdc0.w_ring_int_norsz[25] tdc0.w_ring_norsz[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2940 _091_ a_26431_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2942 VGND _012_ a_9690_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2943 VGND tdc0.w_dly_stop[5] a_3799_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2944 a_21912_6575# _113_ a_21743_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X2945 a_14542_12015# a_14103_12021# a_14457_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2946 VGND _046_ a_4025_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2947 VPWR a_17267_13103# a_17435_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2948 a_24665_8751# a_24131_8757# a_24570_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2949 VPWR a_16771_8751# _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2950 net33 a_17283_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2951 VPWR a_25474_13077# a_25401_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2952 a_22435_10357# a_22726_10657# a_22677_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2953 VGND a_17267_13103# a_17435_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2954 _140_ tdc0.r_ring_ctr[2] a_19715_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2955 VGND net17 tdc1.w_ring_norsz[18] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2957 a_15289_11247# tdc0.r_dly_store_ctr[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2958 a_13161_9071# tdc1.r_dly_store_ring[24] a_12815_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2959 tdc0.w_ring_buf[24] a_9135_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2960 VGND a_20966_5055# a_20924_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2961 VPWR tdc1.r_dly_store_ring[2] a_22351_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2962 a_4423_15101# a_3799_14735# a_4315_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2963 a_11045_4943# a_10055_4943# a_10919_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2964 tdc1.w_ring_norsz[17] net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2965 VGND _111_ a_21511_9447# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X2966 tdc1.r_dly_store_ctr[8] a_12835_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2967 VGND a_9963_8751# _077_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2968 a_7657_3855# a_6467_3855# a_7548_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2969 a_8102_7663# a_7663_7669# a_8017_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2970 a_11426_15599# _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X2971 tdc0.w_ring_norsz[15] tdc0.w_ring_norsz[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2972 VGND a_12835_5211# a_12793_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2973 a_10569_7093# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X2974 a_19142_14013# a_18869_13647# a_19057_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2977 VPWR tdc0.w_ring_norsz[20] a_17037_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2978 a_17392_15823# a_16311_15823# a_17045_16065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2979 a_9058_16189# a_8932_16091# a_8654_16075# VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2982 a_17739_7882# tdc1.w_ring_norsz[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2983 a_3668_12559# _005_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2984 uo_out[4] a_21912_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2985 VPWR tdc0.r_ring_ctr[12] a_3521_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2987 a_12609_9295# a_11619_9295# a_12483_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2988 a_10735_14013# a_9871_13647# a_10478_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2989 a_23569_6281# net65 tdc1.w_ring_int_norsz[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2990 VPWR tdc1.w_ring_int_norsz[14] a_12981_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2992 a_3686_9661# a_3247_9295# a_3601_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2993 VPWR tdc0.w_dly_stop[2] a_2787_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2995 _032_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2996 a_21223_5309# a_20525_4943# a_20966_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2997 VGND a_19867_4703# a_19801_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2998 a_23377_13109# a_23211_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2999 a_22381_14977# a_22163_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3000 a_24765_13897# _077_ a_24849_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3002 tdc1.w_ring_buf[9] a_27903_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3004 a_23726_9813# a_23558_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3005 VGND a_24351_4399# a_24519_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3006 a_17011_3855# a_16495_3855# a_16916_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3007 a_19713_8867# a_19439_9111# a_19631_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3008 tdc1.r_dly_store_ctr[5] a_13203_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3009 uo_out[6] a_11792_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X3010 tdc0.w_ring_buf[25] a_17875_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3011 a_8937_4943# tdc1.r_ring_ctr[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3012 tdc1.r_ring_ctr[4] a_17935_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X3014 a_19437_16065# a_19219_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3015 a_2769_7119# tdc1.r_ring_ctr[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3017 tdc0.r_dly_store_ring[19] a_24243_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3018 VPWR a_12539_9839# _072_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3019 _172_ tdc1.r_ring_ctr[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3020 a_10781_10633# tdc0.r_dly_store_ring[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3022 a_7557_13103# tdc0.r_ring_ctr[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3023 a_6559_8457# net60 a_6813_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3024 tdc0.r_dly_store_ring[19] a_24243_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3025 a_19389_4765# a_19345_4373# a_19223_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3026 a_21151_15823# a_20801_15823# a_21056_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3027 a_19034_10901# a_18866_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3028 VGND a_4588_7637# _623_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X3031 a_9849_8207# a_8859_8207# a_9723_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3032 VGND a_21886_9813# a_21844_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3033 a_17267_13103# a_16403_13109# a_17010_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3034 a_12805_12015# net21 tdc0.w_ring_norsz[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3036 a_18103_10205# tdc0.r_dly_store_ring[5] a_17740_10071# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X3037 a_3855_6031# a_3339_6031# a_3760_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3038 a_3854_8319# a_3686_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3039 a_17935_4703# a_17760_4777# a_18114_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3040 VPWR a_4073_6273# a_3963_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3041 a_21718_8751# a_21445_8757# a_21633_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3044 tdc0.w_ring_buf[1] a_19347_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3045 VGND net21 tdc0.w_ring_norsz[22] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3046 a_3963_5309# _061_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3047 a_8723_11636# tdc0.w_ring_norsz[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3048 a_27411_7093# tdc1.w_dly_stop[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3049 a_22257_9545# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X3050 a_24849_9839# a_25071_9813# a_24683_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3051 tdc0.w_ring_norsz[26] tdc0.w_ring_int_norsz[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3053 a_10310_14013# a_10037_13647# a_10225_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3054 VGND _107_ a_21743_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3055 _066_ _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3056 VPWR _196_ _054_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3057 net26 a_3115_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3058 a_10045_5487# tdc1.r_dly_store_ring[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3059 VPWR tdc1.w_ring_norsz[4] a_20083_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3060 a_24021_14735# a_23855_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3061 VPWR a_14703_12724# tdc0.w_ring_buf[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3062 VGND a_17751_3829# tdc1.r_ring_ctr[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3063 a_23075_10383# a_22855_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3064 VPWR a_5417_4917# _183_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3065 _139_ a_6027_9622# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3066 VGND _196_ _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3067 tdc0.r_ring_ctr[8] a_14899_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X3068 VPWR a_22695_5487# a_22863_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3069 a_17704_12559# a_17305_12559# a_17578_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3070 VGND tdc1.r_dly_store_ctr[10] a_20433_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X3071 a_25373_10159# _085_ a_25071_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3074 _095_ a_21279_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X3075 a_3871_7485# _063_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3076 tdc1.r_dly_store_ctr[8] a_12835_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3077 a_16247_6397# a_15465_6031# a_16163_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3078 a_24159_13103# a_23377_13109# a_24075_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
R41 VPWR tt_um_hpretl_tt06_tdc_v2_90.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3080 VGND a_18059_16375# net9 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3081 VGND _066_ a_21717_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X3082 a_8228_8041# a_7829_7669# a_8102_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3084 a_27790_5487# a_27517_5493# a_27705_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3085 a_21843_8041# a_21707_7881# a_21423_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3086 VGND _147_ _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3087 VGND _112_ a_20729_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3088 a_18869_10383# a_18703_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3090 a_16213_12809# tdc0.w_ring_norsz[1] a_16129_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3091 net22 a_19255_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3092 a_25505_12335# tdc0.r_dly_store_ctr[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X3093 a_7055_12925# a_6357_12559# a_6798_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3094 a_3812_9295# a_3413_9295# a_3686_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3096 a_20175_13103# _077_ a_20353_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3097 VGND net58 tdc0.w_ring_int_norsz[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3098 VPWR _109_ a_20883_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3099 VGND a_25071_10901# a_25029_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3100 a_18003_8573# a_17139_8207# a_17746_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3102 VGND a_24849_9839# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3105 VGND net21 tdc0.w_ring_norsz[31] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3106 VPWR _195_ _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3107 a_9006_7231# a_8838_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3108 VPWR tdc0.w_ring_norsz[12] a_19899_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3109 a_25857_14569# a_24867_14197# a_25731_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3111 VPWR tdc1.w_ring_int_norsz[6] a_16937_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3112 net29 a_9924_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3113 tdc1.w_ring_norsz[8] tdc1.w_ring_int_norsz[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3114 VGND _083_ a_10594_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3115 a_9006_7231# a_8838_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3117 a_7001_6031# a_6835_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3118 a_12333_14569# a_11343_14197# a_12207_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3119 VPWR a_14623_3615# a_14610_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3123 a_22719_10357# net35 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3124 tdc0.w_ring_norsz[3] tdc0.w_ring_norsz[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3126 VPWR a_21886_9813# a_21813_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3128 VGND a_25731_4221# a_25899_4123# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3129 VPWR tdc1.r_ring_ctr[12] a_5907_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.162 ps=1.33 w=1 l=0.15
X3130 VPWR a_4328_7119# a_4503_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3131 a_21423_7895# a_21707_7881# a_21642_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3132 VPWR a_17045_16065# a_16935_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3133 tdc1.w_ring_buf[16] a_7111_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3134 VPWR _068_ a_10087_10411# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3136 tdc0.w_ring_int_norsz[5] net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3138 a_21369_16065# a_21151_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3139 a_22811_3615# a_22636_3689# a_22990_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3140 a_5951_7485# a_5087_7119# a_5694_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3141 VPWR _012_ a_9690_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3142 VGND _157_ a_6191_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3143 a_19032_4765# _024_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3144 VPWR _190_ a_14351_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3145 VGND tdc1.r_ring_ctr[0] a_13797_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3146 a_3108_10927# a_2894_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X3147 VPWR a_29487_8725# a_29403_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3149 a_3789_13897# _158_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3151 a_19505_10205# tdc0.r_dly_store_ring[25] a_19433_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3153 a_8654_14191# a_8215_14197# a_8569_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3154 VGND a_2519_7369# _022_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X3155 a_3870_10749# a_3431_10383# a_3785_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3156 a_14073_4765# tdc1.r_ring_ctr[9] a_14001_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3160 a_14644_5487# _178_ a_14553_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.153 ps=1.3 w=1 l=0.15
X3161 a_24021_14735# a_23855_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3162 VGND net3 a_9411_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3164 a_11115_4007# _168_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X3166 uo_out[5] a_15504_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3167 a_26891_12559# _067_ a_27069_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3169 a_29733_7983# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X3170 VGND tdc0.w_dly_stop[2] a_2787_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3171 VGND tdc0.w_ring_norsz[5] a_16219_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3172 a_23657_5487# tdc1.r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3173 a_3505_11471# tdc0.r_ring_ctr[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3174 a_27036_7637# net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3175 tdc1.w_ring_int_norsz[18] net63 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3177 a_17949_6575# tdc1.w_ring_norsz[21] a_17865_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3178 a_24754_7663# a_24481_7669# a_24669_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3179 _069_ a_10975_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3180 a_15168_4943# _018_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3181 a_15487_10633# _115_ a_15391_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3182 a_3760_4943# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3183 tdc0.w_ring_buf[5] a_16219_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3184 a_20713_4943# tdc1.r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3185 tdc1.w_ring_int_norsz[8] tdc1.w_ring_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3187 a_20727_14735# tdc0.r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3188 VPWR _196_ _049_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3189 a_15005_7119# a_14839_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3190 a_23285_9845# a_23119_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R42 tdc0.g_ring3[28].stg01_55.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3191 VPWR a_14983_14165# net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3192 VGND a_12863_5719# tdc1.r_dly_store_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3193 VPWR net25 a_9953_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3194 a_19867_4703# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3195 VGND a_3854_9407# a_3812_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3196 VPWR net36 a_26615_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3198 a_9740_3855# tdc1.r_ring_ctr[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3200 tdc0.w_ring_int_norsz[10] tdc0.w_ring_norsz[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3201 VPWR tdc1.r_ring_ctr[12] a_5507_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X3202 a_21511_9447# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X3203 VGND a_30254_7895# a_30203_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3204 a_2807_11169# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3205 a_20801_15823# a_20635_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3206 a_9206_6397# a_8767_6031# a_9121_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3207 VPWR a_21716_15823# a_21891_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3209 VPWR a_12007_13077# a_11923_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3210 a_21813_9839# a_21279_9845# a_21718_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3211 _138_ a_10977_9955# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3212 a_25692_8207# _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X3213 a_20617_6575# tdc1.r_dly_store_ctr[12] a_20533_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3214 a_9282_13077# a_9114_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3215 tdc1.w_ring_norsz[12] tdc1.w_ring_norsz[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3216 a_29955_8983# tdc1.r_dly_store_ring[25] a_30101_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X3217 tdc1.r_dly_store_ring[30] a_9799_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3220 a_25677_10927# tdc0.r_dly_store_ring[3] a_25593_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3221 a_7461_10927# tdc0.w_ring_norsz[23] a_7377_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3222 a_25214_5487# a_24941_5493# a_25129_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3223 a_25857_13481# a_24867_13109# a_25731_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3224 VPWR tdc1.w_ring_int_norsz[20] a_23377_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3225 VPWR tdc1.w_ring_norsz[22] a_11885_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3226 a_4111_9661# a_3413_9295# a_3854_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3227 _113_ a_20729_9955# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3228 VGND tdc0.w_dly_stop[3] a_2879_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3229 VGND _075_ a_20613_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X3230 a_25306_4221# a_25033_3855# a_25221_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3231 VPWR a_14967_12015# a_15135_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3232 a_26513_13103# tdc0.r_dly_store_ring[10] a_26431_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3233 VGND net15 a_8399_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3234 a_11609_7663# net16 tdc1.w_ring_norsz[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3235 tdc0.w_ring_buf[22] a_10975_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3237 a_11763_8725# net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X3238 a_6907_14191# _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3239 VGND a_14967_12015# a_15135_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3240 VPWR a_21886_8725# a_21813_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R43 VPWR tt_um_hpretl_tt06_tdc_v2_84.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3241 a_4943_9622# a_4761_9622# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3242 a_16845_2767# a_16679_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3243 a_10699_10633# _066_ a_10781_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3244 a_23565_13103# tdc0.w_ring_buf[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3247 a_21445_7369# tdc1.r_dly_store_ctr[2] a_21361_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3248 _019_ _181_ a_6541_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X3249 a_20327_3615# _048_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3250 VGND net27 a_4903_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3251 VPWR a_18671_14495# a_18658_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3252 _018_ a_14644_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3254 _088_ a_20175_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X3255 a_7091_4221# a_6467_3855# a_6983_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3256 a_21976_3677# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3257 tdc0.w_ring_int_norsz[17] tdc0.w_ring_norsz[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3259 VGND a_11087_5211# a_11045_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3260 a_23469_5493# a_23303_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3261 a_11230_6397# a_10791_6031# a_11145_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3262 VGND tdc0.r_ring_ctr[3] a_20359_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X3264 VPWR a_9963_8751# _077_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3265 a_12231_2741# _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3266 a_4295_10749# a_3431_10383# a_4038_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3267 a_24393_10927# tdc0.w_ring_buf[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3268 VGND net22 _042_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3269 a_22252_15645# _009_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3270 VPWR a_27491_5108# tdc1.w_dly_stop[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3271 tdc0.w_ring_int_norsz[10] net41 a_18249_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3272 tdc1.r_dly_store_ring[27] a_30039_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3273 a_28047_12247# a_28338_12137# a_28289_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3275 VGND net12 tdc0.w_ring_int_norsz[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3276 VGND a_12651_9563# a_12609_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3277 VPWR tdc1.r_ring_ctr[10] a_15481_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3278 tdc0.r_dly_store_ctr[11] a_22679_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3279 VGND _065_ a_19899_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3280 VGND tdc0.r_ring_ctr[7] a_9253_14763# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3281 a_3686_8573# a_3413_8207# a_3601_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3282 VPWR a_20303_5487# a_20471_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3283 a_20303_5487# a_19605_5493# a_20046_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3284 VGND a_9707_13077# a_9665_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3285 a_26149_6575# tdc1.w_ring_norsz[12] a_26065_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3286 a_6078_10749# a_5639_10383# a_5993_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3287 tdc1.w_ring_norsz[20] tdc1.w_ring_norsz[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3288 VPWR tdc0.w_ring_norsz[17] a_15483_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3289 a_17305_12559# a_17139_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3290 a_12621_3855# _175_ _180_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3291 VPWR net20 _045_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3292 a_18029_13647# a_17475_13621# a_17682_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3293 a_11739_6397# a_10957_6031# a_11655_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3294 VGND net25 a_14011_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3295 VPWR net24 a_13735_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3296 a_17611_13647# a_17482_13921# a_17191_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3298 tdc1.w_ring_norsz[2] net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3299 VPWR _075_ a_12529_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3300 a_7699_6397# a_6835_6031# a_7442_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3301 VGND a_17083_9839# a_17251_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3302 tdc0.w_ring_norsz[12] tdc0.w_ring_norsz[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3303 VGND _064_ a_15159_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3304 VGND a_24519_4373# a_24477_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3305 a_9332_6031# a_8933_6031# a_9206_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3307 VPWR a_10699_14735# _152_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3308 VGND a_14710_11989# a_14668_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3309 a_10478_13759# a_10310_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3310 VPWR _069_ a_10045_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3311 a_22728_14735# a_21647_14735# a_22381_14977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3313 VGND a_9891_8475# a_9849_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3314 a_25079_8751# a_24297_8757# a_24995_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3315 a_11505_11471# tdc0.r_dly_store_ring[14] a_11067_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3316 VGND _075_ a_26777_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3317 VGND a_10735_14013# a_10903_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3318 VPWR tdc0.r_ring_ctr[11] a_16127_14557# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X3319 a_20603_13621# net32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3320 a_4420_4943# a_3339_4943# a_4073_5185# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3322 _085_ tdc1.r_dly_store_ring[1] a_24674_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X3323 _191_ a_10699_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X3325 a_21813_8751# a_21279_8757# a_21718_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3326 a_4503_12533# a_4328_12559# a_4682_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3327 VGND a_19310_10495# a_19268_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3328 tdc0.r_dly_store_ring[12] a_20931_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3329 VPWR a_15261_11445# _114_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3330 a_19479_7983# a_19425_7895# a_19379_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X3331 _174_ a_10607_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3332 a_8017_7663# tdc1.w_ring_buf[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3333 VGND tdc1.w_ring_norsz[16] tdc1.w_ring_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3336 a_20798_5309# a_20525_4943# a_20713_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3338 VPWR _113_ a_21912_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X3339 VPWR a_9643_12724# tdc0.w_ring_buf[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3341 tdc0.w_ring_norsz[21] tdc0.w_ring_norsz[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3345 VPWR tdc1.r_dly_store_ring[31] a_10787_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3346 a_12851_7663# a_12153_7669# a_12594_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3347 a_20230_12671# a_20062_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3348 VGND _084_ a_20451_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3349 a_11149_11721# _086_ a_11067_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3350 a_17578_8573# a_17139_8207# a_17493_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3352 VPWR a_14155_4917# _179_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
R44 VPWR tdc0.g_ring3[22].stg01_49.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3353 a_7745_10927# net21 tdc0.w_ring_norsz[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3354 _067_ a_11987_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3355 a_24209_14735# tdc0.r_ring_ctr[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3356 a_16845_2767# a_16679_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3357 a_8912_15599# tdc0.r_ring_ctr[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3358 VPWR a_22438_5461# a_22365_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3359 net12 a_19255_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3360 a_10493_13423# tdc0.r_dly_store_ring[30] a_10147_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3361 tdc1.w_ring_int_norsz[16] net61 a_5277_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3362 _071_ _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3364 VPWR a_4111_8573# a_4279_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3365 VGND a_19034_6549# a_18992_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3366 VGND tdc0.r_dly_store_ring[28] a_20341_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X3367 a_11356_6031# a_10957_6031# a_11230_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3368 a_4038_10495# a_3870_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3369 VGND a_12599_16671# a_12533_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3370 net15 a_9103_4659# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3372 net36 a_23671_15287# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3373 a_13599_5853# a_13379_5865# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3374 a_11713_6691# _127_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3375 a_24029_12559# tdc0.r_dly_store_ring[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3376 VGND a_25899_14165# a_25857_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3377 VPWR a_29119_7637# a_29035_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3378 a_26969_9839# tdc1.w_ring_buf[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3380 tdc0.w_ring_buf[20] a_22843_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3381 a_2601_7369# _184_ a_2519_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3382 VPWR a_4038_10495# a_3965_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3383 a_8639_3689# a_8123_3317# a_8544_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3385 VGND a_26420_11721# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3386 a_15023_13103# _077_ a_15105_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3388 a_12243_15101# a_11619_14735# a_12135_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3389 a_15283_8457# _065_ a_15701_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3391 a_5526_7485# a_5087_7119# a_5441_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3392 a_24021_12021# a_23855_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3393 a_26617_8751# tdc1.w_ring_int_norsz[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3395 VPWR a_24922_7637# a_24849_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3400 VPWR _117_ a_15333_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3401 VPWR _104_ a_25616_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X3402 VPWR _086_ a_6241_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X3403 VGND _195_ _038_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3405 a_13173_12809# net38 tdc0.w_ring_int_norsz[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3407 a_29446_8573# a_29173_8207# a_29361_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3408 a_13161_4777# a_12171_4405# a_13035_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3409 a_25327_12015# _077_ a_25505_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3410 a_20338_11837# a_20065_11471# a_20253_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3411 VGND a_9374_6143# a_9332_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
R45 tdc1.g_ring3[17].stg01_62.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3412 a_28526_9839# a_28253_9845# a_28441_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3413 a_25033_14197# a_24867_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3414 VGND a_16463_12533# net38 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3416 a_5468_11471# a_5069_11471# a_5342_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3417 VPWR a_22912_15657# a_23087_15583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3418 a_24849_13897# tdc0.r_dly_store_ctr[11] a_24765_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3419 VGND tdc0.w_ring_norsz[28] tdc0.w_ring_int_norsz[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3421 a_3601_9295# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3422 a_18866_6575# a_18427_6581# a_18781_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3423 VGND net36 a_26615_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3424 VPWR a_25382_5461# a_25309_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3425 VGND tdc1.w_ring_buf[18] a_22261_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3427 a_21270_12809# _083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3428 VGND tdc0.w_ring_norsz[26] tdc0.w_ring_norsz[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3429 a_12437_6031# _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X3430 a_15023_13103# _077_ a_15105_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3431 VPWR a_25474_3967# a_25401_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3432 a_4503_7093# a_4328_7119# a_4682_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3433 a_22365_5487# a_21831_5493# a_22270_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3436 _193_ a_14197_10389# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3438 VGND a_30856_7895# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3440 a_17704_8207# a_17305_8207# a_17578_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3441 a_11705_8457# tdc1.w_ring_norsz[24] a_11621_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3442 VPWR a_9503_9295# _086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3443 a_22389_12809# tdc0.w_ring_norsz[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3445 VGND tdc1.w_ring_int_norsz[15] tdc1.w_ring_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3446 VPWR tdc1.r_dly_store_ring[22] a_12437_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3447 a_19034_6549# a_18866_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3450 a_17853_5865# a_16863_5493# a_17727_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3451 VPWR net31 a_21279_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3453 VPWR a_22381_14977# a_22271_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3454 tdc0.w_ring_buf[27] a_25971_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3455 a_19327_16189# _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3456 a_8937_4943# tdc1.r_ring_ctr[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3457 VGND a_11398_6143# a_11356_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3458 VGND net15 tdc1.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3461 VPWR net19 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3462 tdc0.r_dly_store_ring[10] a_25899_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3464 a_15569_14511# _157_ a_15351_14423# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3465 a_15263_4943# a_14747_4943# a_15168_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3466 tdc0.r_dly_store_ring[10] a_25899_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3467 a_6907_14191# a_6283_14197# a_6799_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3468 a_9723_8573# a_8859_8207# a_9466_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3469 _069_ a_10975_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3470 tdc0.r_dly_store_ring[4] a_22311_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3471 _115_ a_15207_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3473 a_15005_7119# a_14839_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3474 VPWR a_16209_8751# a_16309_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X3475 VPWR a_3854_8319# a_3781_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3476 a_6241_9622# tdc0.r_dly_store_ring[7] a_6027_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X3477 a_5652_7119# a_5253_7119# a_5526_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3478 a_25071_9813# _085_ a_25373_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3479 a_20152_3689# a_19237_3317# a_19805_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3481 VPWR tdc1.r_dly_store_ctr[0] a_13887_8359# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3482 tdc1.r_ring_ctr[5] a_12231_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3484 a_15465_6031# a_15299_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3486 a_15399_4399# _177_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3488 VPWR a_20327_3615# a_20314_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3489 a_22347_15657# a_21831_15285# a_22252_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3491 tdc0.r_ring_ctr[13] a_7539_14495# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3492 VGND a_27491_5108# tdc1.w_dly_stop[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3493 VPWR _065_ a_18243_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X3495 _011_ _146_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3496 VPWR a_7867_6299# a_7783_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3497 tdc1.r_dly_store_ring[23] a_9891_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3499 a_20165_14735# tdc0.r_ring_ctr[0] a_20083_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X3500 a_14116_13647# a_13717_13647# a_13990_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3501 a_15256_10535# _116_ a_15487_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3502 a_27057_12809# tdc0.r_dly_store_ring[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3503 VGND _083_ a_20889_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X3504 tdc1.w_ring_int_norsz[2] net40 a_23033_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3506 VGND net30 a_15299_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3507 tdc1.w_ring_int_norsz[14] net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3508 a_17543_9661# a_16679_9295# a_17286_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3511 VGND net37 a_13551_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3512 VPWR a_12231_2741# a_12218_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3513 a_16129_12809# tdc0.w_ring_int_norsz[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3514 a_7442_6143# a_7274_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3515 VGND tdc0.w_ring_int_norsz[19] tdc0.w_ring_norsz[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3517 VPWR a_9263_7485# a_9431_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3519 VGND a_18751_8359# _129_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X3520 VGND net4 a_16587_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3521 a_25401_4221# a_24867_3855# a_25306_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3522 tdc1.w_ring_int_norsz[29] net74 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3525 a_13379_5865# a_13243_5705# a_12959_5719# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3527 uo_out[1] a_24849_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3528 tdc0.w_ring_norsz[11] net22 a_21457_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3530 VPWR a_7810_13077# a_7737_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3531 a_14723_4765# tdc1.r_ring_ctr[10] a_14627_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X3533 a_18992_6953# a_18593_6581# a_18866_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3535 tdc1.w_ring_int_norsz[8] net38 a_11073_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3536 a_11582_13077# a_11414_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3537 _037_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3539 tdc0.r_dly_store_ctr[9] a_19735_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3540 _177_ a_13919_4512# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3541 a_4111_9661# a_3247_9295# a_3854_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3542 a_23102_10749# a_22855_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3543 VPWR a_20966_5055# a_20893_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3545 a_4025_12559# a_3981_12801# a_3859_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3546 VPWR a_19735_13915# a_19651_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3547 a_12447_13103# _077_ a_12529_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3548 VPWR net34 a_24315_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3549 VPWR a_17760_4777# a_17935_4703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3550 VGND net40 tdc1.w_ring_int_norsz[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3551 VPWR a_6980_4917# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3552 VGND a_17746_8319# a_17704_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3553 a_12065_10383# tdc0.w_ring_buf[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3554 tdc1.w_ring_int_norsz[0] net77 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3555 a_9313_3689# a_8123_3317# a_9204_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3556 a_24849_9839# _090_ a_24765_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3557 a_16127_14557# tdc0.r_ring_ctr[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X3558 VGND _156_ a_14921_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3559 a_23910_5461# a_23742_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3560 a_22227_9839# a_21445_9845# a_22143_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3561 _093_ a_25327_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X3562 VPWR a_12403_8970# tdc1.w_ring_buf[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3563 tdc0.w_ring_buf[28] a_18151_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3564 a_3781_8573# a_3247_8207# a_3686_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3565 VPWR a_15719_10357# net25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3566 a_5989_12015# tdc0.w_ring_norsz[0] a_5905_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3567 tdc1.r_dly_store_ring[28] a_28383_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3568 a_4824_10217# a_4425_9845# a_4698_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3570 VPWR a_12851_7663# a_13019_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3571 a_17305_12559# a_17139_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3572 a_20341_13103# tdc0.r_dly_store_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3573 a_8653_10217# a_7663_9845# a_8527_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3574 VPWR a_15757_13889# a_15647_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3575 VGND a_24738_8725# a_24696_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3577 VPWR tdc1.r_ring_ctr[9] a_14951_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X3579 VGND a_5694_7231# a_5652_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3580 VGND a_25348_10633# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3581 VGND _195_ _034_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3582 VPWR a_19291_6575# a_19459_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3583 VGND tdc1.w_ring_int_norsz[26] tdc1.w_ring_norsz[26] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3584 tdc1.r_dly_store_ring[2] a_22311_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3585 tdc1.r_dly_store_ring[16] a_8327_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3586 net2 a_855_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3587 VPWR a_19459_10901# a_19375_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3590 a_22289_3285# a_22071_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3591 _151_ a_10239_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3592 a_9379_3615# _054_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3593 tdc1.r_ring_ctr[1] a_22811_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X3594 a_7897_7284# tdc1.w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3595 VPWR tdc1.r_ring_ctr[0] _016_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3596 VPWR a_3799_13103# net24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3597 a_6997_7663# net16 tdc1.w_ring_norsz[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3598 a_20603_13621# net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3599 _077_ a_9963_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3600 VPWR net2 a_3247_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3601 a_20763_11837# a_20065_11471# a_20506_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3602 VPWR a_29614_8319# a_29541_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3603 _086_ a_9503_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3604 a_9849_10159# tdc0.r_dly_store_ctr[7] a_9411_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
R46 VPWR tdc0.g_ring3[27].stg01_54.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3605 VGND tdc0.r_ring_ctr[9] a_15769_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X3606 VPWR tdc0.r_ring_ctr[0] a_20727_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3607 VGND a_3255_11721# _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X3608 a_13809_15823# a_13643_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3609 a_20157_7663# a_19991_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X3610 VPWR a_28694_9813# a_28621_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3611 a_18884_8207# _081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X3612 VPWR ui_in[5] a_15575_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3613 VPWR a_21912_6575# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3614 a_13809_6575# a_13275_6581# a_13714_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3615 a_11509_14197# a_11343_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3617 tdc1.w_ring_buf[9] a_27903_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3618 VPWR tdc0.w_ring_norsz[14] a_7745_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3621 a_6559_8457# tdc1.w_ring_int_norsz[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3622 a_20893_5309# a_20359_4943# a_20798_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3623 VGND net10 a_20635_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3626 a_4423_15101# _044_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3627 a_9577_9839# tdc0.r_dly_store_ring[15] a_9493_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3628 a_22926_10357# a_22719_10357# a_23102_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3629 tdc0.w_ring_norsz[5] tdc0.w_ring_norsz[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3632 VPWR a_17751_3829# a_17738_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3633 VGND tdc0.r_ring_ctr[0] a_18029_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3634 VPWR a_23080_14165# net35 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3635 tdc0.w_ring_int_norsz[3] net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3636 a_15657_3855# tdc1.r_ring_ctr[8] _176_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3637 _083_ a_20083_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3638 tdc1.r_ring_ctr[0] a_20327_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3639 a_7377_10927# net20 tdc0.w_ring_norsz[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3640 VPWR net35 a_26431_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
R47 net45 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3641 _072_ a_12539_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3642 VPWR tdc1.w_ring_buf[0] a_15023_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3643 a_5993_10383# tdc0.w_ring_buf[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3644 a_11329_13103# tdc0.w_ring_buf[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3646 a_22063_8029# a_21843_8041# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3647 a_8933_6031# a_8767_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3650 a_26794_11293# a_26479_11159# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3651 a_19793_5487# tdc1.r_ring_ctr[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3652 a_9871_7369# _076_ a_9953_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3653 _173_ a_9811_4737# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3654 VGND a_4111_8573# a_4279_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3655 a_17882_10205# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X3656 VGND net51 tdc0.w_ring_int_norsz[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3659 VGND a_5602_13759# a_5560_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3660 _016_ tdc1.r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3661 a_15351_14423# _157_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X3663 a_12935_7663# a_12153_7669# a_12851_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3664 a_18658_14191# a_17581_14197# a_18496_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3665 a_4533_14977# a_4315_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3667 a_22227_8751# a_21445_8757# a_22143_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3668 VPWR a_12587_8372# tdc1.w_ring_buf[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3669 a_21743_6895# _108_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3670 tdc1.w_ring_norsz[10] net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3671 VGND a_24995_8751# a_25163_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3672 a_14342_10901# a_14174_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3673 VPWR a_12483_9661# a_12651_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3674 VPWR net35 a_24867_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3675 a_11859_16745# a_11509_16373# a_11764_16733# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3676 VPWR a_9891_8475# a_9807_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3677 a_6980_4917# tdc1.w_ring_buf[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3678 _059_ net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3680 VPWR tdc0.r_ring_ctr[10] a_16677_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3682 _042_ net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3683 tdc1.w_ring_norsz[1] tdc1.w_ring_int_norsz[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3684 a_10512_9545# _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3685 VPWR a_5043_8372# tdc1.w_ring_buf[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3686 VGND tdc1.w_ring_norsz[4] a_20083_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3687 a_11145_6031# tdc1.w_ring_buf[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3688 a_4425_8757# a_4259_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3689 a_11885_10927# net38 tdc0.w_ring_int_norsz[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3690 a_23841_4399# tdc1.r_ring_ctr[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3691 a_29541_8573# a_29007_8207# a_29446_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3692 tdc0.w_ring_int_norsz[27] net54 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3693 a_24213_6281# tdc1.r_dly_store_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3694 a_5805_10383# a_5639_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3695 VPWR tdc0.w_ring_norsz[0] a_5271_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3696 VPWR a_24167_5487# a_24335_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3697 a_28951_9839# a_28253_9845# a_28694_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3698 a_4219_13621# tdc0.r_ring_ctr[12] a_4617_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X3699 a_24167_5487# a_23469_5493# a_23910_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3700 a_22636_3689# a_21555_3317# a_22289_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3701 VGND net33 a_19899_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3703 a_28621_9839# a_28087_9845# a_28526_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3704 a_13901_10933# a_13735_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3705 tdc0.r_dly_store_ring[24] a_10443_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3706 VGND a_20327_3615# tdc1.r_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3707 a_5943_14013# a_5161_13647# a_5859_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3708 a_8803_12015# a_8105_12021# a_8546_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3709 net20 a_3399_12275# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3710 a_4437_12559# a_3247_12559# a_4328_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3711 a_25221_13103# tdc0.w_ring_buf[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3712 a_29077_10217# a_28087_9845# a_28951_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3714 a_10957_6031# a_10791_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3715 tdc0.r_dly_store_ctr[12] a_7223_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3716 VPWR a_17711_9563# a_17627_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3717 a_10487_4765# _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X3718 VPWR a_14059_8983# _076_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3719 a_16732_15823# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3722 VPWR net26 a_6835_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3723 VPWR tdc1.w_ring_norsz[6] a_16577_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3725 VGND net22 tdc0.w_ring_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3726 VPWR tdc0.w_ring_norsz[13] a_13173_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3727 a_8546_11989# a_8378_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3728 VGND a_2840_12533# _622_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X3729 VPWR a_20230_12671# a_20157_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3730 a_9298_8573# a_8859_8207# a_9213_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3731 a_15828_4943# a_14747_4943# a_15481_5185# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3732 a_12610_4399# a_12337_4405# a_12525_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3733 VGND net30 a_10791_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3734 a_10124_9269# _139_ a_10594_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3735 VPWR _070_ a_18335_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3738 _152_ a_10699_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X3739 a_10689_4765# _168_ a_10583_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X3740 _108_ a_20451_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X3741 a_3855_6031# a_3505_6031# a_3760_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3742 a_8017_9839# tdc0.w_ring_buf[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3743 a_8378_12015# a_8105_12021# a_8293_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3744 a_9190_5055# a_9022_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3746 VPWR tdc1.w_ring_norsz[29] a_15023_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3749 VPWR a_20603_13621# a_20610_13921# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3750 a_30389_9071# _072_ a_29955_8983# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3751 a_19605_5493# a_19439_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3752 VPWR tdc1.w_ring_norsz[9] a_27903_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3753 a_3965_14735# a_3799_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3754 a_19291_6575# a_18427_6581# a_19034_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3755 a_27793_8751# tdc1.w_ring_norsz[10] a_27709_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3756 VGND a_10919_5309# a_11087_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3757 a_20506_11583# a_20338_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3760 VGND _067_ a_24293_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3762 a_7723_3829# a_7548_3855# a_7902_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3763 a_27222_9813# a_27054_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3764 VGND _047_ a_2525_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X3765 VGND net27 a_3431_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3766 net20 a_3399_12275# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3768 tdc1.w_ring_norsz[22] tdc1.w_ring_int_norsz[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3769 VGND net23 tdc0.w_ring_norsz[21] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3770 VGND _070_ a_18776_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3772 a_12424_16745# a_11509_16373# a_12077_16341# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3773 a_15115_14735# tdc0.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3775 a_17922_4399# a_16845_4405# a_17760_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3776 a_10359_10927# a_9577_10933# a_10275_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3778 a_19142_10749# a_18869_10383# a_19057_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3779 a_6630_9839# a_6357_9845# a_6545_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3780 VPWR tdc1.r_ring_ctr[7] a_9836_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X3781 VGND tdc1.w_ring_norsz[2] tdc1.w_ring_int_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3782 a_3861_13647# tdc0.r_ring_ctr[13] a_3789_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0683 ps=0.86 w=0.65 l=0.15
X3783 a_17493_8207# tdc1.w_ring_buf[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3785 VPWR net12 a_27535_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3786 VGND a_17935_2741# a_17869_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3787 a_20959_13647# a_20739_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3788 tdc1.r_dly_store_ring[20] a_25807_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3789 _189_ a_13553_8867# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3790 uo_out[4] a_21912_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X3791 uo_out[5] a_15504_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X3792 VGND a_26420_11721# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3794 a_22439_3855# a_22089_3855# a_22344_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3795 a_7551_4399# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3796 a_14159_15823# a_13643_15823# a_14064_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3797 VPWR _080_ a_18877_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X3798 a_8113_11721# net38 tdc0.w_ring_int_norsz[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3799 VGND a_7907_15583# a_7841_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3800 VPWR a_9647_14709# _158_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X3801 a_12809_14735# a_11619_14735# a_12700_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3803 a_17457_2767# a_17413_3009# a_17291_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3805 a_17217_5487# tdc1.r_ring_ctr[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3806 a_8654_16075# a_8932_16091# a_8888_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3807 _064_ a_16587_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3809 a_20947_6397# a_20249_6031# a_20690_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3810 a_29587_7895# tdc1.r_dly_store_ring[11] a_29733_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3811 VPWR net36 a_27351_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3812 a_12426_7663# a_11987_7669# a_12341_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3813 a_24485_8751# tdc1.w_ring_buf[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3814 a_17083_9839# a_16219_9845# a_16826_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3815 VGND tdc0.w_ring_norsz[25] tdc0.w_ring_norsz[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3816 VPWR a_13450_5764# a_13379_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3817 a_11950_14165# a_11782_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3818 a_5441_7119# tdc1.r_ring_ctr[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3819 a_14377_16065# a_14159_15823# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3820 uo_out[7] a_10124_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3823 a_7829_9845# a_7663_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3825 a_25306_14191# a_25033_14197# a_25221_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3826 VPWR a_9371_4007# _029_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X3827 VGND tdc1.r_dly_store_ctr[11] a_18777_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X3829 VGND a_10975_8751# _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3830 _038_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3831 VPWR tdc1.w_ring_norsz[14] a_12539_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3832 VPWR a_12139_4007# _168_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3833 a_13620_9269# _083_ a_14008_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3834 VGND _066_ a_10493_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3835 a_9424_8207# a_9025_8207# a_9298_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3836 VPWR _068_ a_12897_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3837 VPWR a_7223_12827# a_7139_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3838 a_25263_7663# a_24481_7669# a_25179_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3839 VGND a_12483_9661# a_12651_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3842 a_23293_6575# net17 tdc1.w_ring_norsz[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3843 VPWR a_3247_13647# net37 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3844 VGND a_8183_4703# tdc1.r_ring_ctr[12] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3845 a_3963_6397# a_3339_6031# a_3855_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
R48 VGND net63 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3847 a_23087_15583# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3848 tdc1.r_ring_ctr[13] a_4595_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3849 a_21270_12809# _088_ a_21178_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X3852 a_27529_7663# tdc1.w_ring_norsz[27] a_27445_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R49 VPWR tdc0.g_ring3[20].stg01_47.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3854 a_6262_6575# a_5989_6581# a_6177_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3855 a_23818_13077# a_23650_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3856 a_3965_14735# a_3799_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3858 net10 a_14983_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3859 _162_ tdc0.r_ring_ctr[12] a_3861_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.119 ps=1.01 w=0.65 l=0.15
X3860 VPWR a_24462_14847# a_24389_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3862 VGND tdc1.w_ring_int_norsz[3] tdc1.w_ring_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3865 a_16463_12533# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X3867 tdc0.r_dly_store_ring[12] a_20931_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3869 a_19057_13647# tdc0.r_ring_ctr[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3870 VPWR net26 a_5823_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3871 a_15446_7231# a_15278_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3872 tdc1.w_ring_buf[2] a_21003_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3874 VPWR a_5043_10548# tdc0.w_ring_buf[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3876 VPWR a_14724_15823# a_14899_15797# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
R50 VPWR tt_um_hpretl_tt06_tdc_v2_92.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3878 a_14385_8457# tdc1.w_ring_norsz[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3879 a_14909_8751# a_15159_8725# _071_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3881 a_15446_7231# a_15278_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3883 VPWR tdc1.w_ring_norsz[26] a_27443_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3884 a_22653_12015# tdc0.w_ring_norsz[18] a_22569_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3885 tdc1.w_ring_norsz[0] tdc1.w_ring_norsz[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3886 VGND a_5935_11739# a_5893_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3887 a_25493_12015# tdc0.r_dly_store_ring[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3888 VPWR a_27479_9839# a_27647_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3889 a_22547_4221# a_21923_3855# a_22439_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3890 a_20188_12559# a_19789_12559# a_20062_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3891 a_20917_15279# tdc0.r_ring_ctr[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3892 VPWR tdc1.w_ring_norsz[30] a_8491_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3894 VGND a_27958_5461# a_27916_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3895 _077_ a_9963_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3896 VPWR a_4503_12533# a_4490_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3897 _130_ a_11713_6691# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X3898 VGND tdc1.w_ring_norsz[4] tdc1.w_ring_int_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3899 a_9103_4659# net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X3901 VPWR a_19567_14013# a_19735_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3902 VGND a_28291_6549# a_28249_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3903 tdc1.w_ring_norsz[2] tdc1.w_ring_int_norsz[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3905 a_20985_2767# tdc1.r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R51 VGND net71 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3906 VGND _158_ a_6824_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3907 a_8183_4703# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3908 VPWR a_6798_9813# a_6725_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3910 a_12552_8041# a_12153_7669# a_12426_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3912 VGND _182_ a_5449_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X3913 VGND tdc1.w_ring_int_norsz[23] tdc1.w_ring_norsz[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3914 VPWR _124_ a_11878_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X3916 _090_ a_21095_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3917 a_22178_13103# a_21739_13109# a_22093_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3918 a_22271_15101# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3919 a_7841_15657# a_6651_15285# a_7732_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3920 a_13441_6581# a_13275_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3921 a_4195_8573# a_3413_8207# a_4111_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3922 VPWR _193_ a_14008_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X3923 VPWR net31 a_16679_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3925 VGND net31 a_20359_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3926 a_19587_3689# a_19071_3317# a_19492_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3927 VGND a_9466_8319# a_9424_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
R52 net53 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3928 _019_ a_6291_5193# a_6541_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X3930 VGND net19 a_26615_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3931 a_18866_10927# a_18593_10933# a_18781_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3932 a_5069_11471# a_4903_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3933 net8 a_15023_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X3934 _103_ a_23947_12809# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3936 a_16937_13103# a_16403_13109# a_16842_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3937 a_4415_13647# _158_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X3938 tdc0.w_ring_norsz[25] tdc0.w_ring_int_norsz[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3940 VPWR net26 a_8583_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3941 a_10225_13647# tdc0.r_ring_ctr[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3942 VGND net7 a_6467_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3943 VPWR a_6791_11636# tdc0.w_ring_buf[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3944 VPWR a_12077_16341# a_11967_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3945 a_21457_12015# tdc0.w_ring_norsz[27] a_21373_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3946 VPWR _065_ a_19163_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3947 a_14725_11305# a_13735_10933# a_14599_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3948 a_4582_5309# a_3505_4943# a_4420_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3949 a_28694_7637# a_28526_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3952 VPWR _075_ a_24213_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3954 VPWR _067_ a_26329_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3955 a_22271_15101# a_21647_14735# a_22163_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3956 VGND a_6291_5193# _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X3957 VGND a_10018_11989# a_9976_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3958 VPWR tdc0.w_ring_norsz[18] a_26063_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3959 a_21247_15823# a_20801_15823# a_21151_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3960 a_19066_7895# a_19535_7637# a_19479_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X3961 VGND _060_ a_7705_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3962 VGND a_29119_9813# a_29077_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3963 VGND tdc1.w_ring_norsz[20] tdc1.w_ring_int_norsz[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3964 tdc1.w_ring_norsz[11] tdc1.w_ring_int_norsz[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3965 tdc1.r_dly_store_ring[26] a_29119_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3967 a_17555_7284# tdc1.w_ring_norsz[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3970 VPWR net9 a_6283_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3971 a_17119_4221# _057_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3972 VGND tdc1.w_ring_norsz[8] tdc1.w_ring_norsz[24] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3973 a_21307_5309# a_20525_4943# a_21223_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3974 a_8102_9839# a_7663_9845# a_8017_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3975 VPWR a_6119_7387# a_6035_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3976 a_6980_4917# tdc1.w_ring_buf[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3977 a_11219_14887# tdc0.r_ring_ctr[4] a_11393_14763# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3978 VGND net6 a_16771_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
R53 VGND net62 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3979 tdc1.w_ring_buf[27] a_28179_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3981 a_21751_9295# _080_ a_21644_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3982 a_23558_9839# a_23119_9845# a_23473_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3983 net25 a_15719_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3984 VGND net22 tdc0.w_ring_norsz[28] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3985 a_15283_8457# a_15335_8181# _066_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3986 VGND net69 tdc1.w_ring_int_norsz[24] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3987 a_6725_9839# a_6191_9845# a_6630_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3988 VGND a_20810_13621# a_20739_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3990 a_17100_14165# net33 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3991 a_10689_3855# _166_ a_10607_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3992 VPWR a_9103_4659# net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3993 VGND a_21923_4399# _166_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3994 a_22344_3855# _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3996 VGND a_14427_12724# tdc0.w_ring_buf[29] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3997 VPWR tdc1.r_ring_ctr[3] a_22373_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3998 a_20387_5487# a_19605_5493# a_20303_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3999 uo_out[3] a_25348_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4000 VPWR tdc0.w_ring_norsz[5] a_11885_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4002 VPWR a_17251_9813# a_17167_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4003 VGND a_30537_7895# a_30350_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X4004 a_22937_12015# tdc0.w_ring_int_norsz[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4005 tdc1.w_ring_norsz[13] tdc1.w_ring_norsz[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4007 a_17682_13621# a_17475_13621# a_17858_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4009 a_14427_12724# tdc0.w_ring_norsz[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4010 a_5955_9622# a_5773_9622# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4011 _045_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4013 a_12242_5309# a_11969_4943# a_12157_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4014 VGND a_20603_13621# a_20610_13921# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4015 a_21716_15823# a_20635_15823# a_21369_16065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4017 tdc0.r_dly_store_ctr[14] a_6027_13915# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4019 a_6756_10217# a_6357_9845# a_6630_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4020 a_17611_13647# a_17475_13621# a_17191_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4021 VGND net19 tdc1.w_ring_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4022 a_15564_11471# tdc0.r_dly_store_ring[13] a_15261_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X4023 a_18869_15823# a_18703_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4024 VPWR net27 a_2327_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4025 tdc0.r_dly_store_ctr[13] a_8235_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4027 a_26777_13423# tdc0.r_dly_store_ctr[2] a_26431_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4028 a_10018_10901# a_9850_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4029 a_24205_10933# a_24039_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4030 VPWR _131_ a_10395_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4031 VGND a_25348_10633# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4032 tdc0.r_ring_ctr[3] a_23087_15583# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4034 a_11131_9955# _136_ a_11059_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4035 a_13883_3689# a_13533_3317# a_13788_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4036 VPWR net7 a_6467_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4037 VPWR a_6430_6549# a_6357_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4038 _105_ a_25511_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4039 VGND a_18671_14495# a_18605_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4040 VGND a_20735_3017# _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X4041 VGND net38 tdc0.w_ring_int_norsz[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4042 a_9843_14735# _156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X4043 VGND _063_ a_4025_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4044 VGND net26 a_7663_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4045 VPWR _166_ a_11895_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X4046 a_12981_3631# tdc1.r_ring_ctr[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4048 tdc1.w_ring_buf[1] a_23119_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4049 tdc1.w_ring_norsz[27] net18 a_27897_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4050 a_7072_15645# _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4051 _120_ a_13551_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X4052 tdc1.w_ring_norsz[9] tdc1.w_ring_int_norsz[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4054 a_23837_5487# a_23303_5493# a_23742_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4055 a_5823_8457# tdc1.w_ring_norsz[0] a_6077_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4056 VGND net72 tdc1.w_ring_int_norsz[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4057 _074_ _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4059 a_10861_13647# a_9871_13647# a_10735_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4060 a_6888_3855# _029_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4061 a_7829_9845# a_7663_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4062 a_15647_14013# a_15023_13647# a_15539_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4065 a_27038_11989# a_26870_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4066 a_12150_10749# a_11711_10383# a_12065_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4067 VGND net26 a_3247_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4068 a_19692_4777# a_18777_4405# a_19345_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4069 a_20881_14735# tdc0.r_ring_ctr[1] a_20809_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4070 VGND tdc0.w_ring_norsz[31] tdc0.w_ring_int_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4071 a_25033_3855# a_24867_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4073 a_23201_11721# net24 tdc0.w_ring_norsz[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4074 _065_ a_16771_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R54 VGND uio_oe[5] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4076 a_8151_13103# a_7369_13109# a_8067_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4077 a_19695_3311# _048_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4081 a_19310_10495# a_19142_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4083 tdc0.r_dly_store_ring[24] a_10443_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4084 a_16677_14985# _154_ a_16595_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4086 a_18795_13103# _072_ a_18877_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4087 tdc0.r_ring_ctr[7] a_7907_15583# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4088 VGND _196_ _056_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4089 a_28621_8757# a_28455_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4090 VGND tdc0.w_ring_norsz[27] tdc0.w_ring_int_norsz[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4091 VPWR tdc0.w_ring_norsz[6] a_8113_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4092 a_13905_13647# tdc0.r_ring_ctr[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4093 a_22665_8457# tdc1.w_ring_norsz[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4094 VPWR a_10975_8751# _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4096 VPWR a_22636_3689# a_22811_3615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4097 _014_ a_12823_16073# a_13073_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X4099 a_9514_3901# _175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4100 a_9811_4737# tdc1.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4101 VPWR net29 a_13735_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4102 net16 a_14800_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4103 a_27705_5487# tdc1.w_ring_buf[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4104 a_5859_14013# a_4995_13647# a_5602_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4105 tdc1.w_ring_int_norsz[4] net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4106 a_8901_3677# a_8857_3285# a_8735_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4108 a_13243_5705# net30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4109 VPWR _064_ a_15701_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4110 a_23569_12015# net46 tdc0.w_ring_int_norsz[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4111 VGND net15 tdc1.w_ring_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4112 a_5353_12015# net20 tdc0.w_ring_norsz[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4113 tdc0.r_dly_store_ctr[10] a_24427_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4115 a_15753_15599# _152_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4116 a_10147_13103# _077_ a_10229_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4117 a_26251_11471# _092_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
X4118 a_21555_4765# tdc1.r_ring_ctr[2] a_21449_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4120 VGND tdc1.w_ring_norsz[11] tdc1.w_ring_norsz[27] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4121 net23 a_13735_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4122 VPWR a_17682_13621# a_17611_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4123 _156_ a_16127_14557# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X4124 a_15801_13647# a_15757_13889# a_15635_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4125 VPWR a_15828_4943# a_16003_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4126 VPWR _070_ a_19713_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4127 VPWR a_16587_8207# _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4128 a_18776_9071# a_18243_8751# _081_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4129 VPWR net36 a_28087_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4131 VPWR _154_ a_16845_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4132 a_7443_4777# a_6927_4405# a_7348_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4134 VPWR _158_ a_3689_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4135 VGND a_14583_13077# a_14541_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4136 VGND a_12403_8970# tdc1.w_ring_buf[24] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4138 VGND _103_ a_24683_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4139 _067_ a_11987_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4140 VPWR net20 _044_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4141 a_17195_2767# a_16679_2767# a_17100_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4142 a_13991_3311# a_13367_3317# a_13883_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4143 _048_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4144 a_9213_8207# tdc1.w_ring_buf[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4145 VPWR a_8183_4703# a_8170_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4147 VGND _072_ a_11505_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X4149 a_3505_6031# a_3339_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4150 _094_ a_20157_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4151 a_3505_4943# a_3339_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4152 VGND a_16155_7895# _119_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4153 VPWR a_11582_13077# a_11509_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4154 a_6630_12925# a_6357_12559# a_6545_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4155 VGND a_20083_8751# _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4157 tdc0.w_ring_buf[21] a_13459_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4159 a_13814_11471# _086_ a_13645_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X4160 a_21369_16065# a_21151_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4162 VGND net7 a_3339_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4166 VGND net41 tdc0.w_ring_int_norsz[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4167 a_3965_10749# a_3431_10383# a_3870_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4168 _142_ a_20083_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X4169 a_7642_13103# a_7203_13109# a_7557_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4170 a_24094_4373# a_23926_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4171 a_5043_11146# tdc0.w_ring_norsz[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4173 VPWR tdc0.w_ring_int_norsz[14] a_12889_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4174 VPWR tdc0.r_ring_ctr[8] a_15115_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4175 VGND a_15351_14423# _002_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4176 a_29871_7485# a_29173_7119# a_29614_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4177 a_7393_8457# tdc1.w_ring_norsz[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4179 a_2894_10927# a_2807_11169# a_2490_11059# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X4181 VPWR net26 a_5087_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4183 a_14967_12015# a_14103_12021# a_14710_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4184 a_7732_15657# a_6817_15285# a_7385_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4185 a_22821_5865# a_21831_5493# a_22695_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4186 a_25382_5461# a_25214_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4188 a_9945_12015# a_9411_12021# a_9850_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4189 VGND a_22719_10357# a_22726_10657# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4190 tdc0.w_ring_norsz[26] net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4191 a_8289_3317# a_8123_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4192 VGND tdc1.r_dly_store_ring[21] a_16589_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4193 VGND net18 tdc1.w_ring_norsz[26] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4194 a_25033_3855# a_24867_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4195 a_25306_14191# a_24867_14197# a_25221_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4196 VGND net15 _060_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4198 a_14061_8235# net25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X4199 a_14637_12015# a_14103_12021# a_14542_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4200 a_11115_4007# tdc1.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4201 _144_ _141_ a_20917_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4202 VGND _193_ a_14442_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4203 a_19310_5055# a_19142_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4204 a_10124_9269# _139_ a_10512_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4205 a_20253_11471# tdc0.w_ring_buf[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4206 a_7548_3855# a_6467_3855# a_7201_4097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4209 a_24351_4399# a_23653_4405# a_24094_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4210 tdc1.r_dly_store_ctr[5] a_13203_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4211 VGND a_29035_9447# _096_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4212 VGND a_13882_6549# a_13840_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4213 VGND _069_ a_10872_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4214 VPWR a_13887_8359# _186_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4216 net18 a_26615_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X4218 tdc1.w_ring_buf[25] a_28271_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
R55 tt_um_hpretl_tt06_tdc_v2_93.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4219 a_8841_13109# a_8675_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4220 a_8888_16189# a_8451_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4221 _079_ _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X4222 VPWR a_12863_5719# tdc1.r_dly_store_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4223 _035_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4225 VPWR a_12410_5055# a_12337_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4226 a_15193_7119# tdc1.w_ring_buf[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4227 tdc0.w_ring_norsz[9] tdc0.w_ring_int_norsz[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4228 tdc1.r_ring_ctr[12] a_8183_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4229 VPWR net41 a_27351_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X4230 a_12058_9661# a_11785_9295# a_11973_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4231 a_5907_5487# tdc1.r_ring_ctr[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.153 ps=1.3 w=1 l=0.15
X4232 VGND net27 a_7939_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4233 _046_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4235 VGND _144_ _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4236 VGND a_9963_8751# _077_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4237 VPWR a_27951_12247# tdc0.r_dly_store_ring[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4238 a_23389_8457# tdc1.w_ring_norsz[18] a_23305_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4239 VGND _066_ a_15553_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4240 VGND net22 tdc0.w_ring_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4241 tdc1.r_ring_ctr[11] a_16003_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4242 VGND ui_in[5] a_15575_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4243 _058_ net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4244 a_27069_8751# tdc1.w_ring_norsz[25] a_26985_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4246 tdc1.r_ring_ctr[0] a_20327_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4247 a_24462_11989# a_24294_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4248 a_13551_10633# _071_ a_13633_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4249 tdc0.r_dly_store_ctr[12] a_7223_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4250 a_15057_9839# _064_ a_14973_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4251 a_14541_13481# a_13551_13109# a_14415_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4252 a_9595_7663# _071_ a_9677_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4253 a_17095_13799# a_17191_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4255 VGND tdc1.r_dly_store_ring[10] a_29469_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4256 VGND a_24849_9839# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4257 tdc0.r_dly_store_ring[15] a_7223_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4258 VGND tdc0.w_ring_int_norsz[31] tdc0.w_ring_norsz[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4259 a_5720_4943# tdc1.r_ring_ctr[12] a_5417_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X4260 VGND a_29119_7637# a_29077_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4261 a_24294_12015# a_24021_12021# a_24209_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4262 a_19878_5487# a_19605_5493# a_19793_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4263 a_25129_5487# tdc1.w_ring_buf[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4265 VPWR a_15256_10535# _117_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X4266 a_3439_14191# _158_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4267 a_13882_14165# a_13714_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4268 a_15033_3855# _176_ a_14951_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4269 VPWR a_9006_7231# a_8933_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4270 tdc1.r_ring_ctr[7] a_7723_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4271 a_20522_6397# a_20083_6031# a_20437_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4272 VPWR tdc0.w_ring_buf[0] a_18059_16375# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X4275 a_12153_7669# a_11987_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4277 a_27066_11204# a_26866_11049# a_27215_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4278 a_9850_10927# a_9577_10933# a_9765_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4279 VPWR a_7539_14495# a_7526_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4280 tdc1.w_ring_norsz[31] tdc1.w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4281 VPWR tdc0.w_ring_int_norsz[22] a_11417_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4282 tdc0.r_ring_ctr[5] a_12875_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4283 a_6503_10749# a_5639_10383# a_6246_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4284 a_15809_12234# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4286 VGND net20 tdc0.w_ring_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4287 a_26859_11145# net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4288 VGND tdc1.w_ring_int_norsz[16] tdc1.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4289 VGND _175_ a_14073_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4290 a_5249_9129# a_4259_8757# a_5123_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4291 VGND net10 a_13643_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4292 VPWR _085_ a_25071_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4293 a_3526_10927# a_2768_11043# a_2963_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X4294 a_14899_15797# _040_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4295 a_22569_12015# tdc0.w_ring_int_norsz[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4296 a_7894_15279# a_6817_15285# a_7732_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4297 a_6173_10749# a_5639_10383# a_6078_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4298 a_10401_11305# a_9411_10933# a_10275_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
R56 VGND uio_oe[1] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4299 a_23469_5493# a_23303_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4300 a_28897_6575# tdc1.r_dly_store_ring[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4301 VGND net23 tdc0.w_ring_norsz[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4302 tdc1.w_ring_norsz[24] net16 a_12073_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4303 tdc0.w_ring_buf[10] a_24775_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4304 a_15025_7779# _119_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4307 a_25306_13103# a_24867_13109# a_25221_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4309 a_9677_7983# tdc1.r_dly_store_ring[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4310 VGND _086_ a_24683_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4311 a_27866_6549# a_27698_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4312 a_13921_7983# _076_ a_13511_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4314 VPWR a_2511_14191# net28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4315 a_6739_13897# tdc0.r_ring_ctr[13] a_6521_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4316 a_11792_12015# _125_ a_11706_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4317 a_9411_9839# _071_ a_9589_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4318 a_9167_14763# tdc0.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4319 tdc0.w_ring_int_norsz[26] tdc0.w_ring_norsz[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4320 tdc1.w_ring_norsz[30] net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4321 VGND a_8270_9813# a_8228_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4322 a_21844_10217# a_21445_9845# a_21718_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4323 VPWR a_19735_10651# a_19651_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4325 a_28253_7669# a_28087_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4326 tdc1.r_dly_store_ring[1] a_24151_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4328 a_17836_14557# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4329 a_25639_5487# a_24941_5493# a_25382_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4330 a_28809_8751# tdc1.w_ring_buf[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4331 tdc1.r_dly_store_ring[19] a_25071_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4332 a_22443_15657# a_21997_15285# a_22347_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4333 tdc1.r_dly_store_ctr[13] a_6855_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4334 a_8653_8041# a_7663_7669# a_8527_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4335 a_3413_8207# a_3247_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4336 VGND a_23726_9813# a_23684_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4337 a_28897_6575# tdc1.r_dly_store_ring[12] a_28813_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4338 _074_ a_14794_9922# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X4339 _071_ a_15159_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4340 VPWR a_26479_11159# tdc0.r_dly_store_ring[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4341 a_16968_13481# a_16569_13109# a_16842_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4342 a_16289_6031# a_15299_6031# a_16163_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4343 VPWR _069_ a_27057_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X4344 VPWR tdc1.w_ring_norsz[28] a_26053_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4345 a_13511_7895# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
R57 net49 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4348 _116_ a_15023_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4349 a_9963_5487# _077_ a_10045_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4350 VPWR a_30039_7387# a_29955_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R58 tt_um_hpretl_tt06_tdc_v2_89.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4352 a_15990_5309# a_14913_4943# a_15828_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4353 a_24683_10159# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4354 VGND tdc1.w_ring_norsz[29] a_15023_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4355 VGND a_11987_9839# _067_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4356 VGND tdc1.w_ring_norsz[9] a_27903_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4357 VGND _121_ a_15420_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4358 VGND a_9503_9295# _086_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4359 a_4880_14735# a_3965_14735# a_4533_14977# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4360 a_10512_9545# _134_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4361 VGND a_20655_12827# a_20613_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4363 a_16937_7369# tdc1.w_ring_norsz[22] a_16853_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4365 a_19655_8235# _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4367 a_21721_3317# a_21555_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4368 a_20648_6031# a_20249_6031# a_20522_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4369 VPWR a_25899_14165# a_25815_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4371 VGND net35 a_23211_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4373 VGND _055_ a_7245_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4374 VPWR tdc1.w_ring_norsz[31] a_6733_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4375 a_13905_13103# tdc0.w_ring_buf[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4376 a_21285_14985# _140_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4377 VPWR tdc1.w_ring_norsz[12] a_27167_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4378 a_19893_15823# a_18703_15823# a_19784_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4380 a_17191_13621# a_17475_13621# a_17410_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4381 _069_ a_10975_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4382 a_28694_9813# a_28526_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4383 a_24849_9839# a_25071_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4384 VPWR a_12375_14165# a_12291_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4385 a_6246_10495# a_6078_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4386 a_18866_10927# a_18427_10933# a_18781_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4387 VGND a_4463_10651# a_4421_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4389 _065_ a_16771_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4390 tdc1.r_dly_store_ring[31] a_9431_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4391 VPWR a_5123_9839# a_5291_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4392 tdc1.w_ring_int_norsz[23] net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4393 a_3201_11293# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X4396 VPWR net15 _063_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4397 VPWR a_6246_10495# a_6173_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4398 VPWR tdc0.r_ring_ctr[4] a_10881_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4399 VGND net12 a_27535_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4400 VPWR a_8723_11636# tdc0.w_ring_buf[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4402 a_10919_5309# a_10221_4943# a_10662_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4404 a_3115_9813# net28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X4405 VGND tdc0.r_ring_ctr[2] a_20881_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4406 _015_ _153_ a_16017_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X4407 VGND a_16595_14985# _001_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X4409 VPWR tdc1.w_ring_int_norsz[21] a_17581_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4410 a_29871_7485# a_29007_7119# a_29614_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4411 a_4866_8725# a_4698_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4412 VPWR _066_ a_9677_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4413 a_11782_14191# a_11343_14197# a_11697_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4414 a_19142_14013# a_18703_13647# a_19057_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4415 VGND _081_ a_19741_8235# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4416 VPWR net31 a_18703_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4417 a_17811_5487# a_17029_5493# a_17727_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4418 VPWR a_21912_6575# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4420 a_20138_15823# _032_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4421 a_17836_14557# _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4422 a_11965_13481# a_10975_13109# a_11839_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4423 a_7201_4097# a_6983_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4424 VGND tdc1.w_ring_norsz[27] tdc1.w_ring_int_norsz[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4426 tdc0.w_ring_buf[2] a_23855_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4427 net41 a_26983_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X4428 a_20441_12015# net41 tdc0.w_ring_int_norsz[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4430 a_6743_7663# tdc1.w_ring_int_norsz[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4431 a_25815_13103# a_25033_13109# a_25731_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4434 a_11491_2767# a_11141_2767# a_11396_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4435 VPWR a_12226_9407# a_12153_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4437 VGND net43 tdc0.w_ring_int_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4438 VPWR net27 a_7203_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4439 a_25472_8181# _101_ a_25864_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X4440 a_25121_9129# a_24131_8757# a_24995_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4441 a_5602_13759# a_5434_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4442 VPWR tdc0.r_ring_ctr[10] a_15627_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X4443 tdc1.r_dly_store_ctr[2] a_21391_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4444 VGND a_8183_4703# tdc1.r_ring_ctr[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4445 VPWR _076_ a_9963_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4446 VGND a_16279_13621# a_16213_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4447 a_9371_4007# a_9514_3901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X4448 VGND a_5859_14013# a_6027_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4449 a_17191_13621# a_17482_13921# a_17433_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4450 VPWR a_14623_3615# tdc1.r_ring_ctr[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4451 VPWR a_8067_13103# a_8235_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4452 VGND _043_ a_15801_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4453 VGND net25 a_9849_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X4455 VGND _171_ a_9740_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X4456 VGND _041_ a_17089_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4457 VGND a_8067_13103# a_8235_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4458 _121_ a_15025_7779# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X4459 a_11325_7663# tdc1.w_ring_norsz[7] a_11241_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4460 VGND tdc1.w_ring_norsz[14] a_12539_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4461 a_25182_10383# _105_ a_25348_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4462 VGND _123_ a_11435_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4463 tdc0.w_ring_norsz[27] tdc0.w_ring_norsz[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4464 tdc0.w_ring_buf[4] a_20727_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4466 a_29173_8207# a_29007_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4467 VPWR a_24849_9839# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4468 a_24293_12559# tdc0.r_dly_store_ring[19] a_23947_12809# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
R59 tt_um_hpretl_tt06_tdc_v2_87.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4469 VGND net23 tdc0.w_ring_norsz[29] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4470 a_16913_756# ui_in[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4471 a_5123_9839# a_4259_9845# a_4866_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4472 VGND net17 tdc1.w_ring_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4473 a_17010_13077# a_16842_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4474 VGND a_20690_6143# a_20648_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4475 VGND net26 a_5087_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4476 a_2932_14165# net28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4478 _146_ a_10363_15617# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X4479 _057_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4481 a_8971_15965# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4482 a_27958_5461# a_27790_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4483 a_9647_14709# _143_ a_10045_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X4484 a_17303_3133# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4486 tdc1.r_dly_store_ctr[9] a_22863_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4487 a_11969_4943# a_11803_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4488 a_25731_4221# a_24867_3855# a_25474_3967# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4489 VGND _188_ a_13553_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4490 a_4682_12559# _046_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4491 tdc1.w_ring_norsz[0] tdc1.w_ring_int_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X4492 a_10781_10383# tdc0.r_dly_store_ring[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4493 a_18877_8457# tdc1.r_dly_store_ring[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
R60 tdc0.g_ring3[29].stg01_56.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4494 a_9282_13077# a_9114_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4495 a_11877_10383# a_11711_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4496 a_9577_10933# a_9411_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4500 VGND a_5043_10548# tdc0.w_ring_buf[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4501 VPWR a_5123_8751# a_5291_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4502 VPWR net31 a_16863_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4503 a_9757_6031# a_8767_6031# a_9631_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4505 a_20433_8029# _065_ a_20333_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X4506 VGND tdc1.w_ring_norsz[26] a_27443_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4508 VGND tdc1.w_ring_int_norsz[4] tdc1.w_ring_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4509 tdc0.w_ring_int_norsz[0] net59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4510 _110_ a_12447_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4511 VPWR a_8451_15797# tdc0.r_ring_ctr[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X4513 a_10221_4943# a_10055_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4515 a_20735_3017# tdc1.r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4516 a_20889_11471# a_19899_11471# a_20763_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
R61 tt_um_hpretl_tt06_tdc_v2_86.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4517 a_8067_13103# a_7203_13109# a_7810_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4518 VGND tdc1.w_ring_norsz[30] a_8491_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4519 tdc1.w_ring_buf[15] a_7571_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4520 VPWR _175_ _176_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4521 a_12153_9661# a_11619_9295# a_12058_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4522 a_16569_13109# a_16403_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4524 a_7017_14165# a_6799_14569# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4527 tdc0.w_ring_buf[18] a_26063_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4528 a_16935_16189# a_16311_15823# a_16827_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4529 a_18877_13103# tdc0.r_dly_store_ring[9] a_18795_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4532 tdc0.w_ring_int_norsz[28] net55 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4533 tdc1.w_ring_norsz[24] tdc1.w_ring_int_norsz[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4534 a_13840_14569# a_13441_14197# a_13714_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4535 VPWR a_9963_8751# _077_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4537 VPWR _166_ a_10291_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X4538 a_25397_7119# tdc1.r_dly_store_ring[19] a_24959_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4539 _175_ a_11067_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X4541 tdc0.r_dly_store_ring[17] a_17435_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4543 a_17935_2741# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4544 a_8293_12015# tdc0.w_ring_buf[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4545 VGND a_17283_14709# net33 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4546 a_20810_13621# a_20610_13921# a_20959_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4547 VGND a_14983_14165# net10 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4548 a_22855_10383# a_22719_10357# a_22435_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4549 a_14209_9111# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X4550 a_14623_3615# a_14448_3689# a_14802_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4551 a_4588_7637# net15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4552 tdc1.r_dly_store_ring[22] a_11823_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4553 a_10493_10159# tdc0.r_dly_store_ring[23] a_10147_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4554 VGND a_24259_14191# a_24427_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4555 VGND a_4503_12533# a_4437_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4557 a_10229_13103# tdc0.r_dly_store_ctr[14] a_10147_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4559 VPWR a_7699_6397# a_7867_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4560 VGND tdc0.w_ring_int_norsz[15] tdc0.w_ring_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4561 a_19973_5487# a_19439_5493# a_19878_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4563 VPWR a_26615_7119# net18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4564 VGND a_25474_14165# a_25432_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4565 VPWR tdc0.r_ring_ctr[1] a_19715_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X4566 _050_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4567 VGND _086_ a_5236_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X4568 a_17011_3855# a_16661_3855# a_16916_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4569 VGND a_7055_9839# a_7223_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4570 net37 a_3247_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4571 VPWR a_21115_6299# a_21031_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4572 a_3689_14191# tdc0.r_ring_ctr[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4573 VGND a_6791_11636# tdc0.w_ring_buf[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4574 a_14913_4943# a_14747_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4575 a_13633_7369# _084_ a_13551_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4576 VPWR a_21707_7881# a_21714_7785# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4578 a_22547_4221# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4579 a_14342_10901# a_14174_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4580 VGND a_19459_10901# a_19417_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4581 _147_ tdc0.r_ring_ctr[5] a_11343_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4582 VGND _195_ _032_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4583 VPWR a_18703_14735# _195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4585 VPWR _083_ a_24591_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X4586 a_22565_15253# a_22347_15657# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4590 a_24604_11305# a_24205_10933# a_24478_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4591 a_19223_4777# a_18777_4405# a_19127_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4593 a_27698_6575# a_27259_6581# a_27613_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4594 a_14174_10927# a_13901_10933# a_14089_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4595 a_14703_12724# tdc0.w_ring_norsz[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4596 VPWR a_27351_8207# net40 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4597 a_5123_8751# a_4259_8757# a_4866_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4598 a_15627_14709# tdc0.r_ring_ctr[8] a_16025_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X4599 VPWR a_8543_15253# _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X4600 VGND net16 tdc1.w_ring_norsz[23] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4602 VGND _196_ _051_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4604 VGND a_25731_13103# a_25899_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4606 tdc1.w_ring_int_norsz[11] net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4607 VGND a_3024_8725# _621_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4608 VPWR tdc0.r_ring_ctr[11] a_15654_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X4609 tdc1.r_ring_ctr[6] a_9379_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4610 a_12889_12015# tdc0.w_ring_norsz[30] a_12805_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4611 a_9976_12393# a_9577_12021# a_9850_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4614 a_26420_11721# _098_ a_26251_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X4615 _127_ a_9963_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4616 _062_ net15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4617 a_8929_12393# a_7939_12021# a_8803_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4619 a_14668_12393# a_14269_12021# a_14542_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4621 a_6749_12015# tdc0.w_ring_norsz[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4622 a_13919_4512# tdc1.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X4623 a_24683_10159# a_25071_9813# a_24849_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4624 a_25221_14191# tdc0.r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4626 a_18114_4765# _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4627 VGND tdc0.w_ring_norsz[10] tdc0.w_ring_norsz[26] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4628 tdc1.r_dly_store_ctr[7] a_9615_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4630 tdc1.w_ring_int_norsz[6] tdc1.w_ring_norsz[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4632 a_3413_8207# a_3247_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4633 tdc0.r_ring_ctr[0] a_19959_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X4634 VPWR a_24002_14165# a_23929_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4635 a_13717_13647# a_13551_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4636 a_16385_3631# tdc1.r_ring_ctr[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4637 tdc1.r_dly_store_ring[6] a_18171_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4638 VGND net21 tdc0.w_ring_norsz[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4639 VPWR a_25899_4123# a_25815_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4640 VGND a_16331_6299# a_16289_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4641 a_21259_16189# _033_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4642 a_14255_15823# a_13809_15823# a_14159_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4644 VPWR _175_ a_12981_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4645 _082_ a_19655_8235# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X4647 VGND _087_ a_20175_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4649 VGND a_12875_14709# a_12809_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4650 VPWR a_17413_4373# a_17303_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4651 VGND a_9127_16060# a_9058_16189# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4652 VGND net28 a_8675_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4653 a_20825_4105# _163_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4654 VGND net34 a_24867_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4656 tdc0.r_dly_store_ctr[6] a_10903_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4657 a_24849_13897# tdc0.r_dly_store_ctr[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4659 a_29446_7485# a_29007_7119# a_29361_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4660 a_10323_7779# _133_ a_10241_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4662 a_22728_14735# a_21813_14735# a_22381_14977# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4663 _056_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4664 VPWR _143_ a_11049_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4665 a_20729_9955# _110_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4667 a_6541_5193# tdc1.r_ring_ctr[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4668 VGND net27 a_2327_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4669 a_19784_15823# a_18869_15823# a_19437_16065# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4670 a_24213_6031# tdc1.r_dly_store_ctr[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4671 VPWR a_27463_11989# a_27379_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4672 VGND tdc0.r_ring_ctr[11] a_16403_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X4673 a_22086_14013# a_21647_13647# a_22001_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4675 VGND a_24646_6549# a_24604_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4676 a_15281_4105# tdc1.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X4677 VGND a_6430_6549# a_6388_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4678 tdc1.r_dly_store_ctr[15] a_6119_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4679 net23 a_13735_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4680 a_11141_2767# a_10975_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4681 tdc0.w_ring_norsz[17] net23 a_16213_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4683 VGND _148_ a_8912_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X4685 a_8527_9839# a_7829_9845# a_8270_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4686 a_26127_9545# _096_ a_26055_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4687 a_28951_9839# a_28087_9845# a_28694_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4688 a_15189_3855# _176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4689 a_13637_7663# _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X4690 a_12731_3311# _175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4692 VPWR a_5291_9813# a_5207_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4693 a_27813_7663# tdc1.w_ring_int_norsz[27] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4694 _069_ a_10975_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4695 uo_out[1] a_24849_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4696 a_27824_6953# a_27425_6581# a_27698_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4697 tdc1.w_ring_int_norsz[9] tdc1.w_ring_norsz[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4698 tdc0.w_ring_int_norsz[22] net49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4699 VPWR tdc0.r_ring_ctr[1] a_20083_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X4700 a_22068_14735# _008_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4701 tdc1.w_ring_int_norsz[12] net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4702 net39 a_17375_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4703 tdc1.r_dly_store_ring[2] a_22311_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4704 tdc1.r_dly_store_ring[16] a_8327_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4705 VGND a_11763_8725# net30 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4706 tdc1.w_ring_buf[1] a_23119_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4707 VPWR a_8399_3855# _196_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4708 a_17397_5487# a_16863_5493# a_17302_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4709 a_12778_4373# a_12610_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4710 VGND a_25472_8181# _102_ VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X4711 _008_ _141_ a_21285_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4712 VGND a_4595_4917# a_4529_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4713 a_14724_15823# a_13643_15823# a_14377_16065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4716 a_20437_6031# tdc1.w_ring_buf[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4717 tdc0.r_ring_ctr[14] a_4503_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4718 VPWR a_11035_3543# _169_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4719 a_21718_8751# a_21279_8757# a_21633_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4720 a_7526_14191# a_6449_14197# a_7364_14569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4721 VPWR a_24903_10927# a_25071_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4722 a_11417_10927# tdc0.w_ring_norsz[6] a_11333_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4723 a_7734_8751# a_7295_8757# a_7649_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4724 a_3273_11293# a_2894_10927# a_3201_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4726 tdc1.r_dly_store_ctr[12] a_20471_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4729 a_28694_9813# a_28526_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4730 VGND tdc0.w_ring_norsz[4] tdc0.w_ring_int_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4731 a_22926_10357# a_22726_10657# a_23075_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X4733 a_29062_8725# a_28894_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4734 a_29445_9129# a_28455_8757# a_29319_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4737 a_22557_11721# net47 tdc0.w_ring_int_norsz[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4738 a_4117_4943# a_4073_5185# a_3951_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4740 a_6191_14735# _159_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X4741 VGND a_17746_12671# a_17704_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4742 tdc1.r_dly_store_ctr[7] a_9615_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4744 a_3255_11721# _161_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4745 VGND a_10799_16073# _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X4746 a_11782_14191# a_11509_14197# a_11697_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4748 a_10799_16073# _143_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4749 a_20451_6575# _077_ a_20629_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4750 VPWR _083_ a_25493_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X4752 VGND net35 a_24867_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4754 VPWR tdc0.w_ring_norsz[3] a_23763_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4755 a_24209_12015# tdc0.w_ring_buf[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4756 a_23929_14191# a_23395_14197# a_23834_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4757 VGND net8 a_13367_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4758 a_24570_8751# a_24297_8757# a_24485_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4759 a_18781_10927# tdc0.w_ring_buf[28] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4760 VPWR _064_ a_15701_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4763 VGND a_9379_3615# a_9313_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4764 a_11145_6031# tdc1.w_ring_buf[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4765 VPWR tdc1.w_ring_int_norsz[18] a_24021_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4766 net28 a_2511_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4769 a_28714_12015# a_28467_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4771 VGND a_19459_6549# a_19417_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4772 tdc1.w_ring_int_norsz[22] net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4774 a_16301_7663# _066_ a_16155_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X4775 a_23726_9813# a_23558_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4776 tdc1.w_ring_norsz[7] tdc1.w_ring_norsz[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4777 _621_.X a_3024_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4780 VPWR a_12291_6183# _126_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4781 a_12793_4943# a_11803_4943# a_12667_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4782 tdc1.r_dly_store_ring[15] a_8695_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4783 a_14553_5487# tdc1.r_ring_ctr[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X4784 a_24646_6549# a_24478_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4785 a_29173_8207# a_29007_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4786 a_29572_7119# a_29173_7119# a_29446_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4787 VPWR net34 a_24867_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4788 VGND a_23259_7882# tdc1.w_ring_buf[18] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4789 _006_ _161_ a_3505_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X4790 net21 a_3484_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4791 VPWR _195_ _041_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4792 VGND _064_ _074_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4793 a_21349_4943# a_20359_4943# a_21223_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4794 VGND a_11950_14165# a_11908_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4795 VGND _092_ a_26251_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4796 a_17760_2767# a_16679_2767# a_17413_3009# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4797 a_12525_4399# tdc1.r_ring_ctr[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4798 a_8639_3689# a_8289_3317# a_8544_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4799 a_11623_12335# _130_ a_11792_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4800 VPWR a_16463_12533# net38 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4801 a_16757_13103# tdc0.w_ring_buf[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4802 VGND _082_ a_20083_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4803 VPWR a_7017_14165# a_6907_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4804 VPWR net31 a_20083_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4805 VGND net27 a_5639_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4806 a_11141_2767# a_10975_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4807 _190_ a_13814_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X4808 VPWR a_10275_12015# a_10443_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4809 a_4511_13647# tdc0.r_ring_ctr[14] a_4415_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X4810 VPWR a_11987_9839# _067_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4811 tdc0.w_ring_buf[1] a_19347_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4812 a_18003_12925# a_17139_12559# a_17746_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4813 VPWR _066_ a_10229_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4814 tdc0.w_ring_int_norsz[24] tdc0.w_ring_norsz[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4815 a_24052_4777# a_23653_4405# a_23926_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4817 VGND a_10275_12015# a_10443_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4818 a_19220_8457# _128_ a_18877_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X4819 a_19605_5493# a_19439_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4820 VPWR _065_ a_19899_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4822 a_16661_3855# a_16495_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4823 VPWR a_5291_8725# a_5207_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4825 VGND a_9799_6299# a_9757_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4826 VPWR _126_ a_11867_6691# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4827 VGND tdc1.w_ring_int_norsz[19] tdc1.w_ring_norsz[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4828 a_11785_9295# a_11619_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4829 a_17673_12925# a_17139_12559# a_17578_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4830 VPWR a_9103_4659# net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4831 VPWR tdc0.w_ring_int_norsz[7] a_7461_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4832 tdc1.w_ring_norsz[28] net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4834 a_3760_6031# _021_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4835 a_18243_9071# _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X4836 a_12778_4373# a_12610_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4837 VPWR tdc1.r_ring_ctr[13] _182_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4838 a_5055_14709# a_4880_14735# a_5234_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4839 tdc0.r_dly_store_ring[13] a_15135_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4840 a_21844_9129# a_21445_8757# a_21718_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4841 a_26431_13103# _072_ a_26513_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4842 _159_ tdc0.r_ring_ctr[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4843 a_7860_9129# a_7461_8757# a_7734_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4844 a_8780_14569# a_8381_14197# a_8654_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4845 a_23469_7369# tdc1.w_ring_norsz[19] a_23385_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4846 a_27036_7637# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4847 VPWR a_24243_13077# a_24159_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4848 VGND a_24887_15003# a_24845_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4849 VPWR a_28123_6575# a_28291_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4850 a_28123_6575# a_27425_6581# a_27866_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4851 VPWR net8 a_18611_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4853 a_3996_10383# a_3597_10383# a_3870_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4855 VGND tdc1.r_ring_ctr[2] a_20789_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4856 a_6817_15285# a_6651_15285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4857 a_13620_9269# _189_ a_14442_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4858 a_10124_9269# _083_ a_10512_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4859 a_23653_4405# a_23487_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4861 a_21717_7119# tdc1.r_dly_store_ring[18] a_21279_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4862 VPWR tdc0.w_ring_norsz[27] a_25971_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4863 VPWR a_24887_11989# a_24803_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4865 a_15278_7485# a_15005_7119# a_15193_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4866 VGND net44 tdc0.w_ring_int_norsz[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4867 VPWR tdc1.r_ring_ctr[8] a_14155_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X4868 a_28538_12292# a_28331_12233# a_28714_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4869 VGND tdc0.w_ring_norsz[29] tdc0.w_ring_int_norsz[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4870 a_12599_16671# a_12424_16745# a_12778_16733# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4872 a_22455_15279# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4873 a_28951_7663# a_28253_7669# a_28694_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4874 a_16301_10927# net23 tdc0.w_ring_norsz[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4875 a_14377_16065# a_14159_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4876 VPWR a_27036_7637# net17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4877 a_4379_10749# a_3597_10383# a_4295_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4878 a_26251_11471# _093_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4880 a_12587_8372# tdc1.w_ring_norsz[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4881 a_10275_12015# a_9411_12021# a_10018_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4882 a_7710_4221# a_6633_3855# a_7548_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4884 VPWR a_14307_14165# a_14223_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4885 a_18193_14557# a_18149_14165# a_18027_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4886 a_9127_16060# a_8932_16091# a_9437_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X4887 VGND a_11823_6299# a_11781_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4888 _164_ a_20635_4512# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4890 a_28467_12393# a_28331_12233# a_28047_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4892 a_15937_4943# a_14747_4943# a_15828_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4893 VGND net36 a_27351_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4894 VPWR a_29319_8751# a_29487_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4895 a_27069_12559# tdc0.r_dly_store_ring[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4896 _107_ a_28731_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4897 VGND a_29614_7231# a_29572_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4898 a_6813_8457# net15 tdc1.w_ring_norsz[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4899 a_25933_9071# tdc1.r_dly_store_ring[17] _079_ VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4900 VPWR tdc1.w_ring_int_norsz[31] a_8013_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4903 VGND a_22143_9839# a_22311_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4904 a_15256_10535# _114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X4907 a_10662_5055# a_10494_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4910 tdc0.r_ring_ctr[2] a_22903_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4912 VGND a_8971_11989# a_8929_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4913 a_8747_3311# a_8123_3317# a_8639_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4914 a_8838_7485# a_8399_7119# a_8753_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4915 a_21399_10535# tdc0.r_dly_store_ring[20] a_21545_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X4916 a_21356_12559# tdc0.r_dly_store_ring[1] a_21095_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4918 a_27769_5108# tdc1.w_dly_stop[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4919 a_8159_8751# a_7461_8757# a_7902_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4920 tdc0.r_dly_store_ring[5] a_17251_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4921 VGND tdc0.w_ring_int_norsz[12] tdc0.w_ring_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4922 a_19693_10383# a_18703_10383# a_19567_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4923 _124_ a_11435_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X4924 VPWR _143_ a_10239_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4925 a_25348_10633# _104_ a_25182_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X4926 VGND net24 tdc0.w_ring_norsz[27] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4927 tdc1.w_ring_int_norsz[7] net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4930 a_17738_4221# a_16661_3855# a_17576_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4931 VPWR a_17746_12671# a_17673_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4933 a_24393_6575# tdc1.w_ring_buf[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4934 a_6177_6575# tdc1.r_ring_ctr[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4935 a_12410_5055# a_12242_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4936 VPWR a_16279_13621# a_16266_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4937 a_28123_6575# a_27259_6581# a_27866_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4939 a_19723_15279# tdc0.r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4940 a_16661_3855# a_16495_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4941 a_8611_7663# a_7829_7669# a_8527_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4942 a_16209_14557# tdc0.r_ring_ctr[8] a_16127_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X4943 VGND net31 a_21279_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4944 a_3484_13077# net24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4945 a_14101_3285# a_13883_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4947 tdc1.r_ring_ctr[12] a_8183_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4948 VPWR _067_ a_18877_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4949 VPWR a_8971_15965# a_8932_16091# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4950 tdc1.r_ring_ctr[3] a_23179_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4951 a_22636_3689# a_21721_3317# a_22289_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
D0 VGND _110_ sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X4953 VGND a_23087_15583# a_23021_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4954 tdc1.w_ring_int_norsz[15] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4955 a_14447_4943# tdc1.r_ring_ctr[10] a_14351_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X4956 net17 a_27036_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4958 a_28253_9845# a_28087_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4960 _099_ a_18501_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4961 VGND a_15335_8181# _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4962 VGND a_29955_8983# _073_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4963 VPWR a_3392_8725# _620_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4964 VGND _035_ a_22609_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4965 _060_ net15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4966 net35 a_23080_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4967 tdc1.w_ring_int_norsz[1] tdc1.w_ring_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4969 a_13717_13647# a_13551_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4970 a_8105_12021# a_7939_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4971 VGND tdc0.w_ring_int_norsz[21] tdc0.w_ring_norsz[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4972 VGND net20 _046_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4974 VGND _171_ _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4975 a_20327_3615# a_20152_3689# a_20506_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4976 a_27951_12247# a_28047_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4977 VPWR _138_ a_10512_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X4979 net24 a_3799_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4980 a_13599_6196# tdc1.w_ring_norsz[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4981 _165_ a_21279_4765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X4982 VGND net26 a_5823_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4983 a_2525_11293# a_2490_11059# a_2287_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X4984 VGND tdc0.w_ring_buf[26] a_28885_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4985 VPWR a_23179_3829# a_23166_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4986 a_10018_10901# a_9850_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4987 VGND a_11792_12015# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4989 VPWR a_21399_10535# _109_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4990 a_3601_9295# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4991 tdc0.w_ring_int_norsz[4] net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4993 a_8159_8751# a_7295_8757# a_7902_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4994 VGND tdc1.w_ring_norsz[26] tdc1.w_ring_norsz[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4996 _027_ _169_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4997 VPWR a_11709_3009# a_11599_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4998 tdc1.w_ring_norsz[30] tdc1.w_ring_int_norsz[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5000 a_24435_4399# a_23653_4405# a_24351_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5001 VPWR _086_ a_24765_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5002 a_6204_10383# a_5805_10383# a_6078_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5004 VGND a_5231_4631# _020_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5005 tdc0.w_ring_int_norsz[26] net53 a_18249_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5006 VPWR a_10018_11989# a_9945_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5007 VPWR tdc0.w_ring_norsz[24] a_9135_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5008 a_25125_7369# tdc1.r_dly_store_ctr[3] a_25041_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5010 a_15553_11247# tdc0.r_dly_store_ring[21] a_15207_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5011 a_20538_13647# a_20223_13799# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5012 a_7093_4405# a_6927_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5013 VGND a_5417_4917# _183_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5015 a_13645_11721# tdc0.r_dly_store_ctr[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5017 a_15504_9295# _117_ a_15420_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5018 a_8964_7119# a_8565_7119# a_8838_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5019 VPWR a_26420_11721# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5020 a_17413_3009# a_17195_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5021 VGND _152_ a_15269_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X5022 a_11763_8725# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X5023 a_27421_12393# a_26431_12021# a_27295_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5024 a_22741_6281# net66 tdc1.w_ring_int_norsz[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5025 tdc1.r_dly_store_ring[30] a_9799_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5028 _051_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5030 VPWR _086_ a_4761_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X5031 a_12905_16073# _152_ a_12823_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5032 tdc1.w_ring_int_norsz[17] tdc1.w_ring_norsz[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5033 a_24861_13647# tdc0.r_dly_store_ctr[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X5034 VGND net34 a_24315_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5035 a_16017_16073# tdc0.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X5036 tdc0.r_ring_ctr[11] a_16279_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X5038 a_4237_9295# a_3247_9295# a_4111_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5040 VGND a_17740_10071# _122_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X5042 _086_ a_9503_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5043 a_26247_6281# _075_ a_26329_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5044 a_24131_6281# _077_ a_24213_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5045 a_26870_12015# a_26597_12021# a_26785_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5046 _072_ a_12539_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5047 tdc1.w_ring_buf[20] a_22935_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5048 VGND net38 tdc0.w_ring_int_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5049 VPWR a_19437_16065# a_19327_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5050 VGND a_19567_10749# a_19735_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5051 VGND tdc1.w_ring_norsz[12] a_27167_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5052 tdc0.w_ring_norsz[10] net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5053 a_23749_14191# tdc0.r_ring_ctr[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5056 net19 a_27411_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5057 VGND a_24243_13077# a_24201_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5058 VGND _195_ _035_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5062 tdc1.w_ring_int_norsz[9] net39 a_14385_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5063 a_25493_12015# tdc0.r_dly_store_ctr[10] a_25409_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5064 a_4880_14735# a_3799_14735# a_4533_14977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5065 a_17497_6575# net19 tdc1.w_ring_norsz[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5066 VGND a_10975_8751# _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X5067 a_8543_15253# a_8686_15395# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X5068 VGND tdc0.w_ring_norsz[1] a_19347_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5069 VGND net9 a_6283_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R62 net69 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5071 a_22001_13647# tdc0.r_ring_ctr[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5072 a_4682_7119# _063_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5073 VGND a_8723_11636# tdc0.w_ring_buf[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5075 a_11219_14887# tdc0.r_ring_ctr[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X5076 a_17405_12015# net56 tdc0.w_ring_int_norsz[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5078 a_10607_3855# _168_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5079 tdc1.r_dly_store_ring[5] a_17711_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5080 a_9127_16060# a_8971_15965# a_9272_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X5081 tdc1.r_dly_store_ring[19] a_25071_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5082 _040_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5083 VPWR _196_ _048_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5084 VPWR a_6521_13621# _160_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5085 a_14599_10927# a_13901_10933# a_14342_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5086 a_23983_9839# a_23119_9845# a_23726_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5087 VPWR a_15446_7231# a_15373_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5088 tdc1.r_dly_store_ring[27] a_30039_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5089 a_14174_10927# a_13735_10933# a_14089_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5090 a_24903_6575# a_24039_6581# a_24646_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5091 a_6687_6575# a_5823_6581# a_6430_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5092 a_20503_15253# _142_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X5093 tdc0.w_ring_buf[2] a_23855_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5094 a_20429_5865# a_19439_5493# a_20303_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5097 VGND net37 a_23671_15287# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
R63 net59 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5098 VGND a_21391_5211# a_21349_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5099 VGND _196_ _057_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5101 VGND a_9723_8573# a_9891_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5103 a_13729_7119# tdc1.r_dly_store_ctr[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X5105 tdc1.w_ring_norsz[4] tdc1.w_ring_norsz[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5106 _098_ a_25973_9301# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X5107 VGND a_10124_9269# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5109 VGND a_11219_14887# _145_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5110 a_15504_9295# _122_ a_15772_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5111 a_20253_11471# tdc0.w_ring_buf[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5112 VGND a_5510_11583# a_5468_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5113 VPWR net33 a_21739_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5114 VPWR a_9707_13077# a_9623_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5115 VPWR a_24849_9839# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5116 a_11049_16073# tdc0.r_ring_ctr[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5117 a_14265_6953# a_13275_6581# a_14139_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5118 VGND _065_ _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X5120 VPWR a_28951_7663# a_29119_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5121 a_7443_4777# a_7093_4405# a_7348_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5122 tdc0.w_dly_stop[5] a_3155_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5123 a_29361_7119# tdc1.w_ring_buf[27] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5124 _100_ a_24959_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5125 a_27353_8751# tdc1.w_ring_int_norsz[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5128 VPWR a_22603_13103# a_22771_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5129 _026_ a_16135_3311# a_16385_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X5130 tdc0.w_ring_buf[4] a_20727_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5131 VPWR net34 a_24131_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5133 VGND a_17739_7882# tdc1.w_ring_buf[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5134 a_12575_10749# a_11711_10383# a_12318_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5135 VGND a_22603_13103# a_22771_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5136 tdc0.w_ring_norsz[25] net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5138 a_16913_756# ui_in[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5139 tdc1.r_ring_ctr[10] a_17935_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X5140 a_27769_5108# tdc1.w_dly_stop[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5141 VPWR a_28291_6549# a_28207_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5142 a_24021_7369# tdc1.w_ring_norsz[3] a_23937_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5143 a_12977_8041# a_11987_7669# a_12851_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5144 VGND a_15543_7895# _118_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5145 a_12245_10749# a_11711_10383# a_12150_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5147 VPWR net7 a_19071_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5148 VPWR a_13620_9269# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5150 VGND a_24903_10927# a_25071_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5151 VPWR net34 a_23487_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5152 VGND a_22811_3615# tdc1.r_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5153 a_12341_7663# tdc1.w_ring_buf[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5154 a_15373_7485# a_14839_7119# a_15278_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5155 a_15525_4943# a_15481_5185# a_15359_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5157 a_20065_11471# a_19899_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5158 VGND tdc0.w_ring_norsz[22] tdc0.w_ring_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5159 tdc0.w_ring_norsz[30] tdc0.w_ring_norsz[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5160 a_24201_13481# a_23211_13109# a_24075_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5161 VPWR a_9247_14165# a_9163_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5162 VPWR _069_ a_15105_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5163 VPWR a_9282_13077# a_9209_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5164 a_23818_13077# a_23650_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5165 a_18781_6575# tdc1.w_ring_buf[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5166 a_5507_6005# tdc1.r_ring_ctr[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X5167 VPWR a_8327_8725# a_8243_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5168 a_20635_4512# tdc1.r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5169 a_4425_8757# a_4259_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5170 VPWR a_22289_3285# a_22179_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5171 a_22654_10383# a_22339_10535# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5172 VGND net3 _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5173 tdc1.w_ring_norsz[22] net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5175 VPWR a_14767_10901# a_14683_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5177 a_17095_13799# a_17191_13621# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5178 a_9765_10927# tdc0.w_ring_buf[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5179 VGND tdc0.w_ring_int_norsz[28] tdc0.w_ring_norsz[28] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5180 a_23650_13103# a_23377_13109# a_23565_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5182 tdc1.w_ring_buf[0] a_5547_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5183 a_30101_9071# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X5184 a_7201_4097# a_6983_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5185 VPWR _166_ a_22649_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5186 tdc1.w_ring_buf[11] a_27903_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5187 a_22603_13103# a_21739_13109# a_22346_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5188 VGND a_14158_13759# a_14116_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5190 a_19034_6549# a_18866_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5191 VGND _042_ a_18193_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5193 tdc1.r_dly_store_ring[10] a_27647_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5195 VPWR a_4533_14977# a_4423_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5199 a_22273_13103# a_21739_13109# a_22178_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5200 _111_ a_20065_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X5201 VPWR tdc0.r_ring_ctr[3] a_20083_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X5203 a_13243_5705# net30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5204 VPWR _064_ a_14059_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X5205 a_10735_14013# a_10037_13647# a_10478_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5206 VGND _056_ a_14145_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5208 VPWR tdc1.r_ring_ctr[4] a_16217_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5210 a_8849_6575# net76 tdc1.w_ring_int_norsz[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
R64 tdc1.g_ring3[26].stg01_71.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5211 tdc1.r_dly_store_ring[5] a_17711_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5212 VPWR a_16463_12533# net38 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5213 a_8197_7663# a_7663_7669# a_8102_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5214 a_7551_4399# a_6927_4405# a_7443_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5215 VGND a_16163_6397# a_16331_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5216 a_17470_5461# a_17302_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5217 a_12337_4405# a_12171_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5218 a_12226_9407# a_12058_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5219 VGND a_24646_10901# a_24604_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5221 VGND a_8695_7637# a_8653_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5222 VPWR tdc1.r_ring_ctr[14] a_5507_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X5223 a_12318_10495# a_12150_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5224 a_20571_12925# a_19789_12559# a_20487_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5225 a_12226_9407# a_12058_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5226 a_17543_9661# a_16845_9295# a_17286_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5228 VGND tdc0.r_ring_ctr[0] _000_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5229 a_18149_14165# a_17931_14569# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5230 VPWR a_12318_10495# a_12245_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5232 a_16573_9839# tdc0.w_ring_buf[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5233 VPWR a_4420_6031# a_4595_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5234 VGND net28 a_7663_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5235 VGND a_12231_2741# a_12165_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5236 VGND tdc0.w_ring_int_norsz[5] tdc0.w_ring_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5237 _154_ a_15115_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5238 a_22270_5487# a_21997_5493# a_22185_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5239 VGND tdc0.w_ring_norsz[2] tdc0.w_ring_int_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5240 VGND a_15703_7485# a_15871_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5241 a_12875_14709# a_12700_14735# a_13054_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5242 a_18593_6581# a_18427_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5243 a_5985_13647# a_4995_13647# a_5859_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5244 a_26597_12021# a_26431_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5245 VPWR tdc0.r_ring_ctr[2] a_20727_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5247 VPWR tdc0.w_ring_norsz[22] a_10975_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5248 a_12667_5309# a_11803_4943# a_12410_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5249 VGND a_13882_14165# a_13840_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5252 a_22347_15657# a_21997_15285# a_22252_15645# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5253 VPWR _195_ _036_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5254 a_4595_4917# a_4420_4943# a_4774_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5257 tdc1.r_dly_store_ring[17] a_25163_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5258 VPWR _068_ a_10975_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5259 a_22086_14013# a_21813_13647# a_22001_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5260 a_9466_8319# a_9298_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5261 a_16845_4405# a_16679_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5262 a_28989_8751# a_28455_8757# a_28894_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5264 a_9715_6397# a_8933_6031# a_9631_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5265 a_12959_5719# a_13243_5705# a_13178_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5268 a_16135_3311# _166_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5269 VPWR net31 a_21831_5493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5270 VPWR tdc1.w_ring_int_norsz[16] a_5823_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5271 a_19153_6281# net19 tdc1.w_ring_norsz[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5272 a_17739_8970# tdc1.w_ring_norsz[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5273 a_13073_16073# tdc0.r_ring_ctr[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5274 VPWR a_6855_6549# a_6771_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5276 tdc1.w_ring_int_norsz[1] net40 a_22665_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5277 VPWR a_15687_15823# _015_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X5278 a_25777_6575# net40 tdc1.w_ring_int_norsz[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5279 a_20889_6895# tdc1.r_dly_store_ring[4] a_20451_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5280 a_7548_3855# a_6633_3855# a_7201_4097# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5281 a_12139_4007# tdc1.r_ring_ctr[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X5282 tdc0.w_ring_int_norsz[23] net50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5283 tdc0.w_ring_int_norsz[30] net57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5284 VGND a_14155_4917# _179_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X5286 uo_out[6] a_11792_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5288 a_17923_12234# tdc0.w_ring_norsz[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5289 VPWR a_22346_13077# a_22273_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R65 tdc1.g_ring3[18].stg01_63.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5290 tdc0.w_dly_stop[5] a_3155_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5291 VGND _054_ a_8901_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5292 a_16845_14985# tdc0.r_ring_ctr[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5293 a_25305_8041# a_24315_7669# a_25179_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5294 a_19379_7983# _064_ a_19275_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X5295 _196_ a_8399_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5296 a_10946_9295# _134_ a_10124_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5298 a_19127_4777# a_18777_4405# a_19032_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5299 a_9379_3615# a_9204_3689# a_9558_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5300 a_9447_5309# a_8749_4943# a_9190_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5301 a_6373_5193# _181_ a_6291_5193# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5302 a_12139_4007# tdc1.r_ring_ctr[4] a_12313_3883# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5304 VGND tdc0.r_ring_ctr[2] _140_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5305 a_14627_4765# _175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X5306 a_12040_14735# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5307 a_14649_6281# net14 a_14565_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5308 tdc1.w_ring_buf[14] a_18151_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5309 VPWR tdc0.r_ring_ctr[7] a_9008_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X5310 a_3668_7119# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5311 VGND a_4279_9563# a_4237_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5312 a_16385_9845# a_16219_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5314 a_5534_4399# _182_ a_5231_4631# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X5315 a_13629_14191# tdc0.r_ring_ctr[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5317 a_14829_4765# tdc1.r_ring_ctr[9] a_14723_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X5319 a_14059_8983# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.34 w=0.42 l=0.15
X5320 a_15769_15823# _153_ a_15687_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5321 a_17119_4221# a_16495_3855# a_17011_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5322 VGND tdc1.w_ring_norsz[9] tdc1.w_ring_norsz[25] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5323 VGND a_24462_14847# a_24420_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5324 a_14155_4917# tdc1.r_ring_ctr[8] a_14553_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X5325 tdc1.w_ring_int_norsz[20] net65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5326 VGND tdc1.r_ring_ctr[7] a_9897_4737# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X5327 VGND a_21327_7895# tdc1.r_dly_store_ring[18] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5329 a_8753_7119# tdc1.w_ring_buf[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5330 VPWR tdc0.w_ring_norsz[28] a_18151_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5331 a_20261_8029# a_19991_7663# a_20157_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5332 a_24683_13647# _077_ a_24861_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5334 a_11613_12559# tdc0.r_dly_store_ctr[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X5335 a_12610_4399# a_12171_4405# a_12525_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5336 a_18169_10137# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5338 a_14267_16189# _040_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5340 VPWR _189_ a_14008_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5341 a_28526_7663# a_28087_7669# a_28441_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5342 a_5871_11146# tdc0.w_ring_norsz[31] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5343 VGND net19 tdc1.w_ring_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5344 VPWR a_10975_8751# _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5345 tdc0.w_dly_stop[2] a_2603_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5346 a_16266_14013# a_15189_13647# a_16104_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5347 net34 a_24276_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5348 a_4985_12015# net20 tdc0.w_ring_norsz[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5349 a_19587_3689# a_19237_3317# a_19492_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5350 VGND net60 tdc1.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5352 _049_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5353 VGND _135_ a_10977_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5354 a_19867_4703# a_19692_4777# a_20046_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5355 tdc1.w_ring_int_norsz[17] net62 a_7393_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5357 net2 a_855_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5358 VGND a_17751_3829# a_17685_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5359 VGND net36 a_28087_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5360 a_3597_10383# a_3431_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5361 VPWR net7 a_3247_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5364 a_24803_15101# a_24021_14735# a_24719_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5365 a_15207_10927# _074_ a_15289_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5366 tdc0.w_ring_buf[16] a_4627_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5367 VGND _086_ a_6248_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X5368 a_7902_3855# _055_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5370 a_11967_16367# a_11343_16373# a_11859_16745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5372 VGND a_17323_8759# net31 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5374 VPWR tdc0.r_ring_ctr[15] a_3337_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5375 VPWR tdc0.w_ring_norsz[28] a_17405_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5376 VPWR _195_ _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5377 a_27411_7093# tdc1.w_dly_stop[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X5378 a_7897_7284# tdc1.w_ring_norsz[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5379 a_14415_13103# a_13717_13109# a_14158_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5380 VGND a_17567_15797# a_17501_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5381 a_17273_3855# a_17229_4097# a_17107_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5383 VPWR a_9924_14165# net29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5385 a_29181_9545# _072_ a_29035_9447# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X5386 _043_ net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5387 a_18671_14495# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5388 VPWR tdc0.w_ring_norsz[20] a_22843_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5389 tdc1.w_ring_norsz[11] net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5390 VPWR net3 a_9503_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5391 _182_ tdc1.r_ring_ctr[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5392 a_22511_14013# a_21813_13647# a_22254_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5393 a_14293_6281# tdc1.w_ring_norsz[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5394 a_17037_10927# net48 tdc0.w_ring_int_norsz[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5395 _047_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5396 VPWR net34 a_28455_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5397 _187_ a_12815_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5398 a_14090_9295# _194_ a_13620_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5399 a_19235_4399# a_18611_4405# a_19127_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5400 VPWR a_11792_12015# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5401 a_6704_14557# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5403 VPWR tdc0.r_ring_ctr[1] a_19973_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5405 tdc1.w_ring_buf[31] a_7295_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5406 a_13633_10633# tdc0.r_dly_store_ring[8] a_13551_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5408 _095_ a_21279_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5410 a_13201_5487# a_12863_5719# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5414 a_4073_6273# a_3855_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5415 a_10241_7779# _132_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5416 tdc0.w_ring_norsz[9] net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5419 a_9665_13481# a_8675_13109# a_9539_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5420 VPWR a_17100_14165# net32 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5421 tdc0.r_ring_ctr[9] a_17567_15797# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X5422 a_13714_6575# a_13441_6581# a_13629_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5423 a_22167_3689# a_21721_3317# a_22071_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5424 a_10275_10927# a_9577_10933# a_10018_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5425 a_26506_11721# _093_ a_26420_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5427 VPWR tdc1.r_ring_ctr[0] a_20817_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5428 a_11795_6691# _129_ a_11713_6691# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5429 VPWR _184_ a_2769_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5432 a_12736_4777# a_12337_4405# a_12610_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5434 a_20083_14735# tdc0.r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5435 tdc1.w_ring_norsz[28] tdc1.w_ring_int_norsz[28] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5436 a_4328_7119# a_3247_7119# a_3981_7361# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5437 a_28652_8041# a_28253_7669# a_28526_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5438 a_18991_8207# _080_ a_18884_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X5439 a_18243_9071# _065_ a_18243_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5440 VGND a_6671_10651# a_6629_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5441 VGND tdc1.w_ring_int_norsz[6] tdc1.w_ring_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5442 a_12897_8751# tdc1.r_dly_store_ring[16] a_12815_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5444 a_19695_3311# a_19071_3317# a_19587_3689# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5445 a_3024_8725# net26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5446 tdc0.w_ring_norsz[4] tdc0.w_ring_norsz[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5447 VPWR a_12835_5211# a_12751_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5448 VPWR a_19066_7895# _128_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X5449 VGND _067_ a_25933_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.266 pd=2.12 as=0.091 ps=0.93 w=0.65 l=0.15
X5450 VPWR tdc1.r_ring_ctr[1] a_20985_3017# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5451 VGND tdc0.w_ring_buf[27] a_27413_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5453 _008_ _140_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5454 _044_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5455 VGND net64 tdc1.w_ring_int_norsz[19] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5456 a_12397_14735# a_12353_14977# a_12231_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5457 a_7737_13103# a_7203_13109# a_7642_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5458 a_26145_7369# net73 tdc1.w_ring_int_norsz[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5460 tdc0.r_dly_store_ring[16] a_5935_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5461 a_3763_12559# a_3247_12559# a_3668_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5463 a_21998_6575# _108_ a_21912_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5464 a_22543_9295# _080_ a_22447_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.107 ps=0.98 w=0.65 l=0.15
X5465 a_25409_12015# _086_ a_25327_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5467 a_7699_6397# a_7001_6031# a_7442_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5468 VGND net15 _061_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5469 tdc1.w_ring_buf[3] a_24223_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5471 a_14089_10927# tdc0.w_ring_buf[21] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5472 a_8822_14165# a_8654_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5473 VGND tdc0.w_ring_norsz[27] a_25971_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5476 a_6704_14557# _004_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5477 a_6545_12559# tdc0.r_ring_ctr[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5478 a_17283_14709# net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X5479 a_3789_13647# _158_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5480 VPWR tdc1.w_ring_norsz[2] a_23845_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5482 VPWR a_5055_14709# tdc0.r_ring_ctr[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5484 VGND a_6980_4917# net7 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5485 a_13991_3311# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5486 VGND tdc1.r_dly_store_ctr[8] a_13921_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X5487 VPWR a_11067_4399# _175_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5488 a_18087_12925# a_17305_12559# a_18003_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5490 tdc0.w_ring_norsz[2] net22 a_22653_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5491 VPWR net36 a_29007_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5492 a_8654_14191# a_8381_14197# a_8569_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5493 VPWR _166_ a_11115_4007# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5494 a_10505_3311# _172_ _028_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5495 tdc1.w_ring_norsz[1] net17 a_23021_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5497 VPWR tdc0.w_ring_norsz[23] a_7755_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5498 a_26785_12015# tdc0.w_ring_buf[18] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5499 VGND _070_ a_18335_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5500 a_5449_4719# _183_ a_5231_4631# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
R66 VGND uio_out[1] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5502 _135_ a_10087_10411# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X5503 a_14909_8751# _065_ a_14655_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5504 VGND _090_ a_24683_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5505 VPWR a_2287_10901# tdc0.r_ring_ctr[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X5506 a_20353_13423# tdc0.r_dly_store_ctr[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X5507 a_24137_7663# tdc1.w_ring_norsz[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5508 a_4420_6031# a_3505_6031# a_4073_6273# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5510 a_15105_13103# tdc0.r_dly_store_ring[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5511 tdc1.w_ring_int_norsz[16] net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5512 VPWR tdc0.w_ring_norsz[26] a_19255_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5513 net31 a_17323_8759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X5514 VGND a_25807_5461# a_25765_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5516 VPWR tdc1.w_ring_norsz[10] a_26789_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5517 tdc0.w_ring_int_norsz[11] tdc0.w_ring_norsz[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5518 VGND a_11582_13077# a_11540_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
R67 VGND net56 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5519 VGND net30 a_12171_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5520 VGND a_8822_14165# a_8780_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5522 VGND net25 a_10217_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X5523 VGND a_18003_12925# a_18171_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R68 net74 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5524 VPWR a_10443_10901# a_10359_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5525 VGND a_8183_4703# a_8117_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5526 a_12862_15101# a_11785_14735# a_12700_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5527 VPWR net9 a_11343_16373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5528 VGND a_28123_6575# a_28291_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5529 a_18593_10933# a_18427_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5531 a_11839_13103# a_11141_13109# a_11582_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5532 a_26781_9845# a_26615_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5533 a_18501_7663# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X5534 VPWR a_29119_9813# a_29035_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5535 a_9029_13103# tdc0.w_ring_buf[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5536 VGND tdc0.w_ring_norsz[9] tdc0.w_ring_norsz[25] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5537 a_11414_13103# a_10975_13109# a_11329_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5539 a_19310_13759# a_19142_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5540 a_5342_11837# a_5069_11471# a_5257_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5541 VPWR a_14448_3689# a_14623_3615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5543 VGND net7 a_6927_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5544 _017_ _177_ a_15649_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X5545 a_17869_2767# a_16679_2767# a_17760_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5547 a_18671_14495# a_18496_14569# a_18850_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5548 _134_ a_10241_7779# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X5549 a_19433_10205# a_19163_9839# a_19329_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5550 tdc1.r_dly_store_ring[25] a_30039_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5551 a_9272_16189# a_9058_16189# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X5552 a_3686_9661# a_3413_9295# a_3601_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5554 VPWR tdc0.r_ring_ctr[0] a_18029_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5555 a_18877_8457# _081_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X5556 a_13599_6196# tdc1.w_ring_norsz[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5558 VPWR a_14011_9839# _075_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5559 tdc0.w_ring_norsz[6] tdc0.w_ring_int_norsz[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5560 VGND net21 tdc0.w_ring_norsz[30] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5561 a_8747_3311# _054_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5562 a_13990_13103# a_13551_13109# a_13905_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5563 VPWR a_19567_10749# a_19735_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5564 VGND a_20083_8751# _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5565 a_21825_15823# a_20635_15823# a_21716_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5567 a_6449_14197# a_6283_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5568 VGND a_20230_12671# a_20188_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5569 VGND net31 a_16863_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5570 a_25731_13103# a_24867_13109# a_25474_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5571 _133_ a_9595_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5572 a_20319_13621# a_20610_13921# a_20561_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5573 a_28621_8757# a_28455_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5575 tdc1.r_dly_store_ring[4] a_21115_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5576 VPWR net8 a_14747_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5577 a_15504_9295# _122_ a_15333_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5578 net5 a_16219_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5579 a_16573_9839# tdc0.w_ring_buf[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5580 tdc0.w_ring_norsz[28] tdc0.w_ring_norsz[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5581 VGND _084_ a_25182_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5584 a_5703_6031# _181_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X5585 VGND a_14800_6549# net16 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5587 VPWR tdc0.w_ring_int_norsz[16] a_5069_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5588 a_22304_13481# a_21905_13109# a_22178_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5589 VGND a_4038_10495# a_3996_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5590 VPWR net29 a_9411_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5591 VGND net29 a_11711_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5593 _012_ _148_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5594 VPWR a_27411_7093# net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5595 VGND a_27479_9839# a_27647_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5596 VPWR a_17375_7637# net39 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5597 VPWR net29 a_14103_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
R69 VGND net60 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5598 VGND tdc1.w_ring_norsz[1] tdc1.w_ring_norsz[17] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5600 a_5905_6031# tdc1.r_ring_ctr[13] a_5799_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X5601 VPWR a_17923_12234# tdc0.w_ring_buf[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R70 VPWR tdc1.g_ring3[24].stg01_69.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5602 a_21545_10383# _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X5603 VGND net11 tdc0.w_ring_int_norsz[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5606 VGND a_5123_8751# a_5291_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5607 VGND net20 _045_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5608 VPWR a_13882_6549# a_13809_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5609 VGND a_21223_5309# a_21391_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5610 _166_ a_21923_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X5611 a_20169_9295# a_19899_9295# a_20065_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5612 tdc0.w_ring_norsz[24] tdc0.w_ring_int_norsz[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5613 a_12077_16341# a_11859_16745# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5614 a_25182_10383# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X5615 VPWR a_13735_12559# net23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5616 VPWR tdc0.r_ring_ctr[12] a_4219_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X5617 a_12981_6575# tdc1.w_ring_norsz[30] a_12897_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5619 a_20338_11837# a_19899_11471# a_20253_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5620 a_20487_12925# a_19623_12559# a_20230_12671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5622 a_24131_6281# _077_ a_24213_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5623 a_22925_6575# net17 tdc1.w_ring_norsz[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5624 a_26247_6281# _075_ a_26329_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5625 VGND a_10699_14735# _152_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5626 VPWR net32 a_18703_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5627 a_14415_14013# a_13551_13647# a_14158_13759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5628 VPWR a_4111_9661# a_4279_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5629 a_20445_4105# tdc1.r_ring_ctr[2] _163_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5630 a_9459_8970# tdc1.w_ring_norsz[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5632 VGND _185_ _021_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5633 VGND net6 a_14794_9922# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5634 a_11435_12559# _075_ a_11613_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5635 a_13035_4399# a_12171_4405# a_12778_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5636 VGND net7 a_3247_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5637 tdc0.w_ring_buf[12] a_19899_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5638 a_20157_12925# a_19623_12559# a_20062_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5640 tdc1.w_ring_buf[20] a_22935_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5641 VPWR net7 a_21555_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5642 _085_ _084_ a_24591_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5643 VGND a_9503_9295# _086_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X5644 VGND tdc0.w_ring_int_norsz[29] tdc0.w_ring_norsz[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5645 a_9121_6031# tdc1.w_ring_buf[30] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5647 a_11923_13103# a_11141_13109# a_11839_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5648 a_14085_14013# a_13551_13647# a_13990_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5649 a_8228_10217# a_7829_9845# a_8102_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5652 VPWR a_11087_5211# a_11003_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5653 tdc1.r_dly_store_ctr[3] a_24519_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5654 a_12815_8751# _067_ a_12897_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5655 a_13551_10633# _071_ a_13633_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5657 a_23684_10217# a_23285_9845# a_23558_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5658 a_5635_5193# tdc1.r_ring_ctr[13] a_5417_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5660 VPWR a_17935_2741# tdc1.r_ring_ctr[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5661 a_14710_11989# a_14542_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5662 a_14158_13759# a_13990_14013# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5663 a_10872_7119# tdc1.r_dly_store_ring[31] a_10569_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X5664 VGND _089_ a_21095_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.172 ps=1.83 w=0.65 l=0.15
X5665 a_12529_13103# tdc0.r_dly_store_ctr[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5667 a_19291_6575# a_18593_6581# a_19034_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5669 a_17118_9661# a_16679_9295# a_17033_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5670 tdc0.r_dly_store_ctr[3] a_24887_15003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5672 VGND _053_ a_11753_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5673 a_24462_11989# a_24294_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5674 VGND a_17555_7284# tdc1.w_ring_buf[21] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5675 VGND tdc0.w_ring_norsz[2] tdc0.w_ring_norsz[18] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5677 VGND a_2511_14191# net28 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5678 VPWR a_9551_15511# _148_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X5679 VPWR a_21511_9447# _112_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X5680 a_24903_10927# a_24039_10933# a_24646_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5681 a_23285_11721# tdc0.w_ring_norsz[3] a_23201_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5685 VGND net16 tdc1.w_ring_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5686 _004_ a_6364_14985# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.327 ps=1.65 w=1 l=0.15
R71 VGND net75 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5688 a_6799_14569# a_6283_14197# a_6704_14557# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5689 a_2519_7369# _184_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5690 tdc0.r_dly_store_ring[7] a_5291_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5693 a_4617_13647# tdc0.r_ring_ctr[13] a_4511_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X5694 VPWR _079_ a_25071_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5695 a_8270_9813# a_8102_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5696 a_24573_10927# a_24039_10933# a_24478_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5697 VPWR _047_ a_2287_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5698 VGND _065_ _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5699 a_14159_15823# a_13809_15823# a_14064_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5701 a_28538_12292# a_28338_12137# a_28687_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5702 VPWR _180_ a_5534_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X5703 a_7661_4373# a_7443_4777# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5704 tdc0.w_ring_buf[3] a_23763_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5705 _185_ tdc1.r_ring_ctr[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.176 ps=1.84 w=0.65 l=0.15
X5708 VGND _081_ a_22543_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X5709 a_28526_9839# a_28087_9845# a_28441_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5711 a_17100_4765# _017_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5712 a_5437_12015# tdc0.w_ring_norsz[16] a_5353_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5713 tdc1.r_dly_store_ctr[9] a_22863_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5714 _153_ tdc0.r_ring_ctr[8] a_15753_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5715 a_8378_12015# a_7939_12021# a_8293_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5716 a_17195_2767# a_16845_2767# a_17100_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5718 VPWR net33 a_21279_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5719 _192_ a_13551_10633# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5720 a_2963_10901# a_2768_11043# a_3273_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X5721 VPWR a_7201_4097# a_7091_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5723 VPWR a_17083_9839# a_17251_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5724 a_15823_14735# _152_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X5726 VPWR a_14158_13759# a_14085_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5728 a_15543_7895# tdc1.r_dly_store_ring[13] a_15717_8001# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5729 _167_ _164_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5730 tdc1.w_ring_norsz[0] net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5731 tdc0.r_dly_store_ctr[2] a_25899_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5733 tdc0.r_dly_store_ctr[11] a_22679_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5734 a_9022_5309# a_8583_4943# a_8937_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5736 a_18866_6575# a_18593_6581# a_18781_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5737 a_7079_3855# a_6633_3855# a_6983_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5738 tdc1.r_dly_store_ring[3] a_25347_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5739 VPWR a_3854_9407# a_3781_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5740 a_12276_10383# a_11877_10383# a_12150_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5741 VGND _037_ a_12397_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5742 tdc1.r_ring_ctr[13] a_4595_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X5743 a_19567_5309# a_18869_4943# a_19310_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5744 VPWR tdc1.w_ring_norsz[20] a_22935_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5745 VPWR net29 a_13551_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5747 VGND net36 a_29007_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5748 VGND _067_ a_11873_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X5749 a_20437_6031# tdc1.w_ring_buf[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5751 VGND a_19034_10901# a_18992_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5752 VPWR a_14427_12724# tdc0.w_ring_buf[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5753 VGND tdc1.w_ring_norsz[24] tdc1.w_ring_norsz[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5754 a_24719_15101# a_23855_14735# a_24462_14847# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5756 a_15289_10927# tdc0.r_dly_store_ctr[5] a_15207_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5757 a_17554_16189# a_16477_15823# a_17392_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5759 tdc1.w_ring_norsz[17] net17 a_23021_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5761 a_17010_13077# a_16842_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5762 a_17244_9295# a_16845_9295# a_17118_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5763 VPWR a_5507_6005# _184_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X5766 _033_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5767 a_14427_12724# tdc0.w_ring_norsz[29] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5768 VGND a_17935_4703# a_17869_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5770 tdc0.r_dly_store_ring[11] a_22771_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5771 VPWR _086_ a_5773_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X5772 VPWR net30 a_10055_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5773 VPWR a_10735_14013# a_10903_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5775 a_24389_15101# a_23855_14735# a_24294_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5776 a_15654_14191# _155_ a_15351_14423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X5777 a_20811_9955# _112_ a_20729_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5778 tdc0.r_dly_store_ring[11] a_22771_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5779 a_20809_14735# tdc0.r_ring_ctr[0] a_20727_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5781 a_22719_10357# net35 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5782 VPWR a_24646_10901# a_24573_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5783 VPWR a_11792_12015# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5785 VPWR a_5055_14709# a_5042_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5786 a_19057_13647# tdc0.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5787 a_28253_7669# a_28087_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5788 _024_ _164_ a_20825_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5789 a_25731_4221# a_25033_3855# a_25474_3967# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5790 VPWR net4 a_16587_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X5791 tdc0.w_ring_buf[22] a_10975_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5792 a_24462_14847# a_24294_15101# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5794 a_17457_4765# a_17413_4373# a_17291_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5795 a_16301_7663# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5796 VGND tdc0.w_ring_int_norsz[8] tdc0.w_ring_norsz[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5797 VGND a_20327_3615# tdc1.r_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5798 _006_ a_3255_11721# a_3505_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X5799 VPWR _152_ a_15115_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5801 VPWR a_22679_13915# a_22595_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5802 a_23947_12809# _072_ a_24029_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5803 a_10395_7779# _132_ a_10323_7779# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5805 _086_ a_9503_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X5806 a_22903_14709# a_22728_14735# a_23082_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5808 VPWR a_13882_14165# a_13809_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5809 VPWR a_24276_9269# net34 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5810 _097_ a_22257_9545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.112 ps=0.995 w=0.65 l=0.15
X5811 _031_ _176_ a_15281_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X5812 VGND a_16003_4917# a_15937_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5813 a_21361_4765# tdc1.r_ring_ctr[0] a_21279_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X5814 VGND a_8270_7637# a_8228_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5815 tdc0.w_ring_norsz[6] net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5816 a_16658_9839# a_16385_9845# a_16573_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5817 a_17303_3133# a_16679_2767# a_17195_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5818 VGND a_27951_12247# tdc0.r_dly_store_ring[26] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5820 VGND _048_ a_19849_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5821 VGND a_15504_9295# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X5822 VGND a_25639_5487# a_25807_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5823 VGND a_16463_12533# net38 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5825 VPWR a_14415_13103# a_14583_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5826 a_17739_8970# tdc1.w_ring_norsz[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5827 a_10147_9839# _076_ a_10229_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5829 a_30021_7983# _072_ a_29587_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5830 VGND tdc1.w_ring_norsz[17] tdc1.w_ring_int_norsz[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5831 a_3781_9661# a_3247_9295# a_3686_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5832 VPWR _069_ a_10229_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5833 VPWR a_13203_4373# a_13119_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5834 a_11333_10927# net21 tdc0.w_ring_norsz[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5835 VGND a_14415_13103# a_14583_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5836 a_21716_15823# a_20801_15823# a_21369_16065# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5839 a_9204_3689# a_8289_3317# a_8857_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5840 VGND net38 tdc1.w_ring_int_norsz[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5841 a_7768_13481# a_7369_13109# a_7642_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5842 a_9148_4943# a_8749_4943# a_9022_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5844 a_12863_5719# a_12959_5719# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5846 VGND a_8695_9813# a_8653_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5848 a_4219_13621# _158_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X5849 VGND net22 tdc0.w_ring_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5850 VGND tdc0.r_ring_ctr[12] a_3439_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5851 VPWR a_2963_10901# a_2894_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X5852 a_10225_13647# tdc0.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
R72 tt_um_hpretl_tt06_tdc_v2_82.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5853 a_23742_5487# a_23469_5493# a_23657_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5854 a_5510_11583# a_5342_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5857 VPWR net22 a_18703_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5858 a_26995_11305# a_26859_11145# a_26575_11159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5859 a_14008_9545# _083_ a_13620_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X5860 a_22068_14735# _008_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5862 VGND _061_ a_4117_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5863 tdc1.r_dly_store_ring[4] a_21115_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5864 VGND a_5767_11837# a_5935_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5865 a_21056_15823# _007_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5866 a_28731_6575# _072_ a_28909_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5867 VGND tdc1.w_ring_int_norsz[12] tdc1.w_ring_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5868 VGND tdc0.w_ring_norsz[12] tdc0.w_ring_int_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5869 a_25432_14569# a_25033_14197# a_25306_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5871 a_19959_15797# _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5872 VGND a_17286_9407# a_17244_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5873 VGND a_18169_10137# a_18103_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5874 a_6587_10749# a_5805_10383# a_6503_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5875 a_6817_15285# a_6651_15285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5876 a_24385_14569# a_23395_14197# a_24259_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5877 a_4613_9839# tdc0.w_ring_buf[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5880 a_24995_8751# a_24297_8757# a_24738_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5881 a_7461_12015# tdc0.w_ring_norsz[15] a_7377_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5882 _196_ a_8399_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5883 VGND a_22811_3615# a_22745_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5884 a_17375_7637# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X5885 a_13809_15823# a_13643_15823# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5889 VGND _186_ a_13553_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5890 _041_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5891 _162_ tdc0.r_ring_ctr[14] a_3789_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.162 ps=1.33 w=1 l=0.15
X5892 VPWR a_7907_15583# a_7894_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5893 _622_.X a_2840_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5894 VGND _155_ a_15569_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X5895 VGND tdc1.w_ring_norsz[24] tdc1.w_ring_int_norsz[25] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5896 tdc0.w_ring_norsz[1] tdc0.w_ring_norsz[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5897 a_17881_7369# tdc1.w_ring_norsz[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5898 VGND tdc0.w_ring_norsz[25] a_17875_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5899 a_14415_13103# a_13551_13109# a_14158_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
R73 tdc0.g_ring3[30].stg01_57.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
R74 tt_um_hpretl_tt06_tdc_v2_88.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5902 a_4073_5185# a_3855_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5903 a_22333_3677# a_22289_3285# a_22167_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5904 VGND tdc1.w_ring_norsz[11] a_27903_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5906 a_24683_10159# _090_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5907 _070_ a_16771_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X5908 a_14085_13103# a_13551_13109# a_13990_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5909 VGND net32 a_18703_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5910 VPWR tdc0.r_ring_ctr[7] a_9167_14763# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5911 _061_ net15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5912 VPWR a_9379_3615# a_9366_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5913 VPWR a_10919_5309# a_11087_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5914 VGND net32 a_16403_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5915 _151_ a_10239_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5916 VGND _125_ a_11623_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5917 VPWR a_12056_2767# a_12231_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5920 a_18199_9878# tdc1.r_dly_store_ring[5] a_17740_10071# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X5921 tdc0.w_ring_buf[24] a_9135_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5922 tdc1.w_ring_buf[14] a_18151_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5923 a_16279_13621# a_16104_13647# a_16458_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5924 a_15649_4399# tdc1.r_ring_ctr[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5925 a_22438_5461# a_22270_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5926 a_26479_11159# a_26575_11159# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5927 VGND tdc0.w_ring_int_norsz[13] tdc0.w_ring_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5929 a_17858_14013# a_17611_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5930 a_17100_2767# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5931 tdc1.r_dly_store_ctr[12] a_20471_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5935 a_17313_10927# net39 tdc0.w_ring_int_norsz[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5936 a_23021_15657# a_21831_15285# a_22912_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5938 VGND net32 a_18427_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5939 VGND tdc1.w_ring_int_norsz[16] tdc1.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5940 a_24995_8751# a_24131_8757# a_24738_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5942 VGND _179_ a_12621_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5945 tdc0.w_dly_stop[2] a_2603_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5946 a_14158_13759# a_13990_14013# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5947 a_27413_11305# a_26859_11145# a_27066_11204# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X5948 VPWR net9 a_6651_15285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5949 VGND a_9190_5055# a_9148_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5950 a_22701_3855# a_22657_4097# a_22535_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5951 a_18981_12015# tdc0.w_ring_int_norsz[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5953 VPWR tdc1.w_ring_norsz[16] a_7111_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5954 a_4425_9845# a_4259_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5955 VPWR net25 a_13633_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5957 VGND a_29319_8751# a_29487_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5958 tdc1.r_dly_store_ring[13] a_14307_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5959 a_29997_7119# a_29007_7119# a_29871_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5961 a_13633_7369# _076_ a_13717_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5963 a_23377_13109# a_23211_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5964 a_24941_5493# a_24775_5493# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5965 tdc0.w_ring_buf[16] a_4627_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5966 a_25221_14191# tdc0.r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5969 a_19567_10749# a_18869_10383# a_19310_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5972 a_9647_14709# _156_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X5973 net29 a_9924_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5974 net23 a_13735_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X5975 a_25432_13481# a_25033_13109# a_25306_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R75 VGND uio_oe[7] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5976 VPWR a_8803_12015# a_8971_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5977 a_15444_13647# _002_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5978 a_24477_4777# a_23487_4405# a_24351_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5979 a_4613_8751# tdc1.w_ring_buf[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5980 VGND a_28383_5461# a_28341_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5981 VPWR a_11987_9839# _067_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5983 a_6002_5807# tdc1.r_ring_ctr[12] _185_ VGND sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.106 ps=0.975 w=0.65 l=0.15
X5984 VGND a_8803_12015# a_8971_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5985 VGND net40 tdc0.w_ring_int_norsz[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5987 a_6630_12925# a_6191_12559# a_6545_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5988 VGND tdc0.r_ring_ctr[10] a_16595_14985# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5990 a_5069_12015# net42 a_4985_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5991 VPWR a_14158_13077# a_14085_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5992 a_11035_3543# _168_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X5993 a_21279_4765# tdc1.r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5994 a_11396_2767# _027_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5997 a_7745_12015# net38 tdc0.w_ring_int_norsz[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5998 a_4503_12533# _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6000 VPWR a_18171_8475# a_18087_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6003 a_22093_13103# tdc0.w_ring_buf[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6006 a_9589_10159# tdc0.r_dly_store_ring[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6008 a_12778_16733# _036_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6009 uo_out[0] a_13620_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6010 a_22425_14735# a_22381_14977# a_22259_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6011 VGND a_21707_7881# a_21714_7785# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6012 VPWR a_16826_9813# a_16753_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6014 VPWR tdc1.r_ring_ctr[15] a_2601_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6015 tdc0.w_ring_int_norsz[1] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6017 a_22089_3855# a_21923_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6018 a_7369_13109# a_7203_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6020 _194_ a_5015_9622# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X6021 a_19481_15823# a_19437_16065# a_19315_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6023 a_23561_14197# a_23395_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6025 a_11067_11471# _083_ a_11245_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X6026 a_15701_8457# _065_ a_15283_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6028 VGND tdc1.w_ring_norsz[2] a_21003_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6029 VGND a_22311_8725# a_22269_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6030 tdc0.r_dly_store_ctr[13] a_8235_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6031 a_18961_6575# a_18427_6581# a_18866_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6032 VGND a_5055_14709# a_4989_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X6033 VPWR a_17576_3855# a_17751_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6034 VGND a_8327_8725# a_8285_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6035 tdc0.r_dly_store_ctr[10] a_24427_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6036 VGND a_22438_5461# a_22396_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6038 a_8183_4703# a_8008_4777# a_8362_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6039 a_7661_4373# a_7443_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6040 VGND net29 a_13551_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6041 _152_ a_10699_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X6042 a_14223_6575# a_13441_6581# a_14139_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6043 a_25348_10633# _105_ a_25182_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6044 VGND tdc0.w_ring_int_norsz[27] tdc0.w_ring_norsz[27] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6045 a_19235_4399# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6046 VGND net20 _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6047 VPWR a_10569_7093# _131_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6048 a_4490_7485# a_3413_7119# a_4328_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
R76 tdc0.g_ring1[16].stg02_42.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6049 a_18992_11305# a_18593_10933# a_18866_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6050 _055_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6051 VPWR a_18003_12925# a_18171_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6052 _052_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6053 a_18795_13103# _072_ a_18877_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6054 VPWR tdc1.r_dly_store_ring[29] a_16301_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X6055 VPWR tdc0.w_ring_buf[20] a_23273_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6056 VGND a_6855_6549# a_6813_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6057 tdc0.w_ring_norsz[29] tdc0.w_ring_norsz[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6059 VGND a_28694_9813# a_28652_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6060 VPWR a_23910_5461# a_23837_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6062 tdc0.w_ring_buf[10] a_24775_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6063 VGND tdc0.w_ring_norsz[12] a_19899_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6064 a_19973_15599# tdc0.r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6066 VGND a_8546_11989# a_8504_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6067 _170_ tdc1.r_ring_ctr[4] a_11978_3631# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X6068 a_24002_14165# a_23834_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6070 VPWR a_20503_15253# _143_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6071 a_11509_13103# a_10975_13109# a_11414_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6074 a_27295_12015# a_26597_12021# a_27038_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6075 a_11908_14569# a_11509_14197# a_11782_14191# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6076 a_19268_13647# a_18869_13647# a_19142_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6077 a_10147_13103# _077_ a_10229_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6079 VPWR _121_ a_15333_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X6081 a_3981_7361# a_3763_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6083 a_28809_8751# tdc1.w_ring_buf[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6084 VPWR a_5935_11739# a_5851_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6086 a_14197_10389# _191_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6088 VGND a_24719_15101# a_24887_15003# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6090 a_12725_6031# _075_ a_12291_6183# VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6091 VPWR a_8399_3855# _196_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6092 VPWR net30 a_11987_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6096 VGND a_21914_7940# a_21843_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6097 a_4989_14735# a_3799_14735# a_4880_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6099 a_17317_7369# tdc1.w_ring_norsz[6] a_17233_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6100 a_22890_15101# a_21813_14735# a_22728_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6101 net28 a_2511_14191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X6102 a_17033_9295# tdc1.w_ring_buf[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6103 VGND tdc0.w_ring_norsz[23] a_7755_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6104 VPWR a_23259_7882# tdc1.w_ring_buf[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6105 tdc1.w_ring_norsz[8] net16 a_11705_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6106 a_15719_10357# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6107 tdc1.r_ring_ctr[14] a_4595_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6108 VGND _145_ a_10449_15617# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6109 a_16753_9839# a_16219_9845# a_16658_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6111 VPWR tdc1.r_ring_ctr[8] a_14431_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X6113 a_24343_14191# a_23561_14197# a_24259_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6114 a_21445_8757# a_21279_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6115 a_7461_8757# a_7295_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6116 VGND a_9647_14709# _158_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X6118 VGND a_7442_6143# a_7400_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6119 VGND a_14767_10901# a_14725_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6120 VGND a_14011_9839# _075_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6121 a_9807_8573# a_9025_8207# a_9723_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6122 VPWR a_14431_4373# _178_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X6123 a_16916_3855# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6124 VGND net31 a_16679_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6125 _089_ a_18795_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6127 VPWR net30 a_13275_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6129 a_16309_8867# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X6130 a_22089_3855# a_21923_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6132 VGND a_24427_14165# a_24385_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6133 a_16753_10927# tdc0.w_ring_norsz[5] a_16669_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6134 a_14802_3677# _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6135 a_12587_8372# tdc1.w_ring_norsz[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6136 VGND tdc1.r_ring_ctr[10] a_15399_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6137 _035_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6138 VPWR a_23671_15287# net36 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6139 a_17089_15823# a_17045_16065# a_16923_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6140 tdc0.r_dly_store_ring[15] a_7223_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6141 VGND a_3247_13647# net37 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6142 _053_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6144 VGND tdc1.w_ring_norsz[13] tdc1.w_ring_int_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6145 a_15465_6031# a_15299_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6146 a_27173_9545# tdc1.w_ring_norsz[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6147 VPWR a_12599_16671# a_12586_16367# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6148 VPWR _070_ a_14655_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6149 tdc1.r_ring_ctr[11] a_16003_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6151 VPWR a_22511_14013# a_22679_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6153 a_25033_13109# a_24867_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6154 _058_ net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6155 tdc1.r_dly_store_ring[31] a_9431_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6157 tdc1.w_ring_norsz[9] net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6158 VGND tdc1.w_ring_norsz[28] tdc1.w_ring_int_norsz[29] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6159 net20 a_3399_12275# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X6160 VPWR _143_ a_11343_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X6162 tdc1.w_ring_int_norsz[30] tdc1.w_ring_norsz[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6163 uo_out[7] a_10124_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6164 a_7093_12015# tdc0.w_ring_norsz[31] a_7009_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6165 VGND a_22926_10357# a_22855_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6168 a_17083_9839# a_16385_9845# a_16826_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6169 VPWR a_5043_11146# tdc0.w_ring_buf[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6170 net7 a_6980_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6171 VGND _069_ a_10309_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6172 a_15504_9295# _083_ a_15333_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X6173 VPWR a_21369_16065# a_21259_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6174 VGND tdc0.r_dly_store_ring[12] a_21833_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6175 VGND net35 a_23855_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6176 a_4588_7637# net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6177 a_18605_14569# a_17415_14197# a_18496_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6178 VGND a_23983_9839# a_24151_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6180 a_19057_4943# tdc1.r_ring_ctr[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6181 a_4195_9661# a_3413_9295# a_4111_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6182 _125_ a_11067_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X6185 net5 a_16219_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6186 a_12533_16745# a_11343_16373# a_12424_16745# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6187 _032_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6188 VPWR _071_ a_12539_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6189 VGND _076_ a_9963_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6191 VPWR tdc1.w_ring_norsz[19] a_23569_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6193 _070_ a_16771_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X6194 net9 a_18059_16375# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6195 a_12056_2767# a_10975_2767# a_11709_3009# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6197 a_21157_13647# a_20603_13621# a_20810_13621# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6198 VGND net26 a_8583_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6199 a_9459_8970# tdc1.w_ring_norsz[23] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6200 a_22912_15657# a_21997_15285# a_22565_15253# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6201 a_14951_3855# _176_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X6203 VPWR a_4588_7637# _623_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6205 tdc0.w_ring_norsz[8] tdc0.w_ring_norsz[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6206 uo_out[3] a_25348_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6208 a_19142_5309# a_18703_4943# a_19057_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6209 net19 a_27411_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6210 VGND _050_ a_19389_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6211 VPWR a_3981_7361# a_3871_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6212 VPWR net31 a_17139_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6213 VGND a_12743_10651# a_12701_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6214 a_24075_13103# a_23377_13109# a_23818_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6215 a_19345_4373# a_19127_4777# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6216 a_20810_13621# a_20603_13621# a_20986_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6217 VGND a_12667_5309# a_12835_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6219 VPWR net13 a_7009_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6220 VPWR a_2807_11169# a_2768_11043# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6221 a_24276_9269# net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
R77 tdc1.g_ring3[19].stg01_64.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6223 a_18613_12015# tdc0.w_ring_int_norsz[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6224 a_22912_15657# a_21831_15285# a_22565_15253# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6225 a_21826_6575# _107_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X6226 VGND _109_ a_20729_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6227 a_16827_15823# a_16311_15823# a_16732_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6228 a_24294_12015# a_23855_12021# a_24209_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6229 VPWR a_9631_6397# a_9799_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6231 _084_ net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6233 a_19291_10927# a_18427_10933# a_19034_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6234 VPWR tdc0.w_ring_norsz[4] a_17313_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
R78 VGND uio_out[3] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6236 a_25306_4221# a_24867_3855# a_25221_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
R79 tdc1.g_ring3[30].stg01_75.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6237 a_3668_7119# _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6238 VPWR tdc1.r_ring_ctr[0] a_20445_4105# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X6240 a_22185_5487# tdc1.r_ring_ctr[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6241 VGND _059_ a_15525_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6242 VGND tdc0.w_ring_norsz[21] tdc0.w_ring_int_norsz[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6244 a_18593_6581# a_18427_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6246 VGND _075_ a_24477_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6247 VPWR a_18059_16375# net9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6248 a_22637_13647# a_21647_13647# a_22511_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6249 VGND _067_ a_26593_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6250 tdc1.w_ring_buf[15] a_7571_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6251 _011_ _147_ a_11809_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6252 a_7557_13103# tdc0.r_ring_ctr[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6253 tdc0.w_ring_int_norsz[25] net52 a_12729_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6255 VPWR a_20046_5461# a_19973_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6257 _623_.X a_4588_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
R80 tdc0.g_ring3[16].stg01_43.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6259 net14 a_12539_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6261 VGND net29 a_9411_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6263 VPWR net10 a_16311_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6266 VPWR net35 a_23855_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6268 tdc0.r_dly_store_ring[3] a_25071_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6269 a_20257_13103# _077_ a_20341_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6271 VGND net31 a_21831_5493# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6272 a_27613_6575# tdc1.w_ring_buf[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6273 a_15168_4943# _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6274 VPWR a_19310_13759# a_19237_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6275 a_7377_12015# net21 tdc0.w_ring_norsz[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6276 VGND tdc0.w_ring_norsz[10] a_24775_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6277 a_23926_4399# a_23653_4405# a_23841_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6278 a_10018_11989# a_9850_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6280 VGND a_15335_8181# _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6281 _054_ _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6282 VPWR net27 a_6191_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6283 a_15481_5185# a_15263_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6285 tdc1.r_dly_store_ring[0] a_4279_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6286 VPWR a_10903_13915# a_10819_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6287 a_5236_9295# tdc1.r_dly_store_ring[0] a_5015_9622# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6288 a_13633_10633# tdc0.r_dly_store_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6289 a_20525_4943# a_20359_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6290 VGND tdc0.r_ring_ctr[4] a_10799_16073# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6291 a_5859_14013# a_5161_13647# a_5602_13759# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6292 a_14116_13481# a_13717_13109# a_13990_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6294 a_8933_6031# a_8767_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6295 VGND a_2963_10901# a_2894_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X6296 VGND _174_ a_11067_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X6297 tdc1.r_ring_ctr[9] a_17751_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X6298 a_5434_14013# a_4995_13647# a_5349_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6299 VGND a_26479_11159# tdc0.r_dly_store_ring[27] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6300 VPWR a_28331_12233# a_28338_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6301 a_9531_5309# a_8749_4943# a_9447_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6302 a_19268_4943# a_18869_4943# a_19142_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6303 VGND _124_ a_11623_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6304 a_17576_3855# a_16495_3855# a_17229_4097# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6305 _000_ tdc0.r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6306 a_9924_14165# net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X6307 tdc0.w_ring_buf[20] a_22843_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6308 VGND a_13035_4399# a_13203_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6309 tdc1.r_dly_store_ring[17] a_25163_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6310 a_22212_13647# a_21813_13647# a_22086_14013# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6311 a_19692_4777# a_18611_4405# a_19345_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6312 tdc1.r_dly_store_ring[24] a_12651_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6315 VGND _034_ a_22425_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6316 VGND net19 _059_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6317 a_7649_8751# tdc1.w_ring_buf[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6318 a_19127_4777# a_18611_4405# a_19032_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6319 a_4219_13621# tdc0.r_ring_ctr[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X6320 VGND _165_ a_21923_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X6321 a_20230_12671# a_20062_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6322 a_14703_12724# tdc0.w_ring_norsz[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6323 a_21423_7895# a_21714_7785# a_21665_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6324 a_3413_12559# a_3247_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6325 VGND _032_ a_19481_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6327 VGND a_12851_7663# a_13019_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6328 VGND a_3484_13077# net21 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6329 a_7189_6031# tdc1.r_ring_ctr[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6330 VPWR a_17435_13077# a_17351_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6332 a_7181_10217# a_6191_9845# a_7055_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6334 tdc1.r_dly_store_ctr[1] a_24335_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6335 a_24570_8751# a_24131_8757# a_24485_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6337 VPWR a_14011_9839# _075_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6338 a_24021_12021# a_23855_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6339 a_15197_14735# tdc0.r_ring_ctr[8] a_15115_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6340 tdc0.w_ring_norsz[18] net24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6341 _036_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6342 VPWR a_19034_10901# a_18961_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6343 a_4595_4917# _061_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6344 VGND a_19291_6575# a_19459_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6345 a_25432_3855# a_25033_3855# a_25306_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6346 a_5805_10383# a_5639_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6347 a_4038_10495# a_3870_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6349 tdc0.r_dly_store_ring[14] a_10443_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6350 a_23749_14191# tdc0.r_ring_ctr[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6352 a_23937_7369# net17 tdc1.w_ring_norsz[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6355 a_9953_7369# tdc1.r_dly_store_ctr[15] a_9871_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6357 VPWR a_13599_6196# tdc1.w_ring_buf[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6358 tdc0.r_dly_store_ring[14] a_10443_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6359 a_29733_7663# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
R81 net58 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6360 VPWR a_4219_13621# _161_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X6361 a_10957_6031# a_10791_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6362 VGND tdc1.w_ring_norsz[20] a_22935_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6363 a_27425_6581# a_27259_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6364 a_4613_9839# tdc0.w_ring_buf[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6365 _092_ a_26891_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6366 VGND net26 a_6835_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6367 a_23273_10383# a_22719_10357# a_22926_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6368 VGND tdc1.w_ring_norsz[25] a_28271_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6370 a_14223_14191# a_13441_14197# a_14139_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6371 a_5015_9622# tdc1.r_dly_store_ring[0] a_4943_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X6372 tdc0.r_ring_ctr[4] a_12599_16671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6374 a_23087_15583# a_22912_15657# a_23266_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6375 tdc0.w_ring_int_norsz[9] tdc0.w_ring_norsz[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6376 VPWR a_22565_15253# a_22455_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6377 a_11623_12335# _124_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
X6378 a_19375_6575# a_18593_6581# a_19291_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6379 VPWR tdc1.w_ring_int_norsz[26] a_27793_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6381 VGND tdc1.w_ring_norsz[0] tdc1.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6383 a_13054_14735# _037_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6384 VPWR tdc0.r_ring_ctr[12] _159_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6385 VPWR tdc1.w_ring_norsz[12] a_25777_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6386 VPWR a_30254_7895# a_30203_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6387 VGND a_21891_15797# a_21825_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X6388 _177_ a_13919_4512# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X6389 VGND net45 tdc0.w_ring_int_norsz[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6390 VPWR _143_ a_9647_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X6391 a_29181_9545# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X6392 VGND tdc0.w_ring_norsz[4] tdc0.w_ring_norsz[20] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6394 a_2765_11293# a_2287_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X6395 VPWR a_5767_11837# a_5935_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6396 a_11709_3009# a_11491_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6397 a_13635_8867# _188_ a_13553_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6398 a_26781_6575# tdc1.w_ring_norsz[28] a_26697_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6399 tdc0.w_ring_int_norsz[2] tdc0.w_ring_norsz[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6400 a_18776_9071# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X6403 a_22695_5487# a_21831_5493# a_22438_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6404 VPWR a_17935_4703# a_17922_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6405 VPWR tdc1.w_ring_int_norsz[13] a_18869_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6406 a_16595_14985# _154_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6407 a_13728_11471# _077_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6408 _004_ a_6364_14985# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6409 VPWR _075_ a_20341_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6410 VGND a_19310_5055# a_19268_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6411 a_14983_14165# tdc0.w_ring_buf[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6412 a_21637_9545# tdc0.r_dly_store_ring[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X6413 a_16385_10927# tdc0.w_ring_norsz[21] a_16301_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6414 VGND a_8451_15797# tdc0.r_ring_ctr[6] VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X6415 a_16732_15823# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6416 a_10359_12015# a_9577_12021# a_10275_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6418 VPWR a_17739_7882# tdc1.w_ring_buf[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6420 VGND a_15504_9295# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6421 a_11709_3009# a_11491_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6422 a_13450_5764# a_13250_5609# a_13599_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6423 VGND _064_ _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6424 tdc1.w_ring_buf[0] a_5547_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6425 tdc1.r_dly_store_ring[3] a_25347_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6426 a_13629_6575# tdc1.w_ring_buf[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6427 tdc0.r_dly_store_ring[4] a_22311_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6428 VGND _115_ a_15256_10535# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6429 VPWR tdc0.w_ring_int_norsz[3] a_22917_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6430 VPWR net35 a_23395_14197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6431 a_20333_8029# _064_ a_20261_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
R82 tdc1.g_ring3[16].stg01_61.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6432 a_10977_9955# _136_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6434 a_29871_8573# a_29173_8207# a_29614_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6435 a_24696_9129# a_24297_8757# a_24570_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6436 VGND net1 a_26983_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6437 _088_ a_20175_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6439 VGND a_16587_8207# _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6440 a_4529_4943# a_3339_4943# a_4420_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
R83 VGND net70 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6442 a_17167_9839# a_16385_9845# a_17083_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6444 _001_ _154_ a_16845_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X6445 VPWR tdc0.w_ring_norsz[4] a_20727_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6446 VPWR a_24259_14191# a_24427_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6447 a_18496_14569# a_17581_14197# a_18149_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6448 VGND a_25474_3967# a_25432_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6449 VGND a_10124_9269# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X6450 a_27817_8457# tdc1.w_ring_norsz[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6451 a_10239_14735# _145_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6452 VGND _083_ a_15772_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
R84 tt_um_hpretl_tt06_tdc_v2_81.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6454 a_24646_6549# a_24478_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6455 VGND a_9282_13077# a_9240_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6457 a_6430_6549# a_6262_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6458 a_14008_9545# _194_ a_13620_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6459 VPWR _151_ a_10699_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6461 VGND _106_ a_28731_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6462 VGND net18 tdc1.w_ring_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R85 net68 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6463 a_10291_4373# _168_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X6464 VPWR _161_ a_4249_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6465 tdc1.r_dly_store_ring[24] a_12651_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6467 tdc1.w_ring_norsz[10] net17 a_27437_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6468 a_17302_5487# a_17029_5493# a_17217_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6469 a_10045_14735# _145_ a_9939_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X6470 a_24462_14847# a_24294_15101# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6471 a_23377_6575# tdc1.w_ring_norsz[4] a_23293_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6472 a_4698_9839# a_4425_9845# a_4613_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6473 a_13717_7369# tdc1.r_dly_store_ctr[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6474 tdc1.w_ring_norsz[16] net15 a_6077_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6475 VGND tdc0.r_ring_ctr[0] a_19723_15279# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6476 tdc0.w_ring_buf[30] a_8583_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6478 a_13533_3317# a_13367_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6479 VPWR a_21327_7895# tdc1.r_dly_store_ring[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6480 a_9539_13103# a_8841_13109# a_9282_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6481 tdc0.r_dly_store_ctr[14] a_6027_13915# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6482 a_9114_13103# a_8675_13109# a_9029_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6483 VGND _057_ a_17273_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6484 VPWR tdc1.r_dly_store_ring[13] a_15543_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6485 _142_ a_20083_14735# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X6486 a_19881_12015# tdc0.w_ring_norsz[28] a_19797_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6487 a_3854_9407# a_3686_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6488 a_24251_5487# a_23469_5493# a_24167_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6489 VGND a_23080_14165# net35 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6490 a_27951_12247# a_28047_12247# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6491 a_7385_15253# a_7167_15657# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6492 a_13450_5764# a_13243_5705# a_13626_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6493 VPWR tdc0.r_ring_ctr[8] a_15627_14709# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
R86 VPWR tdc1.g_ring3[20].stg01_65.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6494 VPWR net28 a_6191_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6495 VPWR a_13620_9269# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6496 a_25474_14165# a_25306_14191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6499 tdc1.w_ring_int_norsz[30] net75 a_14293_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6500 VGND _192_ a_14197_10389# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6501 a_14724_15823# a_13809_15823# a_14377_16065# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6502 VPWR net35 a_23855_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6503 a_17740_10071# tdc1.r_dly_store_ring[5] a_17882_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6504 a_16127_14557# tdc0.r_ring_ctr[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X6505 VPWR _075_ a_26513_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6507 VGND net31 a_17139_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6508 a_20506_3677# _048_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6509 VGND tdc0.w_ring_norsz[3] tdc0.w_ring_int_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6511 net32 a_17100_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6512 VGND tdc0.w_ring_norsz[18] a_26063_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6513 tdc1.w_ring_buf[28] a_27075_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6514 VGND _097_ a_25973_9301# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6515 a_10449_15617# _143_ a_10363_15617# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6518 a_9551_15511# _145_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X6519 _173_ a_9811_4737# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X6520 a_5989_6581# a_5823_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6521 a_24259_14191# a_23395_14197# a_24002_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6522 a_19066_7895# a_19425_7895# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X6525 a_6743_7663# tdc1.w_ring_norsz[16] a_6997_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6526 a_6895_14569# a_6449_14197# a_6799_14569# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6527 _063_ net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6528 a_7577_11721# tdc0.w_ring_norsz[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6529 a_7072_15645# _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6531 a_17229_4097# a_17011_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6532 VGND a_13887_8359# _186_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X6534 a_26529_8457# tdc1.w_ring_norsz[26] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6535 VGND a_14011_9839# _075_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6538 a_14064_15823# _014_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6539 a_20533_6575# _084_ a_20451_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6540 a_13797_5865# a_13243_5705# a_13450_5764# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6541 VGND a_9631_6397# a_9799_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6542 tdc1.w_ring_norsz[21] tdc1.w_ring_norsz[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6544 VGND net34 a_24131_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6545 a_8865_10927# tdc0.w_ring_norsz[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6546 a_9025_8207# a_8859_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6547 VPWR a_6027_13915# a_5943_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6548 VGND a_19735_13915# a_19693_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6550 a_15906_6143# a_15738_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6551 a_11867_6691# _127_ a_11795_6691# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6552 a_3763_7119# a_3247_7119# a_3668_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6554 VGND a_17435_13077# a_17393_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6555 a_15906_6143# a_15738_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6556 VGND tdc1.w_ring_norsz[18] tdc1.w_ring_norsz[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6557 a_16669_10927# net23 tdc0.w_ring_norsz[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6558 VPWR a_8008_4777# a_8183_4703# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6559 VGND a_11115_4007# _171_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6560 a_18690_8751# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6561 VGND a_23179_3829# a_23113_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X6562 net36 a_23671_15287# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X6563 VPWR a_10291_4373# _181_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X6564 VGND net9 a_11343_16373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6565 VPWR net7 a_8123_3317# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6568 a_3526_10927# a_2807_11169# a_2963_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X6569 VPWR tdc0.r_ring_ctr[8] a_12905_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6570 _147_ tdc0.r_ring_ctr[4] a_11426_15599# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X6571 a_16845_9295# a_16679_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6572 _010_ _143_ a_11049_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X6573 a_6888_3855# _029_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X6574 VPWR net35 a_23119_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6575 a_6541_4943# tdc1.r_ring_ctr[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6576 a_19057_10383# tdc0.w_ring_buf[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6578 VGND tdc1.w_ring_norsz[16] a_7111_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6579 VPWR tdc0.w_ring_norsz[31] a_5629_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6580 a_12586_16367# a_11509_16373# a_12424_16745# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6581 VPWR net34 a_24039_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6582 _189_ a_13553_8867# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X6584 VPWR a_15023_5487# net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6585 a_13626_5487# a_13379_5865# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6586 tdc0.r_ring_ctr[12] a_5055_14709# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X6587 tdc1.r_ring_ctr[8] a_14623_3615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X6588 a_28249_6953# a_27259_6581# a_28123_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6589 VGND a_19291_10927# a_19459_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6591 a_8749_4943# a_8583_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6592 VPWR a_4463_10651# a_4379_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6593 a_3951_4943# a_3505_4943# a_3855_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
R87 uio_oe[6] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6594 VPWR a_26847_9460# tdc1.w_ring_buf[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6595 a_24021_4399# a_23487_4405# a_23926_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6596 VPWR a_25731_13103# a_25899_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6597 a_4698_8751# a_4425_8757# a_4613_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6598 VGND net27 a_6191_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6600 VPWR _195_ _038_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6601 a_21886_9813# a_21718_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6602 VPWR a_4595_4917# a_4582_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6603 a_22609_15645# a_22565_15253# a_22443_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6604 tdc0.r_ring_ctr[5] a_12875_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6605 a_3413_9295# a_3247_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6606 VGND tdc1.r_ring_ctr[1] a_20531_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X6607 a_25409_12015# _077_ a_25493_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6610 a_23080_14165# net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X6611 VPWR ui_in[2] a_855_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6612 VGND a_6246_10495# a_6204_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6613 VGND net35 a_26431_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6614 a_6449_14197# a_6283_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6616 a_9623_13103# a_8841_13109# a_9539_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6617 VPWR _171_ a_10505_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6619 _138_ a_10977_9955# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X6622 VPWR tdc0.r_ring_ctr[4] a_11219_14887# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6623 a_22346_13077# a_22178_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6624 VPWR a_30039_8475# a_29955_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6625 VPWR a_15135_11989# a_15051_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6627 VPWR a_22863_5461# a_22779_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6628 tdc1.w_ring_norsz[24] net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6629 a_20763_11837# a_19899_11471# a_20506_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6631 a_19065_12015# tdc0.w_ring_norsz[26] a_18981_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6632 a_3413_12559# a_3247_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6633 a_5507_6005# _181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X6634 a_28441_7663# tdc1.w_ring_buf[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6635 a_11781_6031# a_10791_6031# a_11655_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6636 a_5893_11471# a_4903_11471# a_5767_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6638 a_15105_13423# tdc0.r_dly_store_ctr[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6639 VGND a_13203_4373# a_13161_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6640 VPWR tdc1.r_ring_ctr[3] a_21279_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6641 VPWR tdc1.w_ring_int_norsz[29] a_19237_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6642 a_6521_13621# tdc0.r_ring_ctr[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X6643 a_13629_14191# tdc0.r_ring_ctr[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6644 a_20433_11837# a_19899_11471# a_20338_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6645 VGND _038_ a_8689_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X6646 VPWR a_30856_7895# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6648 VPWR tdc1.w_ring_int_norsz[15] a_7645_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6649 VGND a_12594_7637# a_12552_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6650 tdc0.r_dly_store_ctr[4] a_12375_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6651 a_19057_4943# tdc1.r_ring_ctr[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6653 tdc0.r_dly_store_ring[23] a_8695_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6656 tdc1.w_dly_stop[4] a_27167_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6657 VGND _064_ a_19439_9111# VGND sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X6658 tdc1.r_dly_store_ring[13] a_14307_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6659 a_11601_12809# tdc0.r_dly_store_ring[22] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6661 a_26973_12809# _091_ a_26891_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6662 a_21905_13109# a_21739_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6663 a_17393_13481# a_16403_13109# a_17267_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6664 a_27790_5487# a_27351_5493# a_27705_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6665 VPWR tdc1.r_dly_store_ring[26] a_29181_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X6666 a_15269_14735# tdc0.r_ring_ctr[9] a_15197_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6670 tdc0.r_ring_ctr[10] a_18671_14495# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6671 a_29871_8573# a_29007_8207# a_29614_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6672 VPWR a_7732_15657# a_7907_15583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6673 VGND a_23910_5461# a_23868_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6674 VGND _195_ _041_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6675 VGND a_14583_13915# a_14541_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6676 a_12659_10749# a_11877_10383# a_12575_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6677 a_21259_16189# a_20635_15823# a_21151_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6678 tdc1.w_ring_norsz[6] tdc1.w_ring_norsz[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6680 a_16842_13103# a_16569_13109# a_16757_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6681 VGND net31 a_18703_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6682 VPWR a_17470_5461# a_17397_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6684 VGND a_17895_5461# a_17853_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6685 VPWR a_4866_9813# a_4793_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6686 VGND a_13450_5764# a_13379_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6687 a_30254_7895# a_30350_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X6689 a_9121_6031# tdc1.w_ring_buf[30] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6690 a_27563_9839# a_26781_9845# a_27479_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6691 a_6725_12925# a_6191_12559# a_6630_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6692 VGND _195_ _040_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6693 uo_out[0] a_13620_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6694 tdc0.r_dly_store_ring[3] a_25071_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6695 tdc1.w_ring_buf[16] a_6743_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6698 a_9690_16189# a_8932_16091# a_9127_16060# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X6699 VGND tdc1.r_ring_ctr[5] _170_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6700 VPWR _083_ a_20617_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6701 VGND tdc1.w_ring_norsz[30] tdc1.w_ring_int_norsz[31] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6703 a_14300_11305# a_13901_10933# a_14174_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6704 VGND net32 a_16219_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6705 a_9374_6143# a_9206_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6706 a_18850_14557# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6707 VGND tdc0.w_ring_int_norsz[30] tdc0.w_ring_norsz[30] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6708 a_21886_8725# a_21718_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6710 a_9374_6143# a_9206_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6711 a_7902_8725# a_7734_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6713 VGND _196_ _053_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6714 a_21980_9545# _111_ a_21637_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X6716 VGND tdc1.r_ring_ctr[13] a_5997_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6717 tdc1.w_ring_buf[19] a_23855_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6718 a_20506_11583# a_20338_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6719 VPWR net14 a_18151_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6720 VPWR a_20506_11583# a_20433_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6721 VGND _102_ a_25182_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6722 a_14557_3689# a_13367_3317# a_14448_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6723 a_22687_13103# a_21905_13109# a_22603_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6724 a_22811_3615# _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6725 net41 a_26983_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6726 VGND tdc0.r_ring_ctr[1] a_21157_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6727 a_9850_10927# a_9411_10933# a_9765_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6728 a_6798_9813# a_6630_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6730 a_17931_14569# a_17581_14197# a_17836_14557# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6731 a_8971_15965# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6733 a_7167_15657# a_6651_15285# a_7072_15645# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6734 a_26431_13103# _072_ a_26513_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6735 a_25472_8181# _101_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X6736 VGND tdc1.r_dly_store_ring[9] a_30389_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6737 a_7902_8725# a_7734_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6738 _093_ a_25327_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6739 VPWR net9 a_3247_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6741 a_15757_13889# a_15539_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6743 VPWR _064_ a_20157_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X6744 a_27916_5865# a_27517_5493# a_27790_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6745 tdc0.w_ring_norsz[24] net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6746 VGND net20 tdc0.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6747 a_12218_3133# a_11141_2767# a_12056_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6749 a_4793_9839# a_4259_9845# a_4698_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6750 a_11398_6143# a_11230_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6751 VGND tdc1.w_ring_norsz[12] tdc1.w_ring_int_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6752 VGND tdc1.w_ring_norsz[3] tdc1.w_ring_int_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6753 VPWR tdc0.w_ring_norsz[1] a_19347_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6754 tdc1.w_ring_norsz[15] tdc1.w_ring_norsz[31] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6755 a_15335_8181# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6756 a_14155_4917# tdc1.r_ring_ctr[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X6757 a_10221_4943# a_10055_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6758 a_25137_7119# tdc1.r_dly_store_ctr[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6759 VPWR a_6798_12671# a_6725_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R88 VPWR tdc1.g_ring3[29].stg01_74.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6761 a_22351_9545# _084_ a_22257_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X6763 a_13797_5865# a_13250_5609# a_13450_5764# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6764 _081_ a_18243_8751# a_18776_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6765 VPWR tdc0.r_ring_ctr[12] a_6739_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X6766 a_3686_8573# a_3247_8207# a_3601_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6768 a_12291_6183# tdc1.r_dly_store_ctr[6] a_12437_6281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6769 a_12529_13423# tdc0.r_dly_store_ctr[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6771 VPWR a_4866_8725# a_4793_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6773 a_19651_5309# a_18869_4943# a_19567_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6777 VGND a_29587_7895# _101_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6778 _139_ a_6027_9622# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X6779 a_13979_3689# a_13533_3317# a_13883_3689# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6780 VGND a_5123_9839# a_5291_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6782 VPWR net32 a_18703_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6783 a_18751_8359# tdc1.r_dly_store_ring[6] a_18991_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X6784 VGND _086_ a_25511_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6785 a_2287_10901# a_2490_11059# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X6786 VGND _072_ a_15564_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6787 VGND net34 a_28455_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6788 net20 a_3399_12275# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X6789 tdc0.r_dly_store_ring[1] a_20655_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6791 a_4774_4943# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6792 a_3505_6031# a_3339_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6793 a_16209_8751# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6794 tdc0.w_ring_norsz[20] tdc0.w_ring_int_norsz[20] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6795 a_6430_6549# a_6262_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6796 VPWR a_9723_8573# a_9891_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6797 a_17567_15797# a_17392_15823# a_17746_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6798 VPWR net29 a_9871_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6799 VPWR a_4073_5185# a_3963_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6800 VPWR net5 a_16309_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X6801 _060_ net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6804 a_23293_12015# net40 tdc0.w_ring_int_norsz[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6805 VPWR _152_ a_13073_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6806 tdc1.r_ring_ctr[4] a_17935_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X6807 VPWR tdc1.r_ring_ctr[10] a_14155_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X6809 a_9025_8207# a_8859_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6812 a_6545_9839# tdc0.w_ring_buf[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6813 a_10409_4943# tdc1.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6814 a_3981_7361# a_3763_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6815 VGND tdc0.w_ring_norsz[22] tdc0.w_ring_int_norsz[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6816 a_15261_11445# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X6817 tdc0.w_ring_int_norsz[31] net58 a_7577_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6819 VGND a_14415_14013# a_14583_13915# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6820 a_17746_8319# a_17578_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6821 a_15809_12234# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6822 tdc1.w_ring_norsz[17] tdc1.w_ring_int_norsz[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6824 a_15925_15823# _153_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6825 VPWR a_14377_16065# a_14267_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6826 VPWR a_8159_8751# a_8327_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6828 a_17746_8319# a_17578_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6829 VPWR a_27411_7093# net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X6831 a_13887_8359# tdc1.r_dly_store_ctr[0] a_14061_8235# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6832 VPWR tdc0.w_ring_norsz[21] a_13459_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6833 VGND a_25731_14191# a_25899_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6834 a_23273_10383# a_22726_10657# a_22926_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6835 tdc0.w_ring_int_norsz[8] net38 a_8865_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6837 a_10512_9545# _083_ a_10124_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X6838 uo_out[2] a_26420_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6840 a_9558_3677# _054_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6841 _016_ tdc1.r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6842 a_18496_14569# a_17415_14197# a_18149_14165# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6843 tdc1.r_dly_store_ctr[3] a_24519_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6844 a_6983_3855# a_6467_3855# a_6888_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6845 _068_ a_16309_8867# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X6846 VGND _070_ a_14332_8983# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X6848 VGND a_3799_13103# net24 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6849 a_22917_11721# tdc0.w_ring_norsz[19] a_22833_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6850 a_26513_13103# tdc0.r_dly_store_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6851 a_17760_4777# a_16845_4405# a_17413_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6852 VGND a_26615_7119# net18 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6853 VGND _137_ a_10977_9955# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6855 a_12341_7663# tdc1.w_ring_buf[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6856 a_19798_14735# tdc0.r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X6858 a_26985_8751# tdc1.w_ring_int_norsz[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6859 VPWR _196_ _055_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6860 a_25214_5487# a_24775_5493# a_25129_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6861 VGND _196_ _054_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6862 a_21912_6575# _108_ a_21826_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6863 a_20341_9295# _070_ a_20241_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X6865 a_7810_13077# a_7642_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6867 VGND _068_ a_11045_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6868 a_26420_11721# _098_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X6869 tdc1.w_dly_stop[4] a_27167_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6870 VGND _084_ a_13551_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6871 a_14973_9839# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X6872 a_4793_8751# a_4259_8757# a_4698_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6873 a_5434_14013# a_5161_13647# a_5349_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6874 VPWR _181_ a_5907_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6875 a_5694_7231# a_5526_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6878 VGND a_18703_14735# _195_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6879 a_22143_9839# a_21279_9845# a_21886_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6880 a_22455_15279# a_21831_15285# a_22347_15657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6881 a_22097_12015# net54 tdc0.w_ring_int_norsz[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6882 a_5694_7231# a_5526_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6883 a_3812_8207# a_3413_8207# a_3686_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6886 a_28215_5487# a_27517_5493# a_27958_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
R89 VPWR tdc0.g_ring3[24].stg01_51.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R90 VGND net57 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6887 VPWR a_20327_3615# tdc1.r_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R91 VGND net55 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6890 a_23657_5487# tdc1.r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6891 VGND a_27351_8207# net40 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6892 a_12345_8457# net70 tdc1.w_ring_int_norsz[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6893 tdc0.r_dly_store_ring[23] a_8695_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6894 a_12823_16073# _152_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6895 a_27698_6575# a_27425_6581# a_27613_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6896 tdc1.r_dly_store_ctr[10] a_19735_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6897 a_5042_15101# a_3965_14735# a_4880_14735# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6898 tdc1.w_ring_buf[11] a_27903_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6899 a_30101_8751# _072_ a_29955_8983# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X6900 a_11329_13103# tdc0.w_ring_buf[22] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6901 VPWR a_5859_14013# a_6027_13915# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6902 a_9939_14735# _150_ a_9843_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X6903 VPWR net28 a_8767_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6904 a_19797_12015# net22 tdc0.w_ring_norsz[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R92 uio_out[6] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6905 tdc1.r_ring_ctr[15] a_4503_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6906 VGND tdc0.w_ring_buf[20] a_23273_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6907 a_18785_7369# net41 tdc1.w_ring_int_norsz[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6908 a_29446_8573# a_29007_8207# a_29361_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6909 a_20046_4765# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6910 a_20883_9955# _110_ a_20811_9955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6911 VPWR a_13735_12559# net23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6913 uo_out[5] a_15504_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6914 a_26973_12809# _067_ a_27057_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6915 VPWR _175_ a_13919_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6917 _062_ net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6919 a_3870_10749# a_3597_10383# a_3785_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6920 net14 a_12539_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6921 a_4315_14735# a_3799_14735# a_4220_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6922 a_5043_8372# tdc1.w_ring_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6923 a_3505_11721# tdc0.r_ring_ctr[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6924 a_30856_7895# ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X6926 VGND _086_ a_4761_9622# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X6927 a_15093_12393# a_14103_12021# a_14967_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6931 a_22001_13647# tdc0.r_ring_ctr[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6932 _081_ a_18243_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6933 VPWR _196_ _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6934 a_14710_11989# a_14542_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6935 VGND net23 _043_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6936 VPWR a_18496_14569# a_18671_14495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6938 VGND _052_ a_17457_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6939 a_4328_7119# a_3413_7119# a_3981_7361# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6942 a_22143_8751# a_21445_8757# a_21886_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6943 a_9850_12015# a_9577_12021# a_9765_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
R93 tdc1.stg01_77.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6944 VPWR tdc1.w_ring_int_norsz[16] a_6559_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6945 a_3392_8725# net26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6946 a_21511_9447# _086_ a_21980_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6947 a_8803_12015# a_7939_12021# a_8546_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6949 VGND net33 a_17323_8759# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6950 _082_ a_19655_8235# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X6952 a_14542_12015# a_14269_12021# a_14457_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6953 VPWR a_16163_6397# a_16331_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6954 VGND _071_ a_12539_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6956 a_12165_2767# a_10975_2767# a_12056_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6957 VPWR a_20083_8751# _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6958 a_19854_4399# a_18777_4405# a_19692_4777# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6959 a_24903_6575# a_24205_6581# a_24646_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6960 a_8102_7663# a_7829_7669# a_8017_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6961 a_25121_13647# tdc0.r_dly_store_ctr[3] a_24683_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6962 a_6687_6575# a_5989_6581# a_6430_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6963 a_21843_8041# a_21714_7785# a_21423_7895# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6964 VGND _118_ a_15025_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6965 a_8473_12015# a_7939_12021# a_8378_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6966 a_24259_14191# a_23561_14197# a_24002_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6967 _024_ _163_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6968 a_17669_9295# a_16679_9295# a_17543_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6969 a_27149_9839# a_26615_9845# a_27054_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6970 a_6545_12559# tdc0.r_ring_ctr[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6971 tdc1.r_dly_store_ctr[11] a_17895_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6972 VPWR _195_ _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6973 a_23082_14735# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6974 a_20966_5055# a_20798_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6975 a_21891_15797# a_21716_15823# a_22070_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6976 a_25340_5865# a_24941_5493# a_25214_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6978 VGND _068_ a_10975_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6979 a_28215_5487# a_27351_5493# a_27958_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6980 a_22261_8041# a_21714_7785# a_21914_7940# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6981 a_26575_11159# a_26866_11049# a_26817_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6982 a_11792_12015# _130_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X6984 VPWR a_22811_3615# a_22798_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6985 VGND tdc0.w_ring_int_norsz[23] tdc0.w_ring_norsz[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6986 _075_ a_14011_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6987 tdc0.w_ring_int_norsz[13] net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6988 VPWR a_15809_12234# tdc0.w_ring_buf[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6989 VPWR a_15703_7485# a_15871_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6991 VGND a_13599_6196# tdc1.w_ring_buf[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6992 a_11049_15823# tdc0.r_ring_ctr[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6993 VGND net9 a_6651_15285# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6994 VGND a_3854_8319# a_3812_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6995 a_3399_12275# net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X6996 a_27709_8751# net18 tdc1.w_ring_norsz[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R94 net66 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6998 a_22143_8751# a_21279_8757# a_21886_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7002 tdc1.r_dly_store_ctr[10] a_19735_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7003 a_13379_5865# a_13250_5609# a_12959_5719# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7005 VGND tdc0.w_ring_int_norsz[4] tdc0.w_ring_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7007 _003_ _158_ a_3689_14511# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X7008 a_28894_8751# a_28621_8757# a_28809_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7009 a_25474_13077# a_25306_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7010 VGND _141_ _008_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7011 VGND net20 _044_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7014 a_24941_5493# a_24775_5493# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7017 _038_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7018 VPWR net26 a_4259_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7019 VPWR a_18703_14735# _195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7020 a_29572_8207# a_29173_8207# a_29446_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R95 tdc1.g_ring1[16].stg02_60.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7021 a_4111_8573# a_3413_8207# a_3854_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7022 a_25847_8751# _073_ a_25755_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X7023 a_18776_9071# _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7026 VGND tdc0.w_ring_int_norsz[16] tdc0.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7027 a_18785_6281# net19 tdc1.w_ring_norsz[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7028 a_11587_2767# a_11141_2767# a_11491_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7029 tdc1.w_ring_int_norsz[6] net41 a_17881_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7030 a_18169_10137# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X7031 a_20986_14013# a_20739_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7032 VPWR a_25071_9813# a_24849_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X7033 VPWR a_25639_5487# a_25807_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7035 VPWR _066_ a_15289_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7036 VGND tdc1.w_ring_norsz[22] tdc1.w_ring_int_norsz[23] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7037 a_9209_13103# a_8675_13109# a_9114_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7038 a_10321_14735# _143_ a_10239_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7039 a_25401_14191# a_24867_14197# a_25306_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7041 VGND a_7897_7284# net13 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7042 tdc0.w_ring_norsz[13] tdc0.w_ring_norsz[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7043 VGND net9 a_3247_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7044 _123_ a_10147_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7046 VGND _064_ _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7047 a_8611_9839# a_7829_9845# a_8527_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7049 VPWR a_8546_11989# a_8473_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7051 VGND tdc1.w_ring_int_norsz[18] tdc1.w_ring_norsz[18] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7052 a_29955_7485# a_29173_7119# a_29871_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7053 a_11233_11721# tdc0.r_dly_store_ring[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7054 a_18869_4943# a_18703_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7056 VGND a_12291_6183# _126_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X7057 a_13901_10933# a_13735_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7058 VPWR tdc1.r_dly_store_ctr[10] a_20157_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X7059 a_24591_9545# tdc1.r_dly_store_ring[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X7060 _191_ a_10699_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7061 VGND a_12207_14191# a_12375_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7062 a_21457_7119# tdc1.r_dly_store_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X7064 VPWR net35 a_24039_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7065 a_24209_12015# tdc0.w_ring_buf[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
R96 net65 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7066 VPWR a_26983_8207# net41 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7067 tdc0.w_ring_buf[19] a_23303_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7068 a_23561_14197# a_23395_14197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7069 VGND a_10662_5055# a_10620_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7070 a_19237_5309# a_18703_4943# a_19142_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7071 a_17209_10217# a_16219_9845# a_17083_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7072 VGND tdc0.w_ring_norsz[4] a_20727_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7074 VPWR _038_ a_9272_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X7076 a_22837_14735# a_21647_14735# a_22728_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7077 a_17685_3855# a_16495_3855# a_17576_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7078 a_6997_7663# tdc1.w_ring_norsz[16] a_6743_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7079 a_16923_15823# a_16477_15823# a_16827_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7080 VGND _051_ a_22701_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7081 a_25179_7663# a_24315_7669# a_24922_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7082 tdc0.r_dly_store_ring[9] a_18171_12827# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7083 a_23179_3829# a_23004_3855# a_23358_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7084 VPWR a_19310_10495# a_19237_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7085 a_9765_10927# tdc0.w_ring_buf[24] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7086 VPWR a_12875_14709# a_12862_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7088 a_6248_9295# tdc1.r_dly_store_ring[7] a_6027_9622# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7089 VPWR a_22311_9813# a_22227_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7090 a_11509_16373# a_11343_16373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7091 tdc1.r_ring_ctr[12] a_8183_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7092 a_7907_15583# _039_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7093 tdc1.w_ring_int_norsz[3] net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7094 a_16458_13647# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7095 tdc0.r_dly_store_ring[25] a_19735_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7096 VGND _128_ a_18751_8359# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X7097 a_6798_12671# a_6630_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7098 a_14800_6549# tdc1.w_dly_stop[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X7099 tdc1.r_dly_store_ctr[13] a_6855_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7100 VGND a_23818_13077# a_23776_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7101 tdc0.r_dly_store_ctr[5] a_14307_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7103 VPWR a_27866_6549# a_27793_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7104 VPWR tdc1.w_ring_int_norsz[23] a_11325_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7105 a_20613_12559# a_19623_12559# a_20487_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7106 a_9263_7485# a_8565_7119# a_9006_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7107 a_24029_12809# tdc0.r_dly_store_ring[11] a_23947_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7108 VGND net29 a_9871_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7110 VPWR net25 a_9577_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7111 a_21377_15279# _143_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7112 _034_ _195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7113 tdc0.w_ring_buf[21] a_13459_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7115 VGND a_29614_8319# a_29572_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7116 a_5207_9839# a_4425_9845# a_5123_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7118 a_9647_14709# _145_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X7119 a_22657_4097# a_22439_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7120 tdc1.w_ring_norsz[3] tdc1.w_ring_norsz[19] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7121 tdc1.w_ring_buf[31] a_7295_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7126 a_17410_13647# a_17095_13799# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7127 a_4421_10383# a_3431_10383# a_4295_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7129 VPWR a_25474_14165# a_25401_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7130 a_21633_9839# tdc0.w_ring_buf[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7131 a_5043_11146# tdc0.w_ring_norsz[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7134 VPWR net28 a_7663_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7135 a_20739_13647# a_20603_13621# a_20319_13621# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7137 _071_ a_15159_8725# a_14909_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7138 VGND _195_ _036_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7139 tdc0.w_ring_norsz[11] tdc0.w_ring_int_norsz[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7140 _137_ a_9411_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X7141 VPWR tdc0.w_ring_norsz[2] a_23293_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7143 a_25182_10383# _102_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7144 VGND a_13511_7895# _188_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X7146 a_19977_12559# tdc0.w_ring_buf[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7147 tdc1.w_ring_buf[28] a_27075_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7148 VPWR a_19535_7637# a_19066_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X7149 a_18961_10927# a_18427_10933# a_18866_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7150 a_6027_9622# tdc1.r_dly_store_ring[7] a_5955_9622# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X7151 a_9577_12021# a_9411_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7153 a_13073_15823# tdc0.r_ring_ctr[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7154 a_11877_10383# a_11711_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7155 VGND _149_ _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7156 a_27445_7663# tdc1.w_ring_int_norsz[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7157 VPWR a_8270_7637# a_8197_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7158 VGND a_8971_15965# a_8932_16091# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7159 VGND net15 tdc1.w_ring_norsz[16] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7160 a_14269_12021# a_14103_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7162 VGND a_16771_7663# _070_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7165 VGND net30 a_13275_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7166 a_11540_13481# a_11141_13109# a_11414_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7168 a_11035_3543# _166_ a_11209_3649# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7169 a_10310_14013# a_9871_13647# a_10225_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7170 tdc0.r_ring_ctr[2] a_22903_14709# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X7171 VPWR a_28383_5461# a_28299_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7173 VGND tdc0.w_ring_norsz[8] tdc0.w_ring_norsz[24] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7174 a_6291_5193# _181_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7175 VPWR a_17760_2767# a_17935_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7176 _193_ a_14197_10389# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X7177 a_23947_12809# _072_ a_24029_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7178 a_21413_15823# a_21369_16065# a_21247_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X7179 a_27793_6575# a_27259_6581# a_27698_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7180 _143_ a_20503_15253# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7181 a_22447_9295# tdc1.r_dly_store_ring[2] a_22257_9545# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7184 net27 a_2932_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7185 tdc1.r_dly_store_ctr[1] a_24335_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7186 tdc1.w_ring_buf[3] a_24223_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7188 a_18869_13647# a_18703_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7189 a_17493_8207# tdc1.w_ring_buf[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7190 a_14499_14013# a_13717_13647# a_14415_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7191 VPWR a_17751_3829# tdc1.r_ring_ctr[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7192 a_3854_9407# a_3686_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7193 VGND _069_ a_25949_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X7194 VPWR a_18171_12827# a_18087_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7195 VPWR _196_ _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7196 VPWR a_22311_8725# a_22227_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7198 VPWR net12 a_22097_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7199 a_10761_3855# _168_ a_10689_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7200 VPWR a_30537_7895# a_30350_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7201 a_3963_6397# _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7202 VGND a_26847_9460# tdc1.w_ring_buf[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7203 _010_ a_10799_16073# a_11049_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X7204 a_21707_7881# net33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7205 a_3601_8207# net7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7206 a_19219_15823# a_18703_15823# a_19124_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7207 VPWR net7 a_3339_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7208 a_9466_8319# a_9298_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7209 VGND ui_in[2] a_855_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7211 _030_ a_12731_3311# a_12981_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X7212 VPWR a_28951_9839# a_29119_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7213 VGND a_7223_12827# a_7181_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7214 VGND a_19959_15797# a_19893_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X7217 VPWR a_15481_5185# a_15371_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X7218 a_5207_8751# a_4425_8757# a_5123_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7220 a_5441_7119# tdc1.r_ring_ctr[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7221 VGND a_20487_12925# a_20655_12827# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7223 a_11764_16733# _010_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7224 VPWR tdc1.r_ring_ctr[8] a_13919_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7225 VGND a_27463_11989# a_27421_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7227 VGND _161_ _005_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7230 a_7723_3829# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7231 VGND a_17711_9563# a_17669_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7232 a_24987_10927# a_24205_10933# a_24903_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7233 VPWR tdc0.w_ring_int_norsz[19] a_23285_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7234 _017_ a_15399_4399# a_15649_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X7235 VPWR net15 _062_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7236 a_25949_11247# tdc0.r_dly_store_ring[27] a_25511_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7237 a_12981_3311# tdc1.r_ring_ctr[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7238 VGND a_4295_10749# a_4463_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7239 VPWR tdc0.w_ring_buf[26] a_28885_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7240 a_18777_8029# _065_ a_18677_8029# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X7241 a_10147_9839# _076_ a_10229_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7242 a_7829_7669# a_7663_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7243 tdc1.w_ring_int_norsz[26] tdc1.w_ring_norsz[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7244 a_18877_13103# tdc0.r_dly_store_ring[17] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7247 a_5997_4943# tdc1.r_ring_ctr[12] _182_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7248 a_20464_11471# a_20065_11471# a_20338_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7249 tdc1.w_ring_buf[16] a_6743_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7250 _026_ _166_ a_16385_3631# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X7252 a_14001_4765# tdc1.r_ring_ctr[8] a_13919_4512# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7253 VPWR a_25347_7637# a_25263_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7257 a_10173_10411# tdc0.r_dly_store_ring[31] a_10087_10411# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7258 a_9206_6397# a_8933_6031# a_9121_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7259 tdc1.w_ring_int_norsz[10] net40 a_27173_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7260 tdc1.w_ring_int_norsz[21] net66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7262 a_14139_6575# a_13275_6581# a_13882_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7263 VGND a_17470_5461# a_17428_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7264 a_10409_4943# tdc1.r_ring_ctr[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7265 VPWR a_5871_11146# tdc0.w_ring_buf[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7266 tdc1.r_dly_store_ring[25] a_30039_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7267 tdc0.r_ring_ctr[7] a_7907_15583# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7268 VPWR _196_ _056_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7269 tdc0.r_ring_ctr[11] a_16279_13621# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X7270 VPWR tdc0.w_dly_stop[1] a_2603_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7273 tdc0.r_ring_ctr[9] a_17567_15797# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X7274 VGND tdc0.w_ring_norsz[1] tdc0.w_ring_norsz[17] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7275 _066_ a_15335_8181# a_15283_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7277 VPWR tdc1.w_ring_norsz[2] a_21003_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7279 a_23661_6575# net40 tdc1.w_ring_int_norsz[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7280 a_7561_6575# net15 tdc1.w_ring_norsz[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7281 a_6473_12015# tdc0.w_ring_norsz[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7284 VPWR a_26859_11145# a_26866_11049# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7285 _153_ _152_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7286 VGND tdc1.r_ring_ctr[8] a_12731_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7288 a_20349_10927# net55 tdc0.w_ring_int_norsz[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7289 a_29733_7663# _072_ a_29587_7895# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X7290 a_27897_7663# tdc1.w_ring_norsz[11] a_27813_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7291 VPWR tdc0.w_ring_norsz[16] a_4627_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7292 VGND a_9615_5211# a_9573_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7293 VPWR a_23004_3855# a_23179_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7294 VGND net39 tdc1.w_ring_int_norsz[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7295 a_8197_9839# a_7663_9845# a_8102_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7296 a_12135_14735# a_11619_14735# a_12040_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7297 a_9263_7485# a_8399_7119# a_9006_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7298 VPWR a_25348_10633# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7299 VPWR _173_ a_10607_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7300 VGND tdc1.w_ring_norsz[11] tdc1.w_ring_int_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7301 VGND a_17375_7637# net39 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X7302 a_6077_8457# tdc1.w_ring_norsz[0] a_5823_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R97 net46 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7303 VGND _069_ a_29169_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X7304 tdc1.w_ring_int_norsz[27] tdc1.w_ring_norsz[26] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7307 a_27057_12809# tdc0.r_dly_store_ring[18] a_26973_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7308 a_21721_3317# a_21555_3317# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7309 VGND a_17251_9813# a_17209_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7310 a_9595_7663# _071_ a_9677_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7311 VPWR a_17567_15797# a_17554_16189# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7312 tdc1.w_ring_buf[19] a_23855_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
R98 VPWR tdc0.g_ring3[18].stg01_45.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7313 a_29361_8207# tdc1.w_ring_buf[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7314 a_19805_3285# a_19587_3689# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X7315 a_18129_8207# a_17139_8207# a_18003_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7316 VGND a_6521_13621# _160_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7318 a_12410_5055# a_12242_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7319 a_14267_16189# a_13643_15823# a_14159_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7320 _094_ a_20157_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7321 a_28885_12393# a_28331_12233# a_28538_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7322 VPWR a_16155_7895# _119_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7323 a_17291_4777# a_16845_4405# a_17195_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7324 VPWR net10 a_15023_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7325 VGND a_4595_6005# a_4529_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X7326 a_11141_13109# a_10975_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7327 a_10393_14735# _145_ a_10321_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7328 VGND tdc0.w_ring_int_norsz[0] tdc0.w_ring_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7330 VGND tdc1.w_ring_buf[0] a_15023_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X7331 a_3760_6031# _021_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7332 a_28652_10217# a_28253_9845# a_28526_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7333 VGND net14 a_18151_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7334 VPWR tdc0.w_ring_buf[27] a_27413_11305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7335 a_13788_3677# _030_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X7336 a_24021_8457# tdc1.w_ring_norsz[2] a_23937_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7337 a_27605_10217# a_26615_9845# a_27479_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7338 a_8504_12393# a_8105_12021# a_8378_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7339 a_18003_12925# a_17305_12559# a_17746_12671# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7340 tdc0.r_dly_store_ring[22] a_12007_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7342 tdc0.w_ring_int_norsz[11] net41 a_21009_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7344 VPWR net15 a_8399_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7346 a_18129_12559# a_17139_12559# a_18003_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7347 tdc0.r_dly_store_ring[22] a_12007_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7348 a_19793_5487# tdc1.r_ring_ctr[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7349 a_4117_6031# a_4073_6273# a_3951_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X7350 VGND a_17095_13799# tdc0.r_dly_store_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7351 VPWR a_13243_5705# a_13250_5609# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7352 a_15701_8457# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7353 VPWR a_4279_8475# a_4195_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7354 tdc0.r_dly_store_ctr[7] a_9247_14165# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7355 a_6077_7119# a_5087_7119# a_5951_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7356 a_11973_9295# tdc1.w_ring_buf[24] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7357 a_14089_10927# tdc0.w_ring_buf[21] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7358 a_19275_7983# tdc1.r_dly_store_ring[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
R99 VGND uio_out[5] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7359 a_13717_13109# a_13551_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7360 VPWR tdc1.r_ring_ctr[0] a_13797_5865# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X7362 tdc0.w_ring_norsz[26] net22 a_18697_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7364 a_7189_6031# tdc1.r_ring_ctr[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7365 tdc1.r_ring_ctr[2] a_19867_4703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7366 VGND tdc1.w_ring_norsz[21] tdc1.w_ring_int_norsz[22] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7367 VGND _065_ _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7368 a_16155_7895# tdc1.r_dly_store_ring[21] a_16301_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7369 a_3763_12559# a_3413_12559# a_3668_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7370 VGND tdc1.w_ring_int_norsz[7] tdc1.w_ring_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7371 VPWR a_3024_8725# _621_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7372 tdc0.w_ring_norsz[23] tdc0.w_ring_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7373 _149_ _146_ a_10337_16073# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7374 _141_ a_20727_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7375 a_14290_9111# _064_ a_14209_9111# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X7376 tdc0.r_dly_store_ring[29] a_14583_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7379 a_17922_3133# a_16845_2767# a_17760_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7380 VGND tdc1.w_ring_int_norsz[5] tdc1.w_ring_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7381 VGND net27 a_7203_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7382 a_19124_15823# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7384 _144_ tdc0.r_ring_ctr[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7385 tdc0.w_ring_int_norsz[24] net51 a_7853_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7386 VGND a_12318_10495# a_12276_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7387 a_9765_12015# tdc0.w_ring_buf[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7388 tdc0.r_dly_store_ring[29] a_14583_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7389 VGND tdc1.r_ring_ctr[9] a_15033_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X7391 a_20341_13103# tdc0.r_dly_store_ctr[9] a_20257_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7392 _072_ a_12539_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X7393 a_23841_4399# tdc1.r_ring_ctr[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7394 a_11230_6397# a_10957_6031# a_11145_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7395 tdc1.w_ring_norsz[19] tdc1.w_ring_norsz[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7396 VPWR a_17555_7284# tdc1.w_ring_buf[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7397 VGND tdc0.w_ring_norsz[20] tdc0.w_ring_int_norsz[21] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7398 a_14457_12015# tdc0.w_ring_buf[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7399 a_22344_3855# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7400 VGND a_22863_5461# a_22821_5865# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7401 _083_ a_20083_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7402 a_20249_6031# a_20083_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7403 a_27425_6581# a_27259_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7404 a_19417_6953# a_18427_6581# a_19291_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7405 a_8113_10927# net21 tdc0.w_ring_norsz[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7406 a_3689_14511# tdc0.r_ring_ctr[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7408 a_24478_6575# a_24039_6581# a_24393_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7410 a_6262_6575# a_5823_6581# a_6177_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7412 VPWR net25 a_13717_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7413 _046_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7414 _009_ _144_ a_21377_15279# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7415 _180_ _175_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7416 a_19057_10383# tdc0.w_ring_buf[25] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7417 _195_ a_18703_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7419 a_7055_9839# a_6357_9845# a_6798_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7420 VGND net31 a_20083_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7421 a_25609_8457# tdc1.r_dly_store_ring[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7423 VPWR tdc1.r_ring_ctr[2] a_20635_4512# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X7424 _620_.X a_3392_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7426 a_10217_7119# tdc1.r_dly_store_ctr[7] a_9871_7369# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7427 VGND a_13735_12559# net23 VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X7429 a_17930_3855# _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7430 a_21813_13647# a_21647_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7431 a_11003_5309# a_10221_4943# a_10919_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7432 a_17470_5461# a_17302_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7433 VPWR tdc0.w_ring_int_norsz[31] a_7461_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7436 a_18777_4405# a_18611_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7437 a_15569_14511# tdc0.r_ring_ctr[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7438 VPWR a_2840_12533# _622_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7439 VPWR a_16771_7663# _070_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7440 VGND net23 tdc0.w_ring_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7441 a_18039_14191# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7443 VGND tdc0.w_ring_int_norsz[1] tdc0.w_ring_norsz[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7444 a_10512_9545# _139_ a_10124_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7445 a_14499_13103# a_13717_13109# a_14415_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7446 _174_ a_10607_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7447 tdc1.w_ring_buf[17] a_23855_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7448 a_16025_14735# tdc0.r_ring_ctr[9] a_15919_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X7449 VPWR net35 a_24867_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7450 a_17475_13621# net32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7452 a_12621_10927# net49 tdc0.w_ring_int_norsz[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7453 a_8013_6575# tdc1.w_ring_norsz[15] a_7929_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7454 VGND net29 a_13735_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7455 VPWR net37 a_2511_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7456 a_18869_13647# a_18703_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7457 a_7009_12015# net20 tdc0.w_ring_norsz[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7459 a_16569_13109# a_16403_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7460 VPWR _067_ a_24029_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7461 a_4420_6031# a_3339_6031# a_4073_6273# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7462 VPWR a_7723_3829# a_7710_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7463 VGND net35 a_23395_14197# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7464 VPWR _075_ a_24849_13897# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7465 a_30537_7895# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X7466 tdc1.r_dly_store_ctr[14] a_7867_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7467 VPWR a_9374_6143# a_9301_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7469 a_12483_9661# a_11619_9295# a_12226_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7470 a_17746_12671# a_17578_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7471 VPWR a_14307_6549# a_14223_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7472 a_16301_12015# net23 tdc0.w_ring_norsz[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7473 VGND a_4866_8725# a_4824_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7474 VGND _033_ a_21413_15823# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7475 a_4328_12559# a_3247_12559# a_3981_12801# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7476 a_9677_7663# tdc1.r_dly_store_ring[15] a_9595_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7477 a_13637_7663# _076_ a_13839_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7478 VGND net24 a_13735_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X7479 tdc1.r_dly_store_ring[15] a_8695_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7480 tdc0.w_ring_buf[17] a_15483_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
R100 VGND net77 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7482 a_8686_15395# _152_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X7483 VGND _065_ a_18776_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X7485 a_17217_5487# tdc1.r_ring_ctr[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7486 _104_ a_24683_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X7487 VGND _166_ _025_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7488 VGND a_14139_14191# a_14307_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7489 a_3855_4943# a_3505_4943# a_3760_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7491 a_24646_10901# a_24478_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7492 VPWR net11 a_16669_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7493 uo_out[5] a_15504_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7494 a_11697_14191# tdc0.r_ring_ctr[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7495 a_5231_4631# _183_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X7496 a_24604_6953# a_24205_6581# a_24478_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7497 a_6388_6953# a_5989_6581# a_6262_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7499 a_21642_8029# a_21327_7895# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7501 a_24293_5865# a_23303_5493# a_24167_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7502 VGND net30 a_11987_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7503 _132_ a_9871_7369# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7504 VPWR a_9431_7387# a_9347_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7505 VPWR a_13035_4399# a_13203_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7506 a_13511_7895# _084_ a_13839_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7507 a_13035_4399# a_12337_4405# a_12778_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7508 a_28207_6575# a_27425_6581# a_28123_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7509 _116_ a_15023_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7510 VGND net15 tdc1.w_ring_norsz[31] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7511 a_19631_8867# a_19439_9111# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X7512 VGND a_6027_13915# a_5985_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7513 a_21445_8757# a_21279_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7514 a_7461_8757# a_7295_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7515 VGND a_15261_11445# _114_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7516 a_27242_10927# a_26995_11305# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7517 a_17501_11721# tdc0.w_ring_norsz[25] a_17417_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7518 a_25857_3855# a_24867_3855# a_25731_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7519 VGND tdc1.w_ring_norsz[14] tdc1.w_ring_int_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7520 tdc1.w_ring_norsz[16] tdc1.w_ring_int_norsz[16] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X7522 VPWR net30 a_11803_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7523 VGND net19 tdc1.w_ring_norsz[29] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7524 VPWR a_11398_6143# a_11325_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7525 a_23266_15645# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7527 uo_out[7] a_10124_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7529 a_5417_4917# tdc1.r_ring_ctr[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X7530 tdc0.r_dly_store_ring[6] a_8971_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7531 VGND net40 tdc1.w_ring_int_norsz[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7532 VPWR a_19959_15797# tdc0.r_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7533 a_9643_12724# tdc0.w_ring_norsz[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7534 VGND _086_ a_11067_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7535 tdc0.r_dly_store_ring[6] a_8971_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7536 a_4220_14735# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7538 a_5989_6581# a_5823_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7539 VPWR _082_ a_20083_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7540 VGND _120_ a_15025_7779# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7543 a_9213_8207# tdc1.w_ring_buf[23] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7544 a_16845_14735# tdc0.r_ring_ctr[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7545 tdc1.w_ring_buf[4] a_20083_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7546 a_9301_6397# a_8767_6031# a_9206_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7548 VGND _170_ _027_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7550 a_8270_7637# a_8102_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7551 VPWR a_24462_11989# a_24389_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7552 a_9963_5487# _077_ a_10045_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7553 VPWR a_4328_12559# a_4503_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7554 VGND net14 tdc1.w_ring_norsz[30] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7555 a_10018_11989# a_9850_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7556 VPWR net8 a_16679_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7557 VPWR net34 a_28087_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7558 a_17727_5487# a_17029_5493# a_17470_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7559 a_3981_12801# a_3763_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
R101 VGND uio_out[2] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7561 VGND a_12823_16073# _014_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7562 a_7263_15657# a_6817_15285# a_7167_15657# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7564 VPWR net26 a_3247_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7566 tdc1.w_ring_int_norsz[26] net71 a_27817_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7567 a_18243_8751# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7568 a_11045_10383# tdc0.r_dly_store_ring[24] a_10699_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7570 a_17033_9295# tdc1.w_ring_buf[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7572 a_25041_7369# _075_ a_25125_7369# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7573 VPWR a_6671_10651# a_6587_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7574 a_25306_13103# a_25033_13109# a_25221_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7576 VGND tdc1.r_ring_ctr[11] a_14471_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7577 a_16463_12533# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X7579 a_15420_9295# _117_ a_15504_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7580 a_25182_10383# _104_ a_25348_10633# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7581 a_17375_7637# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X7582 a_19535_7637# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X7583 VGND net34 a_24039_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7585 tdc0.w_ring_int_norsz[14] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7586 a_6364_14985# _159_ a_6273_14985# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.153 ps=1.3 w=1 l=0.15
X7587 VPWR a_19255_14735# net22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7588 a_15359_4943# a_14913_4943# a_15263_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7589 a_8362_4765# _060_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7590 a_9713_15645# _145_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X7591 a_3963_5309# a_3339_4943# a_3855_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7592 VGND a_27647_9813# a_27605_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7593 tdc0.r_dly_store_ring[9] a_18171_12827# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7594 tdc1.r_ring_ctr[5] a_12231_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7595 a_15627_14709# _152_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X7597 tdc0.w_ring_int_norsz[16] net43 a_6473_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7598 VGND net62 tdc1.w_ring_int_norsz[17] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7599 a_11533_3311# _169_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7600 VGND a_18171_8475# a_18129_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7601 VPWR a_22339_10535# tdc0.r_dly_store_ring[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7602 _157_ _152_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7603 a_11325_6397# a_10791_6031# a_11230_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7604 a_19946_16189# a_18869_15823# a_19784_15823# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7606 tdc0.r_dly_store_ctr[2] a_25899_14165# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7607 a_13905_13103# tdc0.w_ring_buf[29] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7609 a_27066_11204# a_26859_11145# a_27242_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7611 VGND net10 a_15023_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7613 VPWR tdc1.w_ring_norsz[11] a_27903_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7614 VGND a_12139_4007# _168_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X7615 VPWR net6 a_14794_9922# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X7616 net8 a_15023_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X7617 a_29403_8751# a_28621_8757# a_29319_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7618 _121_ a_15025_7779# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X7619 VGND _169_ _172_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7620 VPWR tdc1.r_dly_store_ring[17] a_25847_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7621 VGND _083_ a_21356_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
X7622 a_6756_12559# a_6357_12559# a_6630_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7623 VPWR a_17543_9661# a_17711_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7624 a_21813_12015# tdc0.w_ring_norsz[11] a_21729_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7625 a_18249_12015# tdc0.w_ring_norsz[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7627 VGND _190_ a_14197_10389# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7628 VPWR tdc0.w_dly_stop[5] a_3799_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7629 _005_ _162_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7631 VPWR tdc1.w_ring_norsz[25] a_28271_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7633 a_13725_12015# net23 tdc0.w_ring_norsz[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7635 VGND a_25163_8725# a_25121_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7636 a_7055_9839# a_6191_9845# a_6798_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7637 VPWR a_22903_14709# a_22890_15101# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7638 tdc0.w_ring_buf[8] a_11435_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7639 a_6093_14511# tdc0.r_ring_ctr[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7640 VGND a_6119_7387# a_6077_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7641 a_17727_5487# a_16863_5493# a_17470_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7643 a_10045_5487# tdc1.r_dly_store_ctr[14] a_9963_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7645 VGND _150_ a_10393_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7646 a_9022_5309# a_8749_4943# a_8937_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7647 _146_ a_10363_15617# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X7648 VGND a_28215_5487# a_28383_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7650 a_13788_3677# _030_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7652 a_15207_10927# _074_ a_15289_11247# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7653 a_17785_11721# tdc0.w_ring_int_norsz[25] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7654 a_9058_16189# a_8971_15965# a_8654_16075# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X7655 VGND tdc0.w_ring_norsz[3] a_23763_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7656 a_24987_6575# a_24205_6581# a_24903_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
R102 VPWR tdc0.g_ring3[23].stg01_50.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7658 VPWR tdc1.w_ring_int_norsz[0] a_6743_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7659 a_9690_16189# a_8971_15965# a_9127_16060# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X7660 VPWR a_3115_9813# net26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7662 _195_ a_18703_14735# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7663 a_13511_7895# tdc1.r_dly_store_ring[8] a_13637_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X7664 VPWR a_12651_9563# a_12567_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7665 a_14101_3285# a_13883_3689# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7666 VPWR tdc1.w_ring_int_norsz[4] a_23009_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7667 VPWR a_29955_8983# _073_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7668 _110_ a_12447_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7669 a_10245_3311# tdc1.r_ring_ctr[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7670 a_13809_14191# a_13275_14197# a_13714_14191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7671 a_24738_8725# a_24570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7672 VGND _086_ a_5773_9622# VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X7673 VPWR tdc0.w_ring_int_norsz[21] a_16753_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7674 a_4725_12015# tdc0.w_ring_norsz[16] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7675 _022_ _184_ a_2769_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X7676 tdc0.w_ring_int_norsz[18] tdc0.w_ring_norsz[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7679 a_16396_9111# a_16209_8751# a_16309_8867# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X7681 a_5767_11837# a_5069_11471# a_5510_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7682 tdc1.w_dly_stop[1] a_26615_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7683 VPWR net36 a_29007_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7684 uo_out[1] a_24849_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7685 a_4577_14735# a_4533_14977# a_4411_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X7686 VPWR a_15351_14423# _002_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X7687 _091_ a_26431_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7688 a_23201_10927# net41 tdc0.w_ring_int_norsz[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7689 a_27329_12559# tdc0.r_dly_store_ring[26] a_26891_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7691 a_12426_7663# a_12153_7669# a_12341_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7692 a_4613_8751# tdc1.w_ring_buf[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7693 VGND a_19310_13759# a_19268_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7694 a_10589_5309# a_10055_4943# a_10494_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7695 a_27437_8751# tdc1.w_ring_norsz[26] a_27353_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7696 tdc0.w_ring_norsz[17] tdc0.w_ring_int_norsz[17] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7697 VGND a_17010_13077# a_16968_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7700 a_19613_11721# net22 tdc0.w_ring_norsz[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7701 _149_ tdc0.r_ring_ctr[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7702 a_12231_2741# a_12056_2767# a_12410_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7703 a_19741_8235# _080_ a_19655_8235# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7704 a_19329_9839# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X7706 a_22143_9839# a_21445_9845# a_21886_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7707 a_21813_13647# a_21647_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7708 a_24297_8757# a_24131_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7710 tdc1.w_ring_int_norsz[28] net73 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7711 VGND tdc1.w_ring_norsz[27] a_28179_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7712 VGND a_20931_11739# a_20889_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7713 VPWR tdc0.w_ring_int_norsz[15] a_7093_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7714 VPWR net28 a_8399_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7715 a_17267_13103# a_16569_13109# a_17010_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7716 uo_out[3] a_25348_10633# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X7718 a_24738_8725# a_24570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7719 tdc0.r_dly_store_ring[28] a_19459_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7720 a_19237_3317# a_19071_3317# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7721 tdc1.r_dly_store_ring[1] a_24151_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7722 VPWR a_17229_4097# a_17119_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X7723 a_4411_14735# a_3965_14735# a_4315_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7724 a_17475_13621# net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7725 VGND tdc1.w_ring_int_norsz[14] tdc1.w_ring_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7726 VPWR _195_ _032_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7727 a_17283_14709# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X7728 VPWR a_21223_5309# a_21391_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7729 tdc1.r_ring_ctr[12] a_8183_4703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7730 VGND a_5055_14709# tdc0.r_ring_ctr[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7731 a_14983_14165# tdc0.w_ring_buf[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X7733 a_19651_14013# a_18869_13647# a_19567_14013# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7734 tdc1.r_dly_store_ctr[4] a_25899_4123# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7736 a_5349_13647# tdc0.r_ring_ctr[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7737 VGND tdc0.w_ring_norsz[22] a_10975_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7738 tdc1.w_ring_norsz[1] net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7739 _075_ a_14011_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X7740 VPWR tdc0.r_dly_store_ring[13] a_15479_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X7741 VPWR net29 a_10975_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7742 VGND net8 a_18611_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7743 _176_ tdc1.r_ring_ctr[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7744 VGND a_9006_7231# a_8964_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7746 VPWR a_20487_12925# a_20655_12827# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7747 a_20690_6143# a_20522_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7749 a_11241_7663# net16 tdc1.w_ring_norsz[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7750 a_17581_14197# a_17415_14197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7751 a_11601_12809# tdc0.r_dly_store_ctr[6] a_11517_12809# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7752 a_20065_11471# a_19899_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7753 VPWR a_11839_13103# a_12007_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7754 VPWR a_25348_10633# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7755 VGND a_15719_10357# net25 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X7757 _041_ _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7758 VPWR _186_ a_13707_8867# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
R103 tdc0.g_ring3[21].stg01_48.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7759 VPWR tdc0.w_ring_norsz[21] a_12621_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7760 a_27491_5108# tdc1.w_dly_stop[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7761 a_2724_10927# a_2287_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7762 VGND a_11839_13103# a_12007_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7763 tdc1.r_ring_ctr[6] a_9379_3615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7764 VGND net21 tdc0.w_ring_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7765 VGND a_17543_9661# a_17711_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7766 a_26785_12015# tdc0.w_ring_buf[18] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7767 VGND a_9079_14191# a_9247_14165# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7768 a_17578_8573# a_17305_8207# a_17493_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7769 VPWR a_4295_10749# a_4463_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7771 VGND a_19735_5211# a_19693_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7772 a_14448_3689# a_13367_3317# a_14101_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7775 a_2807_11169# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7776 a_18697_12015# tdc0.w_ring_norsz[10] a_18613_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7777 tdc1.r_dly_store_ctr[11] a_17895_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7779 a_14059_8983# a_14332_8983# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7781 VGND net8 a_14747_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7782 a_16385_3311# tdc1.r_ring_ctr[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7783 a_19375_10927# a_18593_10933# a_19291_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7784 tdc1.r_dly_store_ring[29] a_16331_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7785 VGND net23 a_19255_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X7787 a_20257_13103# _087_ a_20175_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7788 VGND a_4111_9661# a_4279_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7789 a_7385_15253# a_7167_15657# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7790 VGND a_28538_12292# a_28467_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7791 VGND net9 a_11619_14735# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7792 VPWR a_8235_13077# a_8151_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7793 VGND a_21912_6575# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7794 VGND a_25899_4123# a_25857_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7797 VGND a_28951_7663# a_29119_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7798 a_24845_12393# a_23855_12021# a_24719_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7799 net40 a_27351_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X7802 _051_ _196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 uio_in[6] VGND 0.182f
C1 uio_in[7] VGND 0.182f
C2 uio_in[4] VGND 0.182f
C3 uio_in[3] VGND 0.182f
C4 uio_in[2] VGND 0.182f
C5 uio_in[1] VGND 0.182f
C6 uio_in[0] VGND 0.182f
C7 ui_in[7] VGND 0.182f
C8 ui_in[6] VGND 0.182f
C9 rst_n VGND 0.182f
C10 ena VGND 0.182f
C11 clk VGND 0.182f
C12 uio_in[5] VGND 0.182f
C13 uio_oe[6] VGND 0.917f
C14 ui_in[3] VGND 0.831f
C15 ui_in[4] VGND 0.83f
C16 ui_in[5] VGND 0.743f
C17 uio_out[6] VGND 0.917f
C18 uio_out[4] VGND 0.917f
C19 uo_out[4] VGND 5.03f
C20 ui_in[0] VGND 1.12f
C21 uo_out[5] VGND 5.04f
C22 uo_out[0] VGND 4.44f
C23 uo_out[7] VGND 5.13f
C24 uo_out[1] VGND 3.47f
C25 uo_out[3] VGND 3.29f
C26 ui_in[2] VGND 0.98f
C27 uo_out[2] VGND 2.97f
C28 uo_out[6] VGND 4.14f
C29 ui_in[1] VGND 0.899f
C30 uio_out[5] VGND 1.13f
C31 uio_oe[4] VGND 1.09f
C32 uio_out[1] VGND 1.09f
C33 uio_oe[5] VGND 1.09f
C34 uio_oe[0] VGND 1.09f
C35 uio_oe[1] VGND 1.09f
C36 uio_oe[2] VGND 1.09f
C37 uio_out[7] VGND 1.09f
C38 uio_oe[3] VGND 1.08f
C39 uio_out[3] VGND 1.09f
C40 uio_oe[7] VGND 1.09f
C41 uio_out[2] VGND 1.09f
C42 uio_out[0] VGND 1.09f
C43 VPWR VGND 2.41p
C44 tt_um_hpretl_tt06_tdc_v2_84.HI VGND 0.415f $ **FLOATING
C45 tt_um_hpretl_tt06_tdc_v2_92.HI VGND 0.415f $ **FLOATING
C46 a_16913_756# VGND 0.524f $ **FLOATING
C47 a_16219_591# VGND 0.524f $ **FLOATING
C48 a_15575_591# VGND 0.524f $ **FLOATING
C49 tt_um_hpretl_tt06_tdc_v2_90.HI VGND 0.415f $ **FLOATING
C50 a_20985_3017# VGND 0.219f $ **FLOATING
C51 a_17303_3133# VGND 0.168f $ **FLOATING
C52 a_17100_2767# VGND 0.259f $ **FLOATING
C53 a_20735_3017# VGND 0.684f $ **FLOATING
C54 a_17760_2767# VGND 0.736f $ **FLOATING
C55 a_17935_2741# VGND 1.13f $ **FLOATING
C56 a_17195_2767# VGND 0.714f $ **FLOATING
C57 _052_ VGND 1.68f $ **FLOATING
C58 a_17413_3009# VGND 0.653f $ **FLOATING
C59 a_16845_2767# VGND 1.57f $ **FLOATING
C60 a_16679_2767# VGND 1.92f $ **FLOATING
C61 a_11599_3133# VGND 0.168f $ **FLOATING
C62 a_11396_2767# VGND 0.259f $ **FLOATING
C63 a_12056_2767# VGND 0.736f $ **FLOATING
C64 a_12231_2741# VGND 0.971f $ **FLOATING
C65 a_11491_2767# VGND 0.714f $ **FLOATING
C66 _053_ VGND 1.6f $ **FLOATING
C67 a_11709_3009# VGND 0.653f $ **FLOATING
C68 a_11141_2767# VGND 1.57f $ **FLOATING
C69 a_10975_2767# VGND 1.92f $ **FLOATING
C70 a_22179_3311# VGND 0.168f $ **FLOATING
C71 a_21976_3677# VGND 0.259f $ **FLOATING
C72 a_19695_3311# VGND 0.168f $ **FLOATING
C73 a_16385_3311# VGND 0.219f $ **FLOATING
C74 a_19492_3677# VGND 0.259f $ **FLOATING
C75 _026_ VGND 1.33f $ **FLOATING
C76 a_13991_3311# VGND 0.168f $ **FLOATING
C77 a_12981_3311# VGND 0.219f $ **FLOATING
C78 a_11895_3311# VGND 0.238f $ **FLOATING
C79 a_13788_3677# VGND 0.259f $ **FLOATING
C80 _027_ VGND 1.27f $ **FLOATING
C81 a_8747_3311# VGND 0.168f $ **FLOATING
C82 a_8544_3677# VGND 0.259f $ **FLOATING
C83 a_22636_3689# VGND 0.736f $ **FLOATING
C84 a_22811_3615# VGND 1.13f $ **FLOATING
C85 a_22071_3689# VGND 0.714f $ **FLOATING
C86 _049_ VGND 1.64f $ **FLOATING
C87 a_22289_3285# VGND 0.653f $ **FLOATING
C88 a_21721_3317# VGND 1.57f $ **FLOATING
C89 _023_ VGND 1.39f $ **FLOATING
C90 a_21555_3317# VGND 1.92f $ **FLOATING
C91 a_20152_3689# VGND 0.736f $ **FLOATING
C92 a_20327_3615# VGND 1.54f $ **FLOATING
C93 a_19587_3689# VGND 0.714f $ **FLOATING
C94 _048_ VGND 1.74f $ **FLOATING
C95 a_19805_3285# VGND 0.653f $ **FLOATING
C96 a_19237_3317# VGND 1.57f $ **FLOATING
C97 _016_ VGND 1.04f $ **FLOATING
C98 a_19071_3317# VGND 1.92f $ **FLOATING
C99 a_16135_3311# VGND 0.684f $ **FLOATING
C100 a_14448_3689# VGND 0.736f $ **FLOATING
C101 a_14623_3615# VGND 1.13f $ **FLOATING
C102 a_13883_3689# VGND 0.714f $ **FLOATING
C103 _056_ VGND 1.64f $ **FLOATING
C104 a_14101_3285# VGND 0.653f $ **FLOATING
C105 a_13533_3317# VGND 1.57f $ **FLOATING
C106 _030_ VGND 1.1f $ **FLOATING
C107 a_13367_3317# VGND 1.92f $ **FLOATING
C108 a_12731_3311# VGND 0.684f $ **FLOATING
C109 _170_ VGND 0.861f $ **FLOATING
C110 a_11035_3543# VGND 0.56f $ **FLOATING
C111 _172_ VGND 0.686f $ **FLOATING
C112 _169_ VGND 1.38f $ **FLOATING
C113 a_9204_3689# VGND 0.736f $ **FLOATING
C114 a_9379_3615# VGND 0.971f $ **FLOATING
C115 a_8639_3689# VGND 0.714f $ **FLOATING
C116 _054_ VGND 1.69f $ **FLOATING
C117 a_8857_3285# VGND 0.653f $ **FLOATING
C118 a_8289_3317# VGND 1.57f $ **FLOATING
C119 _028_ VGND 1.76f $ **FLOATING
C120 a_8123_3317# VGND 1.92f $ **FLOATING
C121 a_25221_3855# VGND 0.23f $ **FLOATING
C122 a_25731_4221# VGND 0.609f $ **FLOATING
C123 a_25899_4123# VGND 0.817f $ **FLOATING
C124 a_25306_4221# VGND 0.626f $ **FLOATING
C125 a_25474_3967# VGND 0.581f $ **FLOATING
C126 a_25033_3855# VGND 1.43f $ **FLOATING
C127 a_24867_3855# VGND 1.81f $ **FLOATING
C128 a_22547_4221# VGND 0.168f $ **FLOATING
C129 a_22344_3855# VGND 0.259f $ **FLOATING
C130 a_23004_3855# VGND 0.736f $ **FLOATING
C131 a_23179_3829# VGND 0.971f $ **FLOATING
C132 a_22439_3855# VGND 0.714f $ **FLOATING
C133 a_22657_4097# VGND 0.653f $ **FLOATING
C134 a_22089_3855# VGND 1.57f $ **FLOATING
C135 a_21923_3855# VGND 1.92f $ **FLOATING
C136 a_20445_4105# VGND 0.238f $ **FLOATING
C137 a_15189_3855# VGND 0.211f $ **FLOATING
C138 a_17119_4221# VGND 0.168f $ **FLOATING
C139 a_16916_3855# VGND 0.259f $ **FLOATING
C140 _163_ VGND 0.794f $ **FLOATING
C141 a_17576_3855# VGND 0.736f $ **FLOATING
C142 a_17751_3829# VGND 1.13f $ **FLOATING
C143 a_17011_3855# VGND 0.714f $ **FLOATING
C144 _057_ VGND 1.76f $ **FLOATING
C145 a_17229_4097# VGND 0.653f $ **FLOATING
C146 a_16661_3855# VGND 1.57f $ **FLOATING
C147 a_16495_3855# VGND 1.92f $ **FLOATING
C148 _031_ VGND 1.44f $ **FLOATING
C149 tdc1.r_ring_ctr[4] VGND 8.54f $ **FLOATING
C150 a_9740_3855# VGND 0.205f $ **FLOATING
C151 a_7091_4221# VGND 0.168f $ **FLOATING
C152 a_6888_3855# VGND 0.259f $ **FLOATING
C153 a_14951_3855# VGND 0.706f $ **FLOATING
C154 _176_ VGND 1.17f $ **FLOATING
C155 a_12139_4007# VGND 0.56f $ **FLOATING
C156 a_11115_4007# VGND 0.619f $ **FLOATING
C157 a_10607_3855# VGND 0.619f $ **FLOATING
C158 _171_ VGND 1.85f $ **FLOATING
C159 a_9514_3901# VGND 0.443f $ **FLOATING
C160 a_9371_4007# VGND 0.65f $ **FLOATING
C161 a_8399_3855# VGND 0.988f $ **FLOATING
C162 a_7548_3855# VGND 0.736f $ **FLOATING
C163 a_7723_3829# VGND 0.971f $ **FLOATING
C164 a_6983_3855# VGND 0.714f $ **FLOATING
C165 _055_ VGND 1.94f $ **FLOATING
C166 a_7201_4097# VGND 0.653f $ **FLOATING
C167 a_6633_3855# VGND 1.57f $ **FLOATING
C168 _029_ VGND 2.01f $ **FLOATING
C169 a_6467_3855# VGND 1.92f $ **FLOATING
C170 a_23841_4399# VGND 0.23f $ **FLOATING
C171 _051_ VGND 1.69f $ **FLOATING
C172 _025_ VGND 1.27f $ **FLOATING
C173 a_19235_4399# VGND 0.168f $ **FLOATING
C174 a_19032_4765# VGND 0.259f $ **FLOATING
C175 a_17303_4399# VGND 0.168f $ **FLOATING
C176 a_15649_4399# VGND 0.219f $ **FLOATING
C177 a_17100_4765# VGND 0.259f $ **FLOATING
C178 a_12525_4399# VGND 0.23f $ **FLOATING
C179 a_7551_4399# VGND 0.168f $ **FLOATING
C180 a_7348_4765# VGND 0.259f $ **FLOATING
C181 a_5449_4719# VGND 0.171f $ **FLOATING
C182 a_24351_4399# VGND 0.609f $ **FLOATING
C183 a_24519_4373# VGND 0.817f $ **FLOATING
C184 a_23926_4399# VGND 0.626f $ **FLOATING
C185 a_24094_4373# VGND 0.581f $ **FLOATING
C186 a_23653_4405# VGND 1.43f $ **FLOATING
C187 a_23487_4405# VGND 1.81f $ **FLOATING
C188 _196_ VGND 14.5f $ **FLOATING
C189 _167_ VGND 0.686f $ **FLOATING
C190 _164_ VGND 1.72f $ **FLOATING
C191 a_21923_4399# VGND 0.698f $ **FLOATING
C192 _165_ VGND 0.663f $ **FLOATING
C193 a_21279_4765# VGND 0.729f $ **FLOATING
C194 tdc1.r_ring_ctr[3] VGND 2.75f $ **FLOATING
C195 a_20635_4512# VGND 0.619f $ **FLOATING
C196 a_19692_4777# VGND 0.736f $ **FLOATING
C197 a_19867_4703# VGND 0.971f $ **FLOATING
C198 a_19127_4777# VGND 0.714f $ **FLOATING
C199 _050_ VGND 1.74f $ **FLOATING
C200 a_19345_4373# VGND 0.653f $ **FLOATING
C201 a_18777_4405# VGND 1.57f $ **FLOATING
C202 _024_ VGND 1.98f $ **FLOATING
C203 a_18611_4405# VGND 1.92f $ **FLOATING
C204 a_17760_4777# VGND 0.736f $ **FLOATING
C205 a_17935_4703# VGND 0.971f $ **FLOATING
C206 a_17195_4777# VGND 0.714f $ **FLOATING
C207 a_17413_4373# VGND 0.653f $ **FLOATING
C208 a_16845_4405# VGND 1.57f $ **FLOATING
C209 _017_ VGND 1.43f $ **FLOATING
C210 a_16679_4405# VGND 1.92f $ **FLOATING
C211 a_15399_4399# VGND 0.684f $ **FLOATING
C212 _177_ VGND 1.39f $ **FLOATING
C213 a_14431_4373# VGND 0.729f $ **FLOATING
C214 a_13919_4512# VGND 0.619f $ **FLOATING
C215 _175_ VGND 7.7f $ **FLOATING
C216 a_13035_4399# VGND 0.609f $ **FLOATING
C217 a_13203_4373# VGND 0.817f $ **FLOATING
C218 a_12610_4399# VGND 0.626f $ **FLOATING
C219 a_12778_4373# VGND 0.581f $ **FLOATING
C220 a_12337_4405# VGND 1.43f $ **FLOATING
C221 tdc1.r_ring_ctr[5] VGND 2.59f $ **FLOATING
C222 a_12171_4405# VGND 1.81f $ **FLOATING
C223 a_11067_4399# VGND 0.698f $ **FLOATING
C224 _174_ VGND 0.924f $ **FLOATING
C225 _166_ VGND 10.3f $ **FLOATING
C226 _168_ VGND 3.16f $ **FLOATING
C227 _173_ VGND 1.7f $ **FLOATING
C228 a_10291_4373# VGND 0.729f $ **FLOATING
C229 a_9811_4737# VGND 0.56f $ **FLOATING
C230 a_9103_4659# VGND 1.2f $ **FLOATING
C231 a_8008_4777# VGND 0.736f $ **FLOATING
C232 a_8183_4703# VGND 1.54f $ **FLOATING
C233 a_7443_4777# VGND 0.714f $ **FLOATING
C234 a_7661_4373# VGND 0.653f $ **FLOATING
C235 a_7093_4405# VGND 1.57f $ **FLOATING
C236 a_6927_4405# VGND 1.92f $ **FLOATING
C237 a_5231_4631# VGND 0.546f $ **FLOATING
C238 a_20713_4943# VGND 0.23f $ **FLOATING
C239 tdc1.w_dly_stop[4] VGND 0.879f $ **FLOATING
C240 a_27769_5108# VGND 0.524f $ **FLOATING
C241 tdc1.w_dly_stop[2] VGND 0.881f $ **FLOATING
C242 a_27491_5108# VGND 0.524f $ **FLOATING
C243 a_27167_4943# VGND 0.524f $ **FLOATING
C244 tdc1.w_dly_stop[3] VGND 0.761f $ **FLOATING
C245 a_26891_4943# VGND 0.524f $ **FLOATING
C246 tdc1.w_dly_stop[1] VGND 0.683f $ **FLOATING
C247 a_26615_4943# VGND 0.524f $ **FLOATING
C248 a_21223_5309# VGND 0.609f $ **FLOATING
C249 a_21391_5211# VGND 0.817f $ **FLOATING
C250 a_20798_5309# VGND 0.626f $ **FLOATING
C251 a_20966_5055# VGND 0.581f $ **FLOATING
C252 a_20525_4943# VGND 1.43f $ **FLOATING
C253 tdc1.r_ring_ctr[2] VGND 2.95f $ **FLOATING
C254 a_20359_4943# VGND 1.81f $ **FLOATING
C255 a_19057_4943# VGND 0.23f $ **FLOATING
C256 a_19567_5309# VGND 0.609f $ **FLOATING
C257 a_19735_5211# VGND 0.817f $ **FLOATING
C258 a_19142_5309# VGND 0.626f $ **FLOATING
C259 a_19310_5055# VGND 0.581f $ **FLOATING
C260 a_18869_4943# VGND 1.43f $ **FLOATING
C261 a_18703_4943# VGND 1.81f $ **FLOATING
C262 _058_ VGND 1.66f $ **FLOATING
C263 a_15371_5309# VGND 0.168f $ **FLOATING
C264 a_15168_4943# VGND 0.259f $ **FLOATING
C265 a_15828_4943# VGND 0.736f $ **FLOATING
C266 a_16003_4917# VGND 0.971f $ **FLOATING
C267 a_15263_4943# VGND 0.714f $ **FLOATING
C268 a_15481_5185# VGND 0.653f $ **FLOATING
C269 a_14913_4943# VGND 1.57f $ **FLOATING
C270 a_14747_4943# VGND 1.92f $ **FLOATING
C271 _179_ VGND 3.1f $ **FLOATING
C272 a_12157_4943# VGND 0.23f $ **FLOATING
C273 tdc1.r_ring_ctr[10] VGND 4.35f $ **FLOATING
C274 a_14155_4917# VGND 0.729f $ **FLOATING
C275 a_12667_5309# VGND 0.609f $ **FLOATING
C276 a_12835_5211# VGND 0.817f $ **FLOATING
C277 a_12242_5309# VGND 0.626f $ **FLOATING
C278 a_12410_5055# VGND 0.581f $ **FLOATING
C279 a_11969_4943# VGND 1.43f $ **FLOATING
C280 tdc1.r_ring_ctr[8] VGND 6.3f $ **FLOATING
C281 a_11803_4943# VGND 1.81f $ **FLOATING
C282 a_10409_4943# VGND 0.23f $ **FLOATING
C283 a_10919_5309# VGND 0.609f $ **FLOATING
C284 a_11087_5211# VGND 0.817f $ **FLOATING
C285 a_10494_5309# VGND 0.626f $ **FLOATING
C286 a_10662_5055# VGND 0.581f $ **FLOATING
C287 a_10221_4943# VGND 1.43f $ **FLOATING
C288 tdc1.r_ring_ctr[6] VGND 3.92f $ **FLOATING
C289 a_10055_4943# VGND 1.81f $ **FLOATING
C290 a_8937_4943# VGND 0.23f $ **FLOATING
C291 a_9447_5309# VGND 0.609f $ **FLOATING
C292 a_9615_5211# VGND 0.817f $ **FLOATING
C293 a_9022_5309# VGND 0.626f $ **FLOATING
C294 a_9190_5055# VGND 0.581f $ **FLOATING
C295 a_8749_4943# VGND 1.43f $ **FLOATING
C296 tdc1.r_ring_ctr[7] VGND 2.92f $ **FLOATING
C297 a_8583_4943# VGND 1.81f $ **FLOATING
C298 _060_ VGND 1.66f $ **FLOATING
C299 _019_ VGND 1.37f $ **FLOATING
C300 a_6541_5193# VGND 0.219f $ **FLOATING
C301 _182_ VGND 1.07f $ **FLOATING
C302 a_5635_5193# VGND 0.253f $ **FLOATING
C303 _183_ VGND 0.762f $ **FLOATING
C304 a_3963_5309# VGND 0.168f $ **FLOATING
C305 a_3760_4943# VGND 0.259f $ **FLOATING
C306 a_6980_4917# VGND 0.648f $ **FLOATING
C307 a_6291_5193# VGND 0.684f $ **FLOATING
C308 a_5417_4917# VGND 0.55f $ **FLOATING
C309 a_4420_4943# VGND 0.736f $ **FLOATING
C310 a_4595_4917# VGND 0.971f $ **FLOATING
C311 a_3855_4943# VGND 0.714f $ **FLOATING
C312 _061_ VGND 1.66f $ **FLOATING
C313 a_4073_5185# VGND 0.653f $ **FLOATING
C314 a_3505_4943# VGND 1.57f $ **FLOATING
C315 _020_ VGND 1.74f $ **FLOATING
C316 a_3339_4943# VGND 1.92f $ **FLOATING
C317 a_27705_5487# VGND 0.23f $ **FLOATING
C318 a_25129_5487# VGND 0.23f $ **FLOATING
C319 a_23657_5487# VGND 0.23f $ **FLOATING
C320 a_22185_5487# VGND 0.23f $ **FLOATING
C321 a_19793_5487# VGND 0.23f $ **FLOATING
C322 a_17217_5487# VGND 0.23f $ **FLOATING
C323 _059_ VGND 1.71f $ **FLOATING
C324 net8 VGND 9.95f $ **FLOATING
C325 _018_ VGND 1.11f $ **FLOATING
C326 a_14471_5807# VGND 0.171f $ **FLOATING
C327 a_13797_5865# VGND 0.23f $ **FLOATING
C328 a_10045_5487# VGND 0.206f $ **FLOATING
C329 a_5907_5487# VGND 0.184f $ **FLOATING
C330 a_28215_5487# VGND 0.609f $ **FLOATING
C331 a_28383_5461# VGND 0.817f $ **FLOATING
C332 a_27790_5487# VGND 0.626f $ **FLOATING
C333 a_27958_5461# VGND 0.581f $ **FLOATING
C334 a_27517_5493# VGND 1.43f $ **FLOATING
C335 tdc1.w_ring_buf[28] VGND 0.872f $ **FLOATING
C336 a_27351_5493# VGND 1.81f $ **FLOATING
C337 a_27075_5487# VGND 0.524f $ **FLOATING
C338 a_25639_5487# VGND 0.609f $ **FLOATING
C339 a_25807_5461# VGND 0.817f $ **FLOATING
C340 a_25214_5487# VGND 0.626f $ **FLOATING
C341 a_25382_5461# VGND 0.581f $ **FLOATING
C342 a_24941_5493# VGND 1.43f $ **FLOATING
C343 a_24775_5493# VGND 1.81f $ **FLOATING
C344 a_24167_5487# VGND 0.609f $ **FLOATING
C345 a_24335_5461# VGND 0.817f $ **FLOATING
C346 a_23742_5487# VGND 0.626f $ **FLOATING
C347 a_23910_5461# VGND 0.581f $ **FLOATING
C348 a_23469_5493# VGND 1.43f $ **FLOATING
C349 tdc1.r_ring_ctr[1] VGND 6.07f $ **FLOATING
C350 a_23303_5493# VGND 1.81f $ **FLOATING
C351 a_22695_5487# VGND 0.609f $ **FLOATING
C352 a_22863_5461# VGND 0.817f $ **FLOATING
C353 a_22270_5487# VGND 0.626f $ **FLOATING
C354 a_22438_5461# VGND 0.581f $ **FLOATING
C355 a_21997_5493# VGND 1.43f $ **FLOATING
C356 tdc1.r_ring_ctr[9] VGND 7.7f $ **FLOATING
C357 a_21831_5493# VGND 1.81f $ **FLOATING
C358 a_20303_5487# VGND 0.609f $ **FLOATING
C359 a_20471_5461# VGND 0.817f $ **FLOATING
C360 a_19878_5487# VGND 0.626f $ **FLOATING
C361 a_20046_5461# VGND 0.581f $ **FLOATING
C362 a_19605_5493# VGND 1.43f $ **FLOATING
C363 a_19439_5493# VGND 1.81f $ **FLOATING
C364 a_17727_5487# VGND 0.609f $ **FLOATING
C365 a_17895_5461# VGND 0.817f $ **FLOATING
C366 a_17302_5487# VGND 0.626f $ **FLOATING
C367 a_17470_5461# VGND 0.581f $ **FLOATING
C368 a_17029_5493# VGND 1.43f $ **FLOATING
C369 a_16863_5493# VGND 1.81f $ **FLOATING
C370 a_15023_5487# VGND 0.698f $ **FLOATING
C371 a_14644_5487# VGND 0.546f $ **FLOATING
C372 _180_ VGND 5.78f $ **FLOATING
C373 _178_ VGND 1.1f $ **FLOATING
C374 tdc1.r_ring_ctr[11] VGND 3.52f $ **FLOATING
C375 tdc1.r_ring_ctr[0] VGND 8.73f $ **FLOATING
C376 a_13379_5865# VGND 0.581f $ **FLOATING
C377 a_13450_5764# VGND 0.626f $ **FLOATING
C378 a_13250_5609# VGND 1.43f $ **FLOATING
C379 a_13243_5705# VGND 1.81f $ **FLOATING
C380 a_12959_5719# VGND 0.609f $ **FLOATING
C381 a_12863_5719# VGND 0.817f $ **FLOATING
C382 a_9963_5487# VGND 0.804f $ **FLOATING
C383 _185_ VGND 1.53f $ **FLOATING
C384 tdc1.g_ring3[29].stg01_74.HI VGND 0.415f $ **FLOATING
C385 a_27167_6031# VGND 0.524f $ **FLOATING
C386 a_26329_6281# VGND 0.206f $ **FLOATING
C387 a_24213_6281# VGND 0.206f $ **FLOATING
C388 a_26247_6281# VGND 0.804f $ **FLOATING
C389 tdc1.r_dly_store_ring[20] VGND 0.943f $ **FLOATING
C390 tdc1.r_dly_store_ctr[4] VGND 1.53f $ **FLOATING
C391 net74 VGND 1.36f $ **FLOATING
C392 a_24131_6281# VGND 0.804f $ **FLOATING
C393 tdc1.r_dly_store_ctr[1] VGND 0.904f $ **FLOATING
C394 tdc1.r_dly_store_ctr[9] VGND 1.16f $ **FLOATING
C395 a_23855_6031# VGND 0.524f $ **FLOATING
C396 net65 VGND 0.822f $ **FLOATING
C397 tdc1.g_ring3[20].stg01_65.HI VGND 0.415f $ **FLOATING
C398 tdc1.w_ring_buf[20] VGND 1.72f $ **FLOATING
C399 a_22935_6031# VGND 0.524f $ **FLOATING
C400 net66 VGND 0.822f $ **FLOATING
C401 tdc1.g_ring3[21].stg01_66.HI VGND 0.415f $ **FLOATING
C402 a_20437_6031# VGND 0.23f $ **FLOATING
C403 a_20947_6397# VGND 0.609f $ **FLOATING
C404 a_21115_6299# VGND 0.817f $ **FLOATING
C405 a_20522_6397# VGND 0.626f $ **FLOATING
C406 a_20690_6143# VGND 0.581f $ **FLOATING
C407 a_20249_6031# VGND 1.43f $ **FLOATING
C408 a_20083_6031# VGND 1.81f $ **FLOATING
C409 a_15653_6031# VGND 0.23f $ **FLOATING
C410 tdc1.w_ring_int_norsz[29] VGND 3.55f $ **FLOATING
C411 a_16163_6397# VGND 0.609f $ **FLOATING
C412 a_16331_6299# VGND 0.817f $ **FLOATING
C413 a_15738_6397# VGND 0.626f $ **FLOATING
C414 a_15906_6143# VGND 0.581f $ **FLOATING
C415 a_15465_6031# VGND 1.43f $ **FLOATING
C416 a_15299_6031# VGND 1.81f $ **FLOATING
C417 tdc1.w_ring_buf[29] VGND 1.03f $ **FLOATING
C418 a_12437_6281# VGND 0.206f $ **FLOATING
C419 a_11145_6031# VGND 0.23f $ **FLOATING
C420 a_15023_6031# VGND 0.524f $ **FLOATING
C421 tdc1.w_ring_int_norsz[30] VGND 0.722f $ **FLOATING
C422 tdc1.w_ring_norsz[29] VGND 3.75f $ **FLOATING
C423 a_13599_6196# VGND 0.524f $ **FLOATING
C424 tdc1.w_ring_norsz[13] VGND 3.98f $ **FLOATING
C425 tdc1.r_dly_store_ctr[6] VGND 1.58f $ **FLOATING
C426 tdc1.r_dly_store_ring[22] VGND 0.76f $ **FLOATING
C427 a_12291_6183# VGND 0.804f $ **FLOATING
C428 a_11655_6397# VGND 0.609f $ **FLOATING
C429 a_11823_6299# VGND 0.817f $ **FLOATING
C430 a_11230_6397# VGND 0.626f $ **FLOATING
C431 a_11398_6143# VGND 0.581f $ **FLOATING
C432 a_10957_6031# VGND 1.43f $ **FLOATING
C433 a_10791_6031# VGND 1.81f $ **FLOATING
C434 tdc1.r_dly_store_ring[30] VGND 0.831f $ **FLOATING
C435 a_9121_6031# VGND 0.23f $ **FLOATING
C436 a_9631_6397# VGND 0.609f $ **FLOATING
C437 a_9799_6299# VGND 0.817f $ **FLOATING
C438 a_9206_6397# VGND 0.626f $ **FLOATING
C439 a_9374_6143# VGND 0.581f $ **FLOATING
C440 a_8933_6031# VGND 1.43f $ **FLOATING
C441 a_8767_6031# VGND 1.81f $ **FLOATING
C442 tdc1.w_ring_buf[30] VGND 0.872f $ **FLOATING
C443 tdc1.r_dly_store_ctr[14] VGND 1.53f $ **FLOATING
C444 a_7189_6031# VGND 0.23f $ **FLOATING
C445 a_8491_6031# VGND 0.524f $ **FLOATING
C446 a_7699_6397# VGND 0.609f $ **FLOATING
C447 a_7867_6299# VGND 0.817f $ **FLOATING
C448 a_7274_6397# VGND 0.626f $ **FLOATING
C449 a_7442_6143# VGND 0.581f $ **FLOATING
C450 a_7001_6031# VGND 1.43f $ **FLOATING
C451 a_6835_6031# VGND 1.81f $ **FLOATING
C452 a_3963_6397# VGND 0.168f $ **FLOATING
C453 a_3760_6031# VGND 0.259f $ **FLOATING
C454 tdc1.r_ring_ctr[12] VGND 10.5f $ **FLOATING
C455 tdc1.r_ring_ctr[14] VGND 2.56f $ **FLOATING
C456 _181_ VGND 5.09f $ **FLOATING
C457 a_5507_6005# VGND 0.729f $ **FLOATING
C458 a_4420_6031# VGND 0.736f $ **FLOATING
C459 a_4595_6005# VGND 0.971f $ **FLOATING
C460 a_3855_6031# VGND 0.714f $ **FLOATING
C461 _062_ VGND 1.6f $ **FLOATING
C462 a_4073_6273# VGND 0.653f $ **FLOATING
C463 a_3505_6031# VGND 1.57f $ **FLOATING
C464 _021_ VGND 1.08f $ **FLOATING
C465 a_3339_6031# VGND 1.92f $ **FLOATING
C466 a_28897_6575# VGND 0.214f $ **FLOATING
C467 a_28813_6575# VGND 0.167f $ **FLOATING
C468 a_27613_6575# VGND 0.23f $ **FLOATING
C469 tdc1.w_ring_int_norsz[13] VGND 3.87f $ **FLOATING
C470 a_20617_6575# VGND 0.214f $ **FLOATING
C471 a_20533_6575# VGND 0.167f $ **FLOATING
C472 a_24393_6575# VGND 0.23f $ **FLOATING
C473 a_21743_6895# VGND 0.319f $ **FLOATING
C474 tdc1.w_ring_buf[4] VGND 1.02f $ **FLOATING
C475 a_18781_6575# VGND 0.23f $ **FLOATING
C476 a_28731_6575# VGND 0.972f $ **FLOATING
C477 tdc1.r_dly_store_ring[28] VGND 1.2f $ **FLOATING
C478 tdc1.r_dly_store_ring[12] VGND 0.668f $ **FLOATING
C479 _106_ VGND 1.64f $ **FLOATING
C480 a_28123_6575# VGND 0.609f $ **FLOATING
C481 a_28291_6549# VGND 0.817f $ **FLOATING
C482 a_27698_6575# VGND 0.626f $ **FLOATING
C483 a_27866_6549# VGND 0.581f $ **FLOATING
C484 a_27425_6581# VGND 1.43f $ **FLOATING
C485 tdc1.w_ring_buf[12] VGND 1.14f $ **FLOATING
C486 a_27259_6581# VGND 1.81f $ **FLOATING
C487 tdc1.w_ring_int_norsz[12] VGND 0.722f $ **FLOATING
C488 tdc1.w_ring_norsz[28] VGND 2.59f $ **FLOATING
C489 tdc1.w_ring_norsz[12] VGND 2.32f $ **FLOATING
C490 a_24903_6575# VGND 0.609f $ **FLOATING
C491 a_25071_6549# VGND 0.817f $ **FLOATING
C492 a_24478_6575# VGND 0.626f $ **FLOATING
C493 a_24646_6549# VGND 0.581f $ **FLOATING
C494 a_24205_6581# VGND 1.43f $ **FLOATING
C495 tdc1.w_ring_buf[19] VGND 1.08f $ **FLOATING
C496 a_24039_6581# VGND 1.81f $ **FLOATING
C497 tdc1.w_ring_int_norsz[20] VGND 0.878f $ **FLOATING
C498 tdc1.w_ring_int_norsz[4] VGND 0.867f $ **FLOATING
C499 tdc1.w_ring_norsz[20] VGND 1.85f $ **FLOATING
C500 a_21912_6575# VGND 1.33f $ **FLOATING
C501 _108_ VGND 1.1f $ **FLOATING
C502 _107_ VGND 4.44f $ **FLOATING
C503 a_20451_6575# VGND 0.972f $ **FLOATING
C504 tdc1.r_dly_store_ring[4] VGND 1.1f $ **FLOATING
C505 tdc1.r_dly_store_ctr[12] VGND 1.1f $ **FLOATING
C506 a_20083_6575# VGND 0.524f $ **FLOATING
C507 a_19291_6575# VGND 0.609f $ **FLOATING
C508 a_19459_6549# VGND 0.817f $ **FLOATING
C509 a_18866_6575# VGND 0.626f $ **FLOATING
C510 a_19034_6549# VGND 0.581f $ **FLOATING
C511 a_18593_6581# VGND 1.43f $ **FLOATING
C512 tdc1.w_ring_buf[14] VGND 0.906f $ **FLOATING
C513 a_18427_6581# VGND 1.81f $ **FLOATING
C514 a_18151_6575# VGND 0.524f $ **FLOATING
C515 tdc1.w_ring_int_norsz[21] VGND 3.17f $ **FLOATING
C516 tdc1.g_ring3[30].stg01_75.HI VGND 0.415f $ **FLOATING
C517 net75 VGND 1.37f $ **FLOATING
C518 a_13629_6575# VGND 0.23f $ **FLOATING
C519 net14 VGND 4.11f $ **FLOATING
C520 a_14800_6549# VGND 0.648f $ **FLOATING
C521 a_14139_6575# VGND 0.609f $ **FLOATING
C522 a_14307_6549# VGND 0.817f $ **FLOATING
C523 a_13714_6575# VGND 0.626f $ **FLOATING
C524 a_13882_6549# VGND 0.581f $ **FLOATING
C525 a_13441_6581# VGND 1.43f $ **FLOATING
C526 tdc1.w_ring_buf[13] VGND 0.961f $ **FLOATING
C527 a_13275_6581# VGND 1.81f $ **FLOATING
C528 tdc1.w_ring_int_norsz[14] VGND 0.923f $ **FLOATING
C529 a_12539_6575# VGND 0.524f $ **FLOATING
C530 a_11713_6691# VGND 0.665f $ **FLOATING
C531 _126_ VGND 1.04f $ **FLOATING
C532 _127_ VGND 1.58f $ **FLOATING
C533 tdc1.w_ring_buf[22] VGND 1.06f $ **FLOATING
C534 a_11299_6794# VGND 0.524f $ **FLOATING
C535 tdc1.w_ring_norsz[30] VGND 5.09f $ **FLOATING
C536 net76 VGND 1f $ **FLOATING
C537 tdc1.w_ring_norsz[14] VGND 3.13f $ **FLOATING
C538 tdc1.g_ring3[31].stg01_76.HI VGND 0.415f $ **FLOATING
C539 a_6177_6575# VGND 0.23f $ **FLOATING
C540 tdc1.w_ring_int_norsz[31] VGND 0.956f $ **FLOATING
C541 tdc1.w_ring_int_norsz[15] VGND 0.984f $ **FLOATING
C542 a_6687_6575# VGND 0.609f $ **FLOATING
C543 a_6855_6549# VGND 0.817f $ **FLOATING
C544 a_6262_6575# VGND 0.626f $ **FLOATING
C545 a_6430_6549# VGND 0.581f $ **FLOATING
C546 a_5989_6581# VGND 1.43f $ **FLOATING
C547 tdc1.r_ring_ctr[13] VGND 3.66f $ **FLOATING
C548 a_5823_6581# VGND 1.81f $ **FLOATING
C549 a_29361_7119# VGND 0.23f $ **FLOATING
C550 a_29871_7485# VGND 0.609f $ **FLOATING
C551 a_30039_7387# VGND 0.817f $ **FLOATING
C552 a_29446_7485# VGND 0.626f $ **FLOATING
C553 a_29614_7231# VGND 0.581f $ **FLOATING
C554 a_29173_7119# VGND 1.43f $ **FLOATING
C555 a_29007_7119# VGND 1.81f $ **FLOATING
C556 tdc1.g_ring3[28].stg01_73.HI VGND 0.415f $ **FLOATING
C557 tdc1.w_ring_buf[27] VGND 1.11f $ **FLOATING
C558 a_28179_7119# VGND 0.524f $ **FLOATING
C559 a_27903_7119# VGND 0.524f $ **FLOATING
C560 tdc1.w_dly_stop[5] VGND 7.37f $ **FLOATING
C561 a_27411_7093# VGND 1.2f $ **FLOATING
C562 a_26615_7119# VGND 0.698f $ **FLOATING
C563 tdc1.w_ring_int_norsz[28] VGND 0.936f $ **FLOATING
C564 a_25125_7369# VGND 0.214f $ **FLOATING
C565 a_25041_7369# VGND 0.167f $ **FLOATING
C566 tdc1.g_ring3[22].stg01_67.HI VGND 0.415f $ **FLOATING
C567 a_21445_7369# VGND 0.214f $ **FLOATING
C568 a_21361_7369# VGND 0.167f $ **FLOATING
C569 tdc1.w_ring_int_norsz[5] VGND 1.17f $ **FLOATING
C570 net73 VGND 0.931f $ **FLOATING
C571 a_24959_7119# VGND 0.972f $ **FLOATING
C572 tdc1.r_dly_store_ring[19] VGND 0.815f $ **FLOATING
C573 tdc1.r_dly_store_ctr[3] VGND 1.69f $ **FLOATING
C574 a_24223_7119# VGND 0.524f $ **FLOATING
C575 tdc1.w_ring_norsz[3] VGND 2.68f $ **FLOATING
C576 tdc1.w_ring_norsz[19] VGND 2.26f $ **FLOATING
C577 a_21279_7119# VGND 0.972f $ **FLOATING
C578 tdc1.r_dly_store_ctr[2] VGND 1.54f $ **FLOATING
C579 tdc1.w_ring_norsz[4] VGND 3.84f $ **FLOATING
C580 net67 VGND 1.58f $ **FLOATING
C581 a_15193_7119# VGND 0.23f $ **FLOATING
C582 tdc1.w_ring_norsz[21] VGND 2.01f $ **FLOATING
C583 a_17555_7284# VGND 0.524f $ **FLOATING
C584 tdc1.w_ring_int_norsz[22] VGND 0.897f $ **FLOATING
C585 tdc1.w_ring_int_norsz[6] VGND 0.995f $ **FLOATING
C586 a_15703_7485# VGND 0.609f $ **FLOATING
C587 a_15871_7387# VGND 0.817f $ **FLOATING
C588 a_15278_7485# VGND 0.626f $ **FLOATING
C589 a_15446_7231# VGND 0.581f $ **FLOATING
C590 a_15005_7119# VGND 1.43f $ **FLOATING
C591 tdc1.w_ring_buf[21] VGND 1.77f $ **FLOATING
C592 a_14839_7119# VGND 1.81f $ **FLOATING
C593 a_13717_7369# VGND 0.214f $ **FLOATING
C594 a_13633_7369# VGND 0.167f $ **FLOATING
C595 a_13551_7119# VGND 0.972f $ **FLOATING
C596 tdc1.r_dly_store_ctr[5] VGND 1.79f $ **FLOATING
C597 tdc1.r_dly_store_ctr[13] VGND 4.44f $ **FLOATING
C598 tdc1.w_ring_norsz[22] VGND 4.85f $ **FLOATING
C599 net68 VGND 0.822f $ **FLOATING
C600 tdc1.g_ring3[23].stg01_68.HI VGND 0.415f $ **FLOATING
C601 a_10787_7369# VGND 0.253f $ **FLOATING
C602 a_9953_7369# VGND 0.206f $ **FLOATING
C603 a_8753_7119# VGND 0.23f $ **FLOATING
C604 tdc1.r_dly_store_ring[31] VGND 1.07f $ **FLOATING
C605 a_10569_7093# VGND 0.55f $ **FLOATING
C606 a_9871_7369# VGND 0.804f $ **FLOATING
C607 tdc1.r_dly_store_ctr[7] VGND 1.53f $ **FLOATING
C608 a_9263_7485# VGND 0.609f $ **FLOATING
C609 a_9431_7387# VGND 0.817f $ **FLOATING
C610 a_8838_7485# VGND 0.626f $ **FLOATING
C611 a_9006_7231# VGND 0.581f $ **FLOATING
C612 a_8565_7119# VGND 1.43f $ **FLOATING
C613 a_8399_7119# VGND 1.81f $ **FLOATING
C614 tdc1.w_ring_buf[31] VGND 1.42f $ **FLOATING
C615 tdc1.r_dly_store_ctr[15] VGND 2.31f $ **FLOATING
C616 a_5441_7119# VGND 0.23f $ **FLOATING
C617 tdc1.w_ring_norsz[15] VGND 1.73f $ **FLOATING
C618 a_7897_7284# VGND 0.524f $ **FLOATING
C619 a_7571_7119# VGND 0.524f $ **FLOATING
C620 a_7295_7119# VGND 0.524f $ **FLOATING
C621 tdc1.w_ring_norsz[31] VGND 2.54f $ **FLOATING
C622 a_5951_7485# VGND 0.609f $ **FLOATING
C623 a_6119_7387# VGND 0.817f $ **FLOATING
C624 a_5526_7485# VGND 0.626f $ **FLOATING
C625 a_5694_7231# VGND 0.581f $ **FLOATING
C626 a_5253_7119# VGND 1.43f $ **FLOATING
C627 a_5087_7119# VGND 1.81f $ **FLOATING
C628 a_3871_7485# VGND 0.168f $ **FLOATING
C629 a_3668_7119# VGND 0.259f $ **FLOATING
C630 a_4328_7119# VGND 0.736f $ **FLOATING
C631 a_4503_7093# VGND 0.971f $ **FLOATING
C632 a_3763_7119# VGND 0.714f $ **FLOATING
C633 _063_ VGND 1.61f $ **FLOATING
C634 a_3981_7361# VGND 0.653f $ **FLOATING
C635 a_3413_7119# VGND 1.57f $ **FLOATING
C636 a_3247_7119# VGND 1.92f $ **FLOATING
C637 _022_ VGND 1.11f $ **FLOATING
C638 a_2769_7369# VGND 0.219f $ **FLOATING
C639 a_2519_7369# VGND 0.684f $ **FLOATING
C640 tdc1.r_ring_ctr[15] VGND 2.28f $ **FLOATING
C641 _184_ VGND 3.24f $ **FLOATING
C642 a_29733_7663# VGND 0.206f $ **FLOATING
C643 a_30203_7663# VGND 0.227f $ **FLOATING
C644 a_28441_7663# VGND 0.23f $ **FLOATING
C645 a_24669_7663# VGND 0.23f $ **FLOATING
C646 tdc1.w_ring_int_norsz[19] VGND 1.01f $ **FLOATING
C647 tdc1.w_ring_int_norsz[3] VGND 0.962f $ **FLOATING
C648 a_30856_7895# VGND 0.535f $ **FLOATING
C649 a_30537_7895# VGND 0.5f $ **FLOATING
C650 a_30350_7637# VGND 0.578f $ **FLOATING
C651 a_30254_7895# VGND 0.498f $ **FLOATING
C652 tdc1.r_dly_store_ring[11] VGND 0.864f $ **FLOATING
C653 tdc1.r_dly_store_ring[27] VGND 1.1f $ **FLOATING
C654 a_29587_7895# VGND 0.804f $ **FLOATING
C655 a_28951_7663# VGND 0.609f $ **FLOATING
C656 a_29119_7637# VGND 0.817f $ **FLOATING
C657 a_28526_7663# VGND 0.626f $ **FLOATING
C658 a_28694_7637# VGND 0.581f $ **FLOATING
C659 a_28253_7669# VGND 1.43f $ **FLOATING
C660 tdc1.w_ring_buf[11] VGND 1.08f $ **FLOATING
C661 a_28087_7669# VGND 1.81f $ **FLOATING
C662 tdc1.w_ring_norsz[11] VGND 2.58f $ **FLOATING
C663 tdc1.w_ring_norsz[27] VGND 3f $ **FLOATING
C664 net19 VGND 12.5f $ **FLOATING
C665 a_27036_7637# VGND 0.648f $ **FLOATING
C666 a_25179_7663# VGND 0.609f $ **FLOATING
C667 a_25347_7637# VGND 0.817f $ **FLOATING
C668 a_24754_7663# VGND 0.626f $ **FLOATING
C669 a_24922_7637# VGND 0.581f $ **FLOATING
C670 a_24481_7669# VGND 1.43f $ **FLOATING
C671 tdc1.w_ring_buf[3] VGND 1.03f $ **FLOATING
C672 a_24315_7669# VGND 1.81f $ **FLOATING
C673 net64 VGND 1.05f $ **FLOATING
C674 tdc1.g_ring3[19].stg01_64.HI VGND 0.415f $ **FLOATING
C675 a_22261_8041# VGND 0.23f $ **FLOATING
C676 tdc1.r_dly_store_ring[18] VGND 0.997f $ **FLOATING
C677 _094_ VGND 1.08f $ **FLOATING
C678 a_23259_7882# VGND 0.524f $ **FLOATING
C679 tdc1.w_ring_buf[18] VGND 1.1f $ **FLOATING
C680 a_21843_8041# VGND 0.581f $ **FLOATING
C681 a_21914_7940# VGND 0.626f $ **FLOATING
C682 a_21714_7785# VGND 1.43f $ **FLOATING
C683 a_21707_7881# VGND 1.81f $ **FLOATING
C684 a_21423_7895# VGND 0.609f $ **FLOATING
C685 a_21327_7895# VGND 0.817f $ **FLOATING
C686 a_20157_7663# VGND 0.673f $ **FLOATING
C687 tdc1.r_dly_store_ctr[10] VGND 1.98f $ **FLOATING
C688 a_19991_7663# VGND 0.641f $ **FLOATING
C689 a_19535_7637# VGND 0.74f $ **FLOATING
C690 a_19425_7895# VGND 0.768f $ **FLOATING
C691 tdc1.r_dly_store_ring[14] VGND 1.42f $ **FLOATING
C692 _099_ VGND 3.44f $ **FLOATING
C693 a_16301_7663# VGND 0.206f $ **FLOATING
C694 a_13839_7663# VGND 0.167f $ **FLOATING
C695 a_13637_7663# VGND 0.214f $ **FLOATING
C696 tdc1.r_dly_store_ring[13] VGND 1.75f $ **FLOATING
C697 a_19066_7895# VGND 0.711f $ **FLOATING
C698 a_18501_7663# VGND 0.673f $ **FLOATING
C699 tdc1.r_dly_store_ctr[11] VGND 1.85f $ **FLOATING
C700 a_18335_7663# VGND 0.641f $ **FLOATING
C701 tdc1.w_ring_norsz[6] VGND 2.59f $ **FLOATING
C702 a_17739_7882# VGND 0.524f $ **FLOATING
C703 a_17375_7637# VGND 0.698f $ **FLOATING
C704 a_16771_7663# VGND 1.2f $ **FLOATING
C705 tdc1.r_dly_store_ring[21] VGND 1.08f $ **FLOATING
C706 tdc1.r_dly_store_ring[29] VGND 1.38f $ **FLOATING
C707 a_16155_7895# VGND 0.804f $ **FLOATING
C708 a_15543_7895# VGND 0.56f $ **FLOATING
C709 a_15025_7779# VGND 0.665f $ **FLOATING
C710 _118_ VGND 0.77f $ **FLOATING
C711 _119_ VGND 1.07f $ **FLOATING
C712 _120_ VGND 1.18f $ **FLOATING
C713 a_9677_7663# VGND 0.206f $ **FLOATING
C714 a_12341_7663# VGND 0.23f $ **FLOATING
C715 tdc1.r_dly_store_ctr[8] VGND 1.97f $ **FLOATING
C716 tdc1.r_dly_store_ring[8] VGND 0.749f $ **FLOATING
C717 a_13511_7895# VGND 0.972f $ **FLOATING
C718 a_12851_7663# VGND 0.609f $ **FLOATING
C719 a_13019_7637# VGND 0.817f $ **FLOATING
C720 a_12426_7663# VGND 0.626f $ **FLOATING
C721 a_12594_7637# VGND 0.581f $ **FLOATING
C722 a_12153_7669# VGND 1.43f $ **FLOATING
C723 a_11987_7669# VGND 1.81f $ **FLOATING
C724 tdc1.w_ring_int_norsz[7] VGND 3.12f $ **FLOATING
C725 tdc1.w_ring_int_norsz[23] VGND 1.04f $ **FLOATING
C726 a_10241_7779# VGND 0.665f $ **FLOATING
C727 _131_ VGND 0.922f $ **FLOATING
C728 _132_ VGND 0.856f $ **FLOATING
C729 _133_ VGND 0.654f $ **FLOATING
C730 a_6997_7663# VGND 0.329f $ **FLOATING
C731 a_6743_7663# VGND 0.381f $ **FLOATING
C732 a_8017_7663# VGND 0.23f $ **FLOATING
C733 a_9595_7663# VGND 0.804f $ **FLOATING
C734 tdc1.r_dly_store_ring[15] VGND 0.825f $ **FLOATING
C735 a_8527_7663# VGND 0.609f $ **FLOATING
C736 a_8695_7637# VGND 0.817f $ **FLOATING
C737 a_8102_7663# VGND 0.626f $ **FLOATING
C738 a_8270_7637# VGND 0.581f $ **FLOATING
C739 a_7829_7669# VGND 1.43f $ **FLOATING
C740 tdc1.w_ring_buf[15] VGND 1.03f $ **FLOATING
C741 a_7663_7669# VGND 1.81f $ **FLOATING
C742 tdc1.w_ring_int_norsz[0] VGND 1.04f $ **FLOATING
C743 tdc1.g_ring1[16].stg02_60.HI VGND 0.415f $ **FLOATING
C744 tdc1.g_ring3[16].stg01_61.HI VGND 0.415f $ **FLOATING
C745 net77 VGND 1.5f $ **FLOATING
C746 tdc1.stg01_77.HI VGND 0.415f $ **FLOATING
C747 _623_.X VGND 0.226f $ **FLOATING
C748 net61 VGND 1.06f $ **FLOATING
C749 net13 VGND 2.76f $ **FLOATING
C750 a_4588_7637# VGND 0.648f $ **FLOATING
C751 tdc1.g_ring3[27].stg01_72.HI VGND 0.415f $ **FLOATING
C752 a_29361_8207# VGND 0.23f $ **FLOATING
C753 a_29871_8573# VGND 0.609f $ **FLOATING
C754 a_30039_8475# VGND 0.817f $ **FLOATING
C755 a_29446_8573# VGND 0.626f $ **FLOATING
C756 a_29614_8319# VGND 0.581f $ **FLOATING
C757 a_29173_8207# VGND 1.43f $ **FLOATING
C758 a_29007_8207# VGND 1.81f $ **FLOATING
C759 tdc1.w_ring_buf[25] VGND 1.07f $ **FLOATING
C760 a_28271_8207# VGND 0.524f $ **FLOATING
C761 a_27351_8207# VGND 0.648f $ **FLOATING
C762 a_26983_8207# VGND 0.648f $ **FLOATING
C763 tdc1.w_ring_int_norsz[11] VGND 1.09f $ **FLOATING
C764 tdc1.w_ring_int_norsz[27] VGND 1.66f $ **FLOATING
C765 a_25609_8457# VGND 0.191f $ **FLOATING
C766 a_18877_8457# VGND 0.234f $ **FLOATING
C767 _129_ VGND 4.43f $ **FLOATING
C768 a_17493_8207# VGND 0.23f $ **FLOATING
C769 net72 VGND 1.4f $ **FLOATING
C770 _101_ VGND 2.29f $ **FLOATING
C771 _100_ VGND 1.09f $ **FLOATING
C772 tdc1.r_dly_store_ring[3] VGND 0.786f $ **FLOATING
C773 a_25472_8181# VGND 0.847f $ **FLOATING
C774 tdc1.w_ring_int_norsz[18] VGND 0.722f $ **FLOATING
C775 tdc1.w_ring_norsz[18] VGND 2.32f $ **FLOATING
C776 tdc1.w_ring_int_norsz[2] VGND 0.936f $ **FLOATING
C777 tdc1.w_ring_int_norsz[1] VGND 0.722f $ **FLOATING
C778 a_21003_8207# VGND 0.524f $ **FLOATING
C779 tdc1.w_ring_norsz[2] VGND 3.32f $ **FLOATING
C780 a_19655_8235# VGND 0.56f $ **FLOATING
C781 _128_ VGND 0.84f $ **FLOATING
C782 tdc1.r_dly_store_ring[6] VGND 1.08f $ **FLOATING
C783 a_18751_8359# VGND 0.953f $ **FLOATING
C784 a_18003_8573# VGND 0.609f $ **FLOATING
C785 a_18171_8475# VGND 0.817f $ **FLOATING
C786 a_17578_8573# VGND 0.626f $ **FLOATING
C787 a_17746_8319# VGND 0.581f $ **FLOATING
C788 a_17305_8207# VGND 1.43f $ **FLOATING
C789 tdc1.w_ring_buf[6] VGND 1.03f $ **FLOATING
C790 a_17139_8207# VGND 1.81f $ **FLOATING
C791 a_16587_8207# VGND 0.648f $ **FLOATING
C792 a_15701_8457# VGND 0.422f $ **FLOATING
C793 a_15283_8457# VGND 0.495f $ **FLOATING
C794 tdc1.r_dly_store_ctr[0] VGND 2.31f $ **FLOATING
C795 tdc1.g_ring3[24].stg01_69.HI VGND 0.415f $ **FLOATING
C796 tdc1.w_ring_buf[8] VGND 1.03f $ **FLOATING
C797 a_15335_8181# VGND 1.45f $ **FLOATING
C798 a_13887_8359# VGND 0.56f $ **FLOATING
C799 a_12587_8372# VGND 0.524f $ **FLOATING
C800 tdc1.w_ring_norsz[8] VGND 2.78f $ **FLOATING
C801 net16 VGND 9.22f $ **FLOATING
C802 tdc1.w_ring_int_norsz[8] VGND 0.839f $ **FLOATING
C803 tdc1.w_ring_int_norsz[24] VGND 1.1f $ **FLOATING
C804 tdc1.r_dly_store_ring[23] VGND 0.95f $ **FLOATING
C805 a_9213_8207# VGND 0.23f $ **FLOATING
C806 net69 VGND 0.97f $ **FLOATING
C807 a_9723_8573# VGND 0.609f $ **FLOATING
C808 a_9891_8475# VGND 0.817f $ **FLOATING
C809 a_9298_8573# VGND 0.626f $ **FLOATING
C810 a_9466_8319# VGND 0.581f $ **FLOATING
C811 a_9025_8207# VGND 1.43f $ **FLOATING
C812 a_8859_8207# VGND 1.81f $ **FLOATING
C813 a_6813_8457# VGND 0.329f $ **FLOATING
C814 a_6559_8457# VGND 0.381f $ **FLOATING
C815 a_6077_8457# VGND 0.329f $ **FLOATING
C816 a_5823_8457# VGND 0.381f $ **FLOATING
C817 tdc1.w_ring_buf[0] VGND 7f $ **FLOATING
C818 a_3601_8207# VGND 0.23f $ **FLOATING
C819 net60 VGND 1.42f $ **FLOATING
C820 net15 VGND 11.5f $ **FLOATING
C821 tdc1.w_ring_int_norsz[16] VGND 2.87f $ **FLOATING
C822 a_5547_8207# VGND 0.524f $ **FLOATING
C823 tdc1.w_ring_norsz[0] VGND 10.1f $ **FLOATING
C824 tdc1.w_ring_norsz[7] VGND 4.56f $ **FLOATING
C825 a_5043_8372# VGND 0.524f $ **FLOATING
C826 a_4111_8573# VGND 0.609f $ **FLOATING
C827 a_4279_8475# VGND 0.817f $ **FLOATING
C828 a_3686_8573# VGND 0.626f $ **FLOATING
C829 a_3854_8319# VGND 0.581f $ **FLOATING
C830 a_3413_8207# VGND 1.43f $ **FLOATING
C831 net7 VGND 15.7f $ **FLOATING
C832 a_3247_8207# VGND 1.81f $ **FLOATING
C833 a_30101_8751# VGND 0.206f $ **FLOATING
C834 a_28809_8751# VGND 0.23f $ **FLOATING
C835 tdc1.r_dly_store_ring[9] VGND 0.864f $ **FLOATING
C836 tdc1.r_dly_store_ring[25] VGND 0.918f $ **FLOATING
C837 a_29955_8983# VGND 0.804f $ **FLOATING
C838 a_29319_8751# VGND 0.609f $ **FLOATING
C839 a_29487_8725# VGND 0.817f $ **FLOATING
C840 a_28894_8751# VGND 0.626f $ **FLOATING
C841 a_29062_8725# VGND 0.581f $ **FLOATING
C842 a_28621_8757# VGND 1.43f $ **FLOATING
C843 a_28455_8757# VGND 1.81f $ **FLOATING
C844 tdc1.g_ring3[26].stg01_71.HI VGND 0.415f $ **FLOATING
C845 net71 VGND 1.09f $ **FLOATING
C846 a_25847_8751# VGND 0.245f $ **FLOATING
C847 net63 VGND 1.34f $ **FLOATING
C848 a_24485_8751# VGND 0.23f $ **FLOATING
C849 tdc1.w_ring_int_norsz[26] VGND 0.969f $ **FLOATING
C850 tdc1.w_ring_norsz[25] VGND 2.43f $ **FLOATING
C851 tdc1.w_ring_int_norsz[9] VGND 6.8f $ **FLOATING
C852 net18 VGND 4.34f $ **FLOATING
C853 tdc1.w_ring_int_norsz[25] VGND 7.31f $ **FLOATING
C854 tdc1.r_dly_store_ring[17] VGND 0.819f $ **FLOATING
C855 _073_ VGND 2.56f $ **FLOATING
C856 _078_ VGND 2.08f $ **FLOATING
C857 a_24995_8751# VGND 0.609f $ **FLOATING
C858 a_25163_8725# VGND 0.817f $ **FLOATING
C859 a_24570_8751# VGND 0.626f $ **FLOATING
C860 a_24738_8725# VGND 0.581f $ **FLOATING
C861 a_24297_8757# VGND 1.43f $ **FLOATING
C862 tdc1.w_ring_buf[17] VGND 0.872f $ **FLOATING
C863 a_24131_8757# VGND 1.81f $ **FLOATING
C864 a_23855_8751# VGND 0.524f $ **FLOATING
C865 tdc1.g_ring3[18].stg01_63.HI VGND 0.415f $ **FLOATING
C866 tdc1.w_ring_norsz[17] VGND 2.67f $ **FLOATING
C867 a_18690_8751# VGND 0.324f $ **FLOATING
C868 a_21633_8751# VGND 0.23f $ **FLOATING
C869 net17 VGND 8.21f $ **FLOATING
C870 tdc1.w_ring_int_norsz[17] VGND 7.72f $ **FLOATING
C871 a_22143_8751# VGND 0.609f $ **FLOATING
C872 a_22311_8725# VGND 0.817f $ **FLOATING
C873 a_21718_8751# VGND 0.626f $ **FLOATING
C874 a_21886_8725# VGND 0.581f $ **FLOATING
C875 a_21445_8757# VGND 1.43f $ **FLOATING
C876 tdc1.w_ring_buf[2] VGND 1.11f $ **FLOATING
C877 a_21279_8757# VGND 1.81f $ **FLOATING
C878 a_20083_8751# VGND 0.988f $ **FLOATING
C879 _082_ VGND 0.877f $ **FLOATING
C880 a_19631_8867# VGND 0.485f $ **FLOATING
C881 a_19439_9111# VGND 0.478f $ **FLOATING
C882 a_18776_9071# VGND 0.337f $ **FLOATING
C883 a_18243_9071# VGND 0.28f $ **FLOATING
C884 a_14909_8751# VGND 0.393f $ **FLOATING
C885 a_14655_8751# VGND 0.388f $ **FLOATING
C886 a_12897_8751# VGND 0.206f $ **FLOATING
C887 a_18243_8751# VGND 1.14f $ **FLOATING
C888 tdc1.w_ring_norsz[5] VGND 2.74f $ **FLOATING
C889 a_17739_8970# VGND 0.524f $ **FLOATING
C890 a_17323_8759# VGND 0.648f $ **FLOATING
C891 a_16771_8751# VGND 1.2f $ **FLOATING
C892 a_16309_8867# VGND 0.601f $ **FLOATING
C893 net5 VGND 4.77f $ **FLOATING
C894 net4 VGND 4.51f $ **FLOATING
C895 a_16209_8751# VGND 0.488f $ **FLOATING
C896 a_15159_8725# VGND 0.587f $ **FLOATING
C897 a_14332_8983# VGND 0.488f $ **FLOATING
C898 net70 VGND 1.22f $ **FLOATING
C899 a_14059_8983# VGND 0.601f $ **FLOATING
C900 a_13553_8867# VGND 0.665f $ **FLOATING
C901 _186_ VGND 0.96f $ **FLOATING
C902 _188_ VGND 1.08f $ **FLOATING
C903 _187_ VGND 0.753f $ **FLOATING
C904 a_12815_8751# VGND 0.804f $ **FLOATING
C905 tdc1.w_ring_norsz[24] VGND 2.44f $ **FLOATING
C906 a_12403_8970# VGND 0.524f $ **FLOATING
C907 tdc1.g_ring3[25].stg01_70.HI VGND 0.415f $ **FLOATING
C908 tdc1.w_ring_buf[23] VGND 1.09f $ **FLOATING
C909 tdc1.r_dly_store_ring[16] VGND 2.56f $ **FLOATING
C910 net62 VGND 1.18f $ **FLOATING
C911 a_7649_8751# VGND 0.23f $ **FLOATING
C912 a_11763_8725# VGND 0.698f $ **FLOATING
C913 a_10975_8751# VGND 1.2f $ **FLOATING
C914 a_9963_8751# VGND 1.2f $ **FLOATING
C915 tdc1.w_ring_norsz[23] VGND 2.96f $ **FLOATING
C916 a_9459_8970# VGND 0.524f $ **FLOATING
C917 a_8159_8751# VGND 0.609f $ **FLOATING
C918 a_8327_8725# VGND 0.817f $ **FLOATING
C919 a_7734_8751# VGND 0.626f $ **FLOATING
C920 a_7902_8725# VGND 0.581f $ **FLOATING
C921 a_7461_8757# VGND 1.43f $ **FLOATING
C922 a_7295_8757# VGND 1.81f $ **FLOATING
C923 tdc1.g_ring3[17].stg01_62.HI VGND 0.415f $ **FLOATING
C924 a_4613_8751# VGND 0.23f $ **FLOATING
C925 _620_.X VGND 0.226f $ **FLOATING
C926 _621_.X VGND 0.226f $ **FLOATING
C927 a_6743_8751# VGND 0.524f $ **FLOATING
C928 a_5123_8751# VGND 0.609f $ **FLOATING
C929 a_5291_8725# VGND 0.817f $ **FLOATING
C930 a_4698_8751# VGND 0.626f $ **FLOATING
C931 a_4866_8725# VGND 0.581f $ **FLOATING
C932 a_4425_8757# VGND 1.43f $ **FLOATING
C933 tdc1.w_ring_buf[7] VGND 1.16f $ **FLOATING
C934 a_4259_8757# VGND 1.81f $ **FLOATING
C935 a_3392_8725# VGND 0.648f $ **FLOATING
C936 a_3024_8725# VGND 0.648f $ **FLOATING
C937 a_29181_9545# VGND 0.206f $ **FLOATING
C938 tdc1.w_ring_buf[9] VGND 1.17f $ **FLOATING
C939 tdc1.w_ring_int_norsz[10] VGND 1.15f $ **FLOATING
C940 _095_ VGND 3.29f $ **FLOATING
C941 _096_ VGND 1.92f $ **FLOATING
C942 a_24591_9545# VGND 0.238f $ **FLOATING
C943 a_29035_9447# VGND 0.804f $ **FLOATING
C944 a_27903_9295# VGND 0.524f $ **FLOATING
C945 a_27443_9295# VGND 0.524f $ **FLOATING
C946 tdc1.w_ring_norsz[26] VGND 2.58f $ **FLOATING
C947 tdc1.w_ring_norsz[9] VGND 2.54f $ **FLOATING
C948 tdc1.w_ring_norsz[10] VGND 2.51f $ **FLOATING
C949 a_26847_9460# VGND 0.524f $ **FLOATING
C950 a_25973_9301# VGND 0.665f $ **FLOATING
C951 net34 VGND 11.4f $ **FLOATING
C952 _097_ VGND 2.21f $ **FLOATING
C953 a_22351_9545# VGND 0.203f $ **FLOATING
C954 a_21637_9545# VGND 0.234f $ **FLOATING
C955 a_15772_9295# VGND 0.123f $ **FLOATING
C956 a_15420_9295# VGND 0.161f $ **FLOATING
C957 a_14442_9295# VGND 0.161f $ **FLOATING
C958 a_14090_9295# VGND 0.123f $ **FLOATING
C959 a_17033_9295# VGND 0.23f $ **FLOATING
C960 a_24276_9269# VGND 0.648f $ **FLOATING
C961 a_23119_9295# VGND 0.524f $ **FLOATING
C962 tdc1.w_ring_norsz[1] VGND 2.36f $ **FLOATING
C963 a_22257_9545# VGND 0.655f $ **FLOATING
C964 tdc1.r_dly_store_ring[2] VGND 0.911f $ **FLOATING
C965 _111_ VGND 1.33f $ **FLOATING
C966 _080_ VGND 4.04f $ **FLOATING
C967 _081_ VGND 4.42f $ **FLOATING
C968 a_21511_9447# VGND 0.953f $ **FLOATING
C969 a_20065_9661# VGND 0.673f $ **FLOATING
C970 a_19899_9295# VGND 0.641f $ **FLOATING
C971 a_17543_9661# VGND 0.609f $ **FLOATING
C972 a_17711_9563# VGND 0.817f $ **FLOATING
C973 a_17118_9661# VGND 0.626f $ **FLOATING
C974 a_17286_9407# VGND 0.581f $ **FLOATING
C975 a_16845_9295# VGND 1.43f $ **FLOATING
C976 tdc1.w_ring_buf[5] VGND 1.23f $ **FLOATING
C977 a_16679_9295# VGND 1.81f $ **FLOATING
C978 net31 VGND 12.8f $ **FLOATING
C979 a_15333_9545# VGND 0.537f $ **FLOATING
C980 a_14008_9545# VGND 0.537f $ **FLOATING
C981 tdc1.r_dly_store_ring[24] VGND 0.826f $ **FLOATING
C982 a_10946_9295# VGND 0.161f $ **FLOATING
C983 a_10594_9295# VGND 0.123f $ **FLOATING
C984 a_11973_9295# VGND 0.23f $ **FLOATING
C985 a_15504_9295# VGND 1.37f $ **FLOATING
C986 _121_ VGND 1.54f $ **FLOATING
C987 _189_ VGND 1.16f $ **FLOATING
C988 a_13620_9269# VGND 1.37f $ **FLOATING
C989 a_12483_9661# VGND 0.609f $ **FLOATING
C990 a_12651_9563# VGND 0.817f $ **FLOATING
C991 a_12058_9661# VGND 0.626f $ **FLOATING
C992 a_12226_9407# VGND 0.581f $ **FLOATING
C993 a_11785_9295# VGND 1.43f $ **FLOATING
C994 tdc1.w_ring_buf[24] VGND 1.22f $ **FLOATING
C995 a_11619_9295# VGND 1.81f $ **FLOATING
C996 net30 VGND 11.7f $ **FLOATING
C997 a_10512_9545# VGND 0.537f $ **FLOATING
C998 tdc1.w_ring_buf[16] VGND 1.41f $ **FLOATING
C999 tdc1.r_dly_store_ring[7] VGND 1.21f $ **FLOATING
C1000 a_5773_9622# VGND 0.607f $ **FLOATING
C1001 _194_ VGND 4.49f $ **FLOATING
C1002 tdc1.r_dly_store_ring[0] VGND 1.43f $ **FLOATING
C1003 a_4761_9622# VGND 0.607f $ **FLOATING
C1004 tdc0.r_dly_store_ring[0] VGND 0.979f $ **FLOATING
C1005 a_3601_9295# VGND 0.23f $ **FLOATING
C1006 _134_ VGND 1.51f $ **FLOATING
C1007 _139_ VGND 2.53f $ **FLOATING
C1008 a_10124_9269# VGND 1.37f $ **FLOATING
C1009 a_9503_9295# VGND 1.2f $ **FLOATING
C1010 a_7111_9295# VGND 0.524f $ **FLOATING
C1011 tdc1.w_ring_norsz[16] VGND 3.9f $ **FLOATING
C1012 a_6027_9622# VGND 0.59f $ **FLOATING
C1013 a_5015_9622# VGND 0.59f $ **FLOATING
C1014 a_4111_9661# VGND 0.609f $ **FLOATING
C1015 a_4279_9563# VGND 0.817f $ **FLOATING
C1016 a_3686_9661# VGND 0.626f $ **FLOATING
C1017 a_3854_9407# VGND 0.581f $ **FLOATING
C1018 a_3413_9295# VGND 1.43f $ **FLOATING
C1019 a_3247_9295# VGND 1.81f $ **FLOATING
C1020 tdc1.r_dly_store_ring[26] VGND 0.918f $ **FLOATING
C1021 a_28441_9839# VGND 0.23f $ **FLOATING
C1022 tdc1.r_dly_store_ring[10] VGND 1.47f $ **FLOATING
C1023 a_24765_9839# VGND 0.171f $ **FLOATING
C1024 a_26969_9839# VGND 0.23f $ **FLOATING
C1025 a_25373_10159# VGND 0.155f $ **FLOATING
C1026 a_24683_10159# VGND 0.398f $ **FLOATING
C1027 tdc1.r_dly_store_ring[1] VGND 0.964f $ **FLOATING
C1028 a_23473_9839# VGND 0.23f $ **FLOATING
C1029 tdc0.r_dly_store_ring[4] VGND 1.31f $ **FLOATING
C1030 a_21633_9839# VGND 0.23f $ **FLOATING
C1031 _113_ VGND 2.61f $ **FLOATING
C1032 a_28951_9839# VGND 0.609f $ **FLOATING
C1033 a_29119_9813# VGND 0.817f $ **FLOATING
C1034 a_28526_9839# VGND 0.626f $ **FLOATING
C1035 a_28694_9813# VGND 0.581f $ **FLOATING
C1036 a_28253_9845# VGND 1.43f $ **FLOATING
C1037 tdc1.w_ring_buf[26] VGND 1.28f $ **FLOATING
C1038 a_28087_9845# VGND 1.81f $ **FLOATING
C1039 a_27479_9839# VGND 0.609f $ **FLOATING
C1040 a_27647_9813# VGND 0.817f $ **FLOATING
C1041 a_27054_9839# VGND 0.626f $ **FLOATING
C1042 a_27222_9813# VGND 0.581f $ **FLOATING
C1043 a_26781_9845# VGND 1.43f $ **FLOATING
C1044 tdc1.w_ring_buf[10] VGND 1.01f $ **FLOATING
C1045 a_26615_9845# VGND 1.81f $ **FLOATING
C1046 a_24849_9839# VGND 1.43f $ **FLOATING
C1047 _085_ VGND 1.2f $ **FLOATING
C1048 _079_ VGND 1.55f $ **FLOATING
C1049 a_25071_9813# VGND 0.822f $ **FLOATING
C1050 a_23983_9839# VGND 0.609f $ **FLOATING
C1051 a_24151_9813# VGND 0.817f $ **FLOATING
C1052 a_23558_9839# VGND 0.626f $ **FLOATING
C1053 a_23726_9813# VGND 0.581f $ **FLOATING
C1054 a_23285_9845# VGND 1.43f $ **FLOATING
C1055 tdc1.w_ring_buf[1] VGND 1.01f $ **FLOATING
C1056 a_23119_9845# VGND 1.81f $ **FLOATING
C1057 a_22143_9839# VGND 0.609f $ **FLOATING
C1058 a_22311_9813# VGND 0.817f $ **FLOATING
C1059 a_21718_9839# VGND 0.626f $ **FLOATING
C1060 a_21886_9813# VGND 0.581f $ **FLOATING
C1061 a_21445_9845# VGND 1.43f $ **FLOATING
C1062 a_21279_9845# VGND 1.81f $ **FLOATING
C1063 a_20729_9955# VGND 0.665f $ **FLOATING
C1064 _112_ VGND 1.15f $ **FLOATING
C1065 _122_ VGND 1.73f $ **FLOATING
C1066 a_10229_9839# VGND 0.206f $ **FLOATING
C1067 a_9577_9839# VGND 0.214f $ **FLOATING
C1068 a_9493_9839# VGND 0.167f $ **FLOATING
C1069 a_16573_9839# VGND 0.23f $ **FLOATING
C1070 net6 VGND 5.69f $ **FLOATING
C1071 _138_ VGND 1.38f $ **FLOATING
C1072 a_19329_9839# VGND 0.673f $ **FLOATING
C1073 a_19163_9839# VGND 0.641f $ **FLOATING
C1074 _065_ VGND 10.8f $ **FLOATING
C1075 a_18169_10137# VGND 0.607f $ **FLOATING
C1076 tdc0.r_dly_store_ring[5] VGND 0.948f $ **FLOATING
C1077 tdc1.r_dly_store_ring[5] VGND 1.15f $ **FLOATING
C1078 a_17740_10071# VGND 0.59f $ **FLOATING
C1079 a_17083_9839# VGND 0.609f $ **FLOATING
C1080 a_17251_9813# VGND 0.817f $ **FLOATING
C1081 a_16658_9839# VGND 0.626f $ **FLOATING
C1082 a_16826_9813# VGND 0.581f $ **FLOATING
C1083 a_16385_9845# VGND 1.43f $ **FLOATING
C1084 a_16219_9845# VGND 1.81f $ **FLOATING
C1085 a_14794_9922# VGND 0.611f $ **FLOATING
C1086 _064_ VGND 9.76f $ **FLOATING
C1087 _070_ VGND 11.5f $ **FLOATING
C1088 a_14011_9839# VGND 1.2f $ **FLOATING
C1089 a_12539_9839# VGND 1.2f $ **FLOATING
C1090 a_11987_9839# VGND 1.2f $ **FLOATING
C1091 a_10977_9955# VGND 0.665f $ **FLOATING
C1092 _136_ VGND 0.792f $ **FLOATING
C1093 _137_ VGND 1.01f $ **FLOATING
C1094 a_8017_9839# VGND 0.23f $ **FLOATING
C1095 a_6545_9839# VGND 0.23f $ **FLOATING
C1096 tdc0.r_dly_store_ring[7] VGND 1.21f $ **FLOATING
C1097 a_4613_9839# VGND 0.23f $ **FLOATING
C1098 net26 VGND 10.5f $ **FLOATING
C1099 a_10147_9839# VGND 0.804f $ **FLOATING
C1100 tdc0.r_dly_store_ring[23] VGND 1.25f $ **FLOATING
C1101 _076_ VGND 5.59f $ **FLOATING
C1102 a_9411_9839# VGND 0.972f $ **FLOATING
C1103 tdc0.r_dly_store_ring[15] VGND 1.43f $ **FLOATING
C1104 a_8527_9839# VGND 0.609f $ **FLOATING
C1105 a_8695_9813# VGND 0.817f $ **FLOATING
C1106 a_8102_9839# VGND 0.626f $ **FLOATING
C1107 a_8270_9813# VGND 0.581f $ **FLOATING
C1108 a_7829_9845# VGND 1.43f $ **FLOATING
C1109 a_7663_9845# VGND 1.81f $ **FLOATING
C1110 a_7055_9839# VGND 0.609f $ **FLOATING
C1111 a_7223_9813# VGND 0.817f $ **FLOATING
C1112 a_6630_9839# VGND 0.626f $ **FLOATING
C1113 a_6798_9813# VGND 0.581f $ **FLOATING
C1114 a_6357_9845# VGND 1.43f $ **FLOATING
C1115 a_6191_9845# VGND 1.81f $ **FLOATING
C1116 a_5123_9839# VGND 0.609f $ **FLOATING
C1117 a_5291_9813# VGND 0.817f $ **FLOATING
C1118 a_4698_9839# VGND 0.626f $ **FLOATING
C1119 a_4866_9813# VGND 0.581f $ **FLOATING
C1120 a_4425_9845# VGND 1.43f $ **FLOATING
C1121 a_4259_9845# VGND 1.81f $ **FLOATING
C1122 a_3115_9813# VGND 0.698f $ **FLOATING
C1123 a_25182_10383# VGND 0.482f $ **FLOATING
C1124 a_25616_10633# VGND 0.14f $ **FLOATING
C1125 a_25264_10633# VGND 0.171f $ **FLOATING
C1126 a_25348_10633# VGND 1.37f $ **FLOATING
C1127 _102_ VGND 1.58f $ **FLOATING
C1128 _084_ VGND 13.5f $ **FLOATING
C1129 a_23273_10383# VGND 0.23f $ **FLOATING
C1130 a_21545_10633# VGND 0.206f $ **FLOATING
C1131 _109_ VGND 1.04f $ **FLOATING
C1132 tdc0.w_ring_buf[4] VGND 1.18f $ **FLOATING
C1133 tdc0.r_dly_store_ring[25] VGND 1.19f $ **FLOATING
C1134 a_19057_10383# VGND 0.23f $ **FLOATING
C1135 a_22855_10383# VGND 0.581f $ **FLOATING
C1136 a_22926_10357# VGND 0.626f $ **FLOATING
C1137 a_22719_10357# VGND 1.81f $ **FLOATING
C1138 a_22726_10657# VGND 1.43f $ **FLOATING
C1139 a_22435_10357# VGND 0.609f $ **FLOATING
C1140 a_22339_10535# VGND 0.817f $ **FLOATING
C1141 tdc0.r_dly_store_ring[20] VGND 0.877f $ **FLOATING
C1142 a_21399_10535# VGND 0.804f $ **FLOATING
C1143 a_20727_10383# VGND 0.524f $ **FLOATING
C1144 a_19567_10749# VGND 0.609f $ **FLOATING
C1145 a_19735_10651# VGND 0.817f $ **FLOATING
C1146 a_19142_10749# VGND 0.626f $ **FLOATING
C1147 a_19310_10495# VGND 0.581f $ **FLOATING
C1148 a_18869_10383# VGND 1.43f $ **FLOATING
C1149 a_18703_10383# VGND 1.81f $ **FLOATING
C1150 tdc0.w_ring_buf[5] VGND 0.977f $ **FLOATING
C1151 _117_ VGND 1.24f $ **FLOATING
C1152 _193_ VGND 1.4f $ **FLOATING
C1153 _192_ VGND 0.661f $ **FLOATING
C1154 a_13633_10633# VGND 0.206f $ **FLOATING
C1155 a_12065_10383# VGND 0.23f $ **FLOATING
C1156 a_16219_10383# VGND 0.524f $ **FLOATING
C1157 a_15719_10357# VGND 0.698f $ **FLOATING
C1158 a_15256_10535# VGND 0.665f $ **FLOATING
C1159 a_14197_10389# VGND 0.665f $ **FLOATING
C1160 a_13551_10633# VGND 0.804f $ **FLOATING
C1161 net25 VGND 7.77f $ **FLOATING
C1162 _071_ VGND 8.55f $ **FLOATING
C1163 tdc0.r_dly_store_ring[8] VGND 0.786f $ **FLOATING
C1164 a_12575_10749# VGND 0.609f $ **FLOATING
C1165 a_12743_10651# VGND 0.817f $ **FLOATING
C1166 a_12150_10749# VGND 0.626f $ **FLOATING
C1167 a_12318_10495# VGND 0.581f $ **FLOATING
C1168 a_11877_10383# VGND 1.43f $ **FLOATING
C1169 a_11711_10383# VGND 1.81f $ **FLOATING
C1170 tdc0.w_ring_buf[8] VGND 0.872f $ **FLOATING
C1171 _191_ VGND 1.92f $ **FLOATING
C1172 a_10781_10633# VGND 0.206f $ **FLOATING
C1173 _135_ VGND 1.28f $ **FLOATING
C1174 tdc0.w_ring_buf[23] VGND 0.949f $ **FLOATING
C1175 tdc0.r_dly_store_ring[31] VGND 1.99f $ **FLOATING
C1176 a_5993_10383# VGND 0.23f $ **FLOATING
C1177 a_11435_10383# VGND 0.524f $ **FLOATING
C1178 a_10699_10633# VGND 0.804f $ **FLOATING
C1179 _068_ VGND 6.13f $ **FLOATING
C1180 a_10087_10411# VGND 0.56f $ **FLOATING
C1181 a_7755_10383# VGND 0.524f $ **FLOATING
C1182 a_6503_10749# VGND 0.609f $ **FLOATING
C1183 a_6671_10651# VGND 0.817f $ **FLOATING
C1184 a_6078_10749# VGND 0.626f $ **FLOATING
C1185 a_6246_10495# VGND 0.581f $ **FLOATING
C1186 a_5805_10383# VGND 1.43f $ **FLOATING
C1187 a_5639_10383# VGND 1.81f $ **FLOATING
C1188 tdc0.w_ring_buf[7] VGND 1.12f $ **FLOATING
C1189 tdc0.r_dly_store_ctr[15] VGND 3.17f $ **FLOATING
C1190 a_3785_10383# VGND 0.23f $ **FLOATING
C1191 a_5043_10548# VGND 0.524f $ **FLOATING
C1192 a_4295_10749# VGND 0.609f $ **FLOATING
C1193 a_4463_10651# VGND 0.817f $ **FLOATING
C1194 a_3870_10749# VGND 0.626f $ **FLOATING
C1195 a_4038_10495# VGND 0.581f $ **FLOATING
C1196 a_3597_10383# VGND 1.43f $ **FLOATING
C1197 a_3431_10383# VGND 1.81f $ **FLOATING
C1198 net3 VGND 5.88f $ **FLOATING
C1199 a_855_10383# VGND 0.524f $ **FLOATING
C1200 a_27413_11305# VGND 0.23f $ **FLOATING
C1201 a_25677_10927# VGND 0.214f $ **FLOATING
C1202 a_25593_10927# VGND 0.167f $ **FLOATING
C1203 _105_ VGND 1.12f $ **FLOATING
C1204 a_24393_10927# VGND 0.23f $ **FLOATING
C1205 tdc0.w_ring_buf[20] VGND 1.13f $ **FLOATING
C1206 tdc0.r_dly_store_ring[28] VGND 1.64f $ **FLOATING
C1207 a_18781_10927# VGND 0.23f $ **FLOATING
C1208 tdc0.w_ring_buf[25] VGND 1.35f $ **FLOATING
C1209 a_26995_11305# VGND 0.581f $ **FLOATING
C1210 a_27066_11204# VGND 0.626f $ **FLOATING
C1211 a_26866_11049# VGND 1.43f $ **FLOATING
C1212 a_26859_11145# VGND 1.81f $ **FLOATING
C1213 a_26575_11159# VGND 0.609f $ **FLOATING
C1214 a_26479_11159# VGND 0.817f $ **FLOATING
C1215 a_25511_10927# VGND 0.972f $ **FLOATING
C1216 tdc0.r_dly_store_ring[27] VGND 0.827f $ **FLOATING
C1217 tdc0.r_dly_store_ring[3] VGND 0.668f $ **FLOATING
C1218 a_24903_10927# VGND 0.609f $ **FLOATING
C1219 a_25071_10901# VGND 0.817f $ **FLOATING
C1220 a_24478_10927# VGND 0.626f $ **FLOATING
C1221 a_24646_10901# VGND 0.581f $ **FLOATING
C1222 a_24205_10933# VGND 1.43f $ **FLOATING
C1223 tdc0.w_ring_buf[3] VGND 0.872f $ **FLOATING
C1224 a_24039_10933# VGND 1.81f $ **FLOATING
C1225 a_23763_10927# VGND 0.524f $ **FLOATING
C1226 a_22843_10927# VGND 0.524f $ **FLOATING
C1227 tdc0.w_ring_int_norsz[4] VGND 1.11f $ **FLOATING
C1228 a_19899_10927# VGND 0.524f $ **FLOATING
C1229 a_19291_10927# VGND 0.609f $ **FLOATING
C1230 a_19459_10901# VGND 0.817f $ **FLOATING
C1231 a_18866_10927# VGND 0.626f $ **FLOATING
C1232 a_19034_10901# VGND 0.581f $ **FLOATING
C1233 a_18593_10933# VGND 1.43f $ **FLOATING
C1234 tdc0.w_ring_buf[28] VGND 0.872f $ **FLOATING
C1235 a_18427_10933# VGND 1.81f $ **FLOATING
C1236 a_18151_10927# VGND 0.524f $ **FLOATING
C1237 a_17875_10927# VGND 0.524f $ **FLOATING
C1238 tdc0.g_ring3[21].stg01_48.HI VGND 0.415f $ **FLOATING
C1239 a_15289_10927# VGND 0.206f $ **FLOATING
C1240 _115_ VGND 0.941f $ **FLOATING
C1241 a_14089_10927# VGND 0.23f $ **FLOATING
C1242 tdc0.r_dly_store_ring[24] VGND 0.918f $ **FLOATING
C1243 a_9765_10927# VGND 0.23f $ **FLOATING
C1244 a_3108_10927# VGND 0.168f $ **FLOATING
C1245 tdc0.w_ring_buf[31] VGND 1.02f $ **FLOATING
C1246 a_3526_10927# VGND 0.259f $ **FLOATING
C1247 tdc0.w_ring_norsz[4] VGND 4.16f $ **FLOATING
C1248 tdc0.w_ring_norsz[20] VGND 4.79f $ **FLOATING
C1249 net48 VGND 1.23f $ **FLOATING
C1250 tdc0.w_ring_int_norsz[21] VGND 0.722f $ **FLOATING
C1251 tdc0.w_ring_int_norsz[5] VGND 1.17f $ **FLOATING
C1252 a_15207_10927# VGND 0.804f $ **FLOATING
C1253 _066_ VGND 12.4f $ **FLOATING
C1254 tdc0.r_dly_store_ring[21] VGND 0.948f $ **FLOATING
C1255 _074_ VGND 1.9f $ **FLOATING
C1256 a_14599_10927# VGND 0.609f $ **FLOATING
C1257 a_14767_10901# VGND 0.817f $ **FLOATING
C1258 a_14174_10927# VGND 0.626f $ **FLOATING
C1259 a_14342_10901# VGND 0.581f $ **FLOATING
C1260 a_13901_10933# VGND 1.43f $ **FLOATING
C1261 tdc0.w_ring_buf[21] VGND 0.872f $ **FLOATING
C1262 a_13735_10933# VGND 1.81f $ **FLOATING
C1263 a_13459_10927# VGND 0.524f $ **FLOATING
C1264 net39 VGND 8.62f $ **FLOATING
C1265 tdc0.w_ring_norsz[21] VGND 3.17f $ **FLOATING
C1266 tdc0.w_ring_norsz[5] VGND 4.35f $ **FLOATING
C1267 tdc0.w_ring_int_norsz[22] VGND 1.11f $ **FLOATING
C1268 a_10275_10927# VGND 0.609f $ **FLOATING
C1269 a_10443_10901# VGND 0.817f $ **FLOATING
C1270 a_9850_10927# VGND 0.626f $ **FLOATING
C1271 a_10018_10901# VGND 0.581f $ **FLOATING
C1272 a_9577_10933# VGND 1.43f $ **FLOATING
C1273 tdc0.w_ring_buf[24] VGND 0.872f $ **FLOATING
C1274 a_9411_10933# VGND 1.81f $ **FLOATING
C1275 a_9135_10927# VGND 0.524f $ **FLOATING
C1276 tdc0.w_ring_norsz[8] VGND 4.39f $ **FLOATING
C1277 tdc0.w_ring_int_norsz[8] VGND 1.07f $ **FLOATING
C1278 tdc0.w_ring_norsz[7] VGND 3.83f $ **FLOATING
C1279 a_5871_11146# VGND 0.524f $ **FLOATING
C1280 a_5043_11146# VGND 0.524f $ **FLOATING
C1281 a_2894_10927# VGND 0.653f $ **FLOATING
C1282 a_2963_10901# VGND 0.714f $ **FLOATING
C1283 a_2768_11043# VGND 1.57f $ **FLOATING
C1284 a_2807_11169# VGND 1.92f $ **FLOATING
C1285 a_2490_11059# VGND 0.736f $ **FLOATING
C1286 a_2287_10901# VGND 0.971f $ **FLOATING
C1287 a_26251_11471# VGND 0.319f $ **FLOATING
C1288 tdc0.w_ring_buf[27] VGND 1.5f $ **FLOATING
C1289 tdc0.w_ring_int_norsz[20] VGND 0.897f $ **FLOATING
C1290 a_27535_11471# VGND 0.524f $ **FLOATING
C1291 a_26420_11721# VGND 1.33f $ **FLOATING
C1292 _098_ VGND 1.76f $ **FLOATING
C1293 a_25971_11471# VGND 0.524f $ **FLOATING
C1294 a_23855_11471# VGND 0.524f $ **FLOATING
C1295 tdc0.w_ring_norsz[3] VGND 2.37f $ **FLOATING
C1296 net47 VGND 0.822f $ **FLOATING
C1297 tdc0.g_ring3[20].stg01_47.HI VGND 0.415f $ **FLOATING
C1298 tdc0.g_ring3[27].stg01_54.HI VGND 0.415f $ **FLOATING
C1299 tdc0.r_dly_store_ring[12] VGND 1.29f $ **FLOATING
C1300 tdc0.g_ring3[26].stg01_53.HI VGND 0.415f $ **FLOATING
C1301 a_20253_11471# VGND 0.23f $ **FLOATING
C1302 a_20763_11837# VGND 0.609f $ **FLOATING
C1303 a_20931_11739# VGND 0.817f $ **FLOATING
C1304 a_20338_11837# VGND 0.626f $ **FLOATING
C1305 a_20506_11583# VGND 0.581f $ **FLOATING
C1306 a_20065_11471# VGND 1.43f $ **FLOATING
C1307 tdc0.w_ring_buf[12] VGND 0.954f $ **FLOATING
C1308 a_19899_11471# VGND 1.81f $ **FLOATING
C1309 tdc0.w_ring_int_norsz[28] VGND 1.1f $ **FLOATING
C1310 a_15479_11721# VGND 0.253f $ **FLOATING
C1311 tdc0.g_ring3[22].stg01_49.HI VGND 0.415f $ **FLOATING
C1312 _114_ VGND 1.18f $ **FLOATING
C1313 _190_ VGND 1.13f $ **FLOATING
C1314 a_13645_11721# VGND 0.253f $ **FLOATING
C1315 net53 VGND 0.939f $ **FLOATING
C1316 tdc0.w_ring_norsz[25] VGND 2.16f $ **FLOATING
C1317 tdc0.w_ring_int_norsz[9] VGND 2.87f $ **FLOATING
C1318 a_15261_11445# VGND 0.55f $ **FLOATING
C1319 a_13814_11471# VGND 0.55f $ **FLOATING
C1320 net49 VGND 1.38f $ **FLOATING
C1321 tdc0.g_ring3[25].stg01_52.HI VGND 0.415f $ **FLOATING
C1322 tdc0.w_ring_int_norsz[25] VGND 2.81f $ **FLOATING
C1323 a_11233_11721# VGND 0.214f $ **FLOATING
C1324 a_11149_11721# VGND 0.167f $ **FLOATING
C1325 tdc0.g_ring3[23].stg01_50.HI VGND 0.415f $ **FLOATING
C1326 net52 VGND 0.822f $ **FLOATING
C1327 tdc0.w_ring_norsz[24] VGND 4.63f $ **FLOATING
C1328 tdc0.w_ring_int_norsz[6] VGND 0.897f $ **FLOATING
C1329 a_11067_11471# VGND 0.972f $ **FLOATING
C1330 tdc0.g_ring3[24].stg01_51.HI VGND 0.415f $ **FLOATING
C1331 tdc0.w_ring_int_norsz[23] VGND 1.61f $ **FLOATING
C1332 net50 VGND 0.931f $ **FLOATING
C1333 a_8723_11636# VGND 0.524f $ **FLOATING
C1334 tdc0.w_ring_int_norsz[7] VGND 1.14f $ **FLOATING
C1335 tdc0.w_ring_int_norsz[24] VGND 1.43f $ **FLOATING
C1336 tdc0.w_ring_buf[15] VGND 1.46f $ **FLOATING
C1337 tdc0.r_dly_store_ring[16] VGND 3.02f $ **FLOATING
C1338 a_5257_11471# VGND 0.23f $ **FLOATING
C1339 tdc0.w_ring_norsz[6] VGND 3.59f $ **FLOATING
C1340 net51 VGND 1.01f $ **FLOATING
C1341 tdc0.w_ring_norsz[23] VGND 2.39f $ **FLOATING
C1342 a_6791_11636# VGND 0.524f $ **FLOATING
C1343 a_5767_11837# VGND 0.609f $ **FLOATING
C1344 a_5935_11739# VGND 0.817f $ **FLOATING
C1345 a_5342_11837# VGND 0.626f $ **FLOATING
C1346 a_5510_11583# VGND 0.581f $ **FLOATING
C1347 a_5069_11471# VGND 1.43f $ **FLOATING
C1348 a_4903_11471# VGND 1.81f $ **FLOATING
C1349 tdc0.w_ring_buf[16] VGND 1.32f $ **FLOATING
C1350 _047_ VGND 1.93f $ **FLOATING
C1351 _006_ VGND 1.25f $ **FLOATING
C1352 a_3505_11721# VGND 0.219f $ **FLOATING
C1353 a_4627_11471# VGND 0.524f $ **FLOATING
C1354 a_3255_11721# VGND 0.684f $ **FLOATING
C1355 tdc0.r_ring_ctr[15] VGND 2.34f $ **FLOATING
C1356 a_28885_12393# VGND 0.23f $ **FLOATING
C1357 a_25493_12015# VGND 0.214f $ **FLOATING
C1358 a_25409_12015# VGND 0.167f $ **FLOATING
C1359 a_26785_12015# VGND 0.23f $ **FLOATING
C1360 _093_ VGND 1.16f $ **FLOATING
C1361 a_24209_12015# VGND 0.23f $ **FLOATING
C1362 tdc0.w_ring_int_norsz[19] VGND 0.931f $ **FLOATING
C1363 tdc0.w_ring_int_norsz[3] VGND 1.02f $ **FLOATING
C1364 tdc0.w_ring_buf[26] VGND 1.52f $ **FLOATING
C1365 a_28467_12393# VGND 0.581f $ **FLOATING
C1366 a_28538_12292# VGND 0.626f $ **FLOATING
C1367 a_28338_12137# VGND 1.43f $ **FLOATING
C1368 a_28331_12233# VGND 1.81f $ **FLOATING
C1369 a_28047_12247# VGND 0.609f $ **FLOATING
C1370 a_27951_12247# VGND 0.817f $ **FLOATING
C1371 a_27295_12015# VGND 0.609f $ **FLOATING
C1372 a_27463_11989# VGND 0.817f $ **FLOATING
C1373 a_26870_12015# VGND 0.626f $ **FLOATING
C1374 a_27038_11989# VGND 0.581f $ **FLOATING
C1375 a_26597_12021# VGND 1.43f $ **FLOATING
C1376 tdc0.w_ring_buf[18] VGND 0.911f $ **FLOATING
C1377 a_26431_12021# VGND 1.81f $ **FLOATING
C1378 a_26063_12015# VGND 0.524f $ **FLOATING
C1379 a_25327_12015# VGND 0.972f $ **FLOATING
C1380 tdc0.r_dly_store_ring[2] VGND 0.788f $ **FLOATING
C1381 _086_ VGND 18.9f $ **FLOATING
C1382 a_24719_12015# VGND 0.609f $ **FLOATING
C1383 a_24887_11989# VGND 0.817f $ **FLOATING
C1384 a_24294_12015# VGND 0.626f $ **FLOATING
C1385 a_24462_11989# VGND 0.581f $ **FLOATING
C1386 a_24021_12021# VGND 1.43f $ **FLOATING
C1387 tdc0.w_ring_buf[2] VGND 1.01f $ **FLOATING
C1388 a_23855_12021# VGND 1.81f $ **FLOATING
C1389 tdc0.w_ring_norsz[2] VGND 2.33f $ **FLOATING
C1390 tdc0.w_ring_norsz[18] VGND 3.22f $ **FLOATING
C1391 net54 VGND 1.25f $ **FLOATING
C1392 tdc0.w_ring_int_norsz[27] VGND 0.714f $ **FLOATING
C1393 tdc0.w_ring_norsz[27] VGND 4.82f $ **FLOATING
C1394 tdc0.w_ring_int_norsz[11] VGND 0.761f $ **FLOATING
C1395 tdc0.g_ring3[28].stg01_55.HI VGND 0.415f $ **FLOATING
C1396 net55 VGND 1.4f $ **FLOATING
C1397 tdc0.w_ring_norsz[12] VGND 2.35f $ **FLOATING
C1398 net12 VGND 4.82f $ **FLOATING
C1399 tdc0.w_ring_int_norsz[12] VGND 0.831f $ **FLOATING
C1400 a_19255_12015# VGND 0.524f $ **FLOATING
C1401 tdc0.w_ring_norsz[26] VGND 1.4f $ **FLOATING
C1402 tdc0.w_ring_int_norsz[10] VGND 0.917f $ **FLOATING
C1403 tdc0.w_ring_int_norsz[26] VGND 0.962f $ **FLOATING
C1404 net41 VGND 11.7f $ **FLOATING
C1405 tdc0.w_ring_norsz[9] VGND 2.06f $ **FLOATING
C1406 a_17923_12234# VGND 0.524f $ **FLOATING
C1407 tdc0.g_ring3[29].stg01_56.HI VGND 0.415f $ **FLOATING
C1408 tdc0.w_ring_int_norsz[18] VGND 3.53f $ **FLOATING
C1409 tdc0.r_dly_store_ring[13] VGND 0.909f $ **FLOATING
C1410 a_14457_12015# VGND 0.23f $ **FLOATING
C1411 a_11623_12335# VGND 0.319f $ **FLOATING
C1412 tdc0.r_dly_store_ring[14] VGND 1.11f $ **FLOATING
C1413 a_9765_12015# VGND 0.23f $ **FLOATING
C1414 tdc0.r_dly_store_ring[6] VGND 1.64f $ **FLOATING
C1415 a_8293_12015# VGND 0.23f $ **FLOATING
C1416 tdc0.w_ring_norsz[28] VGND 3.61f $ **FLOATING
C1417 net56 VGND 0.931f $ **FLOATING
C1418 tdc0.w_ring_int_norsz[1] VGND 0.722f $ **FLOATING
C1419 a_15809_12234# VGND 0.524f $ **FLOATING
C1420 a_14967_12015# VGND 0.609f $ **FLOATING
C1421 a_15135_11989# VGND 0.817f $ **FLOATING
C1422 a_14542_12015# VGND 0.626f $ **FLOATING
C1423 a_14710_11989# VGND 0.581f $ **FLOATING
C1424 a_14269_12021# VGND 1.43f $ **FLOATING
C1425 a_14103_12021# VGND 1.81f $ **FLOATING
C1426 tdc0.w_ring_int_norsz[29] VGND 2.2f $ **FLOATING
C1427 tdc0.w_ring_int_norsz[13] VGND 3.39f $ **FLOATING
C1428 a_11792_12015# VGND 1.33f $ **FLOATING
C1429 _130_ VGND 3.32f $ **FLOATING
C1430 _125_ VGND 0.993f $ **FLOATING
C1431 a_10975_12015# VGND 0.524f $ **FLOATING
C1432 tdc0.w_ring_norsz[22] VGND 3.62f $ **FLOATING
C1433 a_10275_12015# VGND 0.609f $ **FLOATING
C1434 a_10443_11989# VGND 0.817f $ **FLOATING
C1435 a_9850_12015# VGND 0.626f $ **FLOATING
C1436 a_10018_11989# VGND 0.581f $ **FLOATING
C1437 a_9577_12021# VGND 1.43f $ **FLOATING
C1438 a_9411_12021# VGND 1.81f $ **FLOATING
C1439 a_8803_12015# VGND 0.609f $ **FLOATING
C1440 a_8971_11989# VGND 0.817f $ **FLOATING
C1441 a_8378_12015# VGND 0.626f $ **FLOATING
C1442 a_8546_11989# VGND 0.581f $ **FLOATING
C1443 a_8105_12021# VGND 1.43f $ **FLOATING
C1444 tdc0.w_ring_buf[6] VGND 1.16f $ **FLOATING
C1445 a_7939_12021# VGND 1.81f $ **FLOATING
C1446 tdc0.w_ring_int_norsz[31] VGND 0.923f $ **FLOATING
C1447 tdc0.w_ring_int_norsz[15] VGND 0.878f $ **FLOATING
C1448 tdc0.w_ring_norsz[15] VGND 2.74f $ **FLOATING
C1449 tdc0.w_ring_int_norsz[16] VGND 2.39f $ **FLOATING
C1450 tdc0.w_ring_norsz[16] VGND 4.05f $ **FLOATING
C1451 a_3399_12275# VGND 1.2f $ **FLOATING
C1452 _092_ VGND 1.96f $ **FLOATING
C1453 a_27057_12809# VGND 0.214f $ **FLOATING
C1454 a_26973_12809# VGND 0.167f $ **FLOATING
C1455 a_24029_12809# VGND 0.206f $ **FLOATING
C1456 a_26891_12559# VGND 0.972f $ **FLOATING
C1457 tdc0.r_dly_store_ring[26] VGND 1.05f $ **FLOATING
C1458 tdc0.r_dly_store_ring[18] VGND 1.23f $ **FLOATING
C1459 a_24775_12559# VGND 0.524f $ **FLOATING
C1460 tdc0.w_ring_norsz[10] VGND 4.65f $ **FLOATING
C1461 a_23947_12809# VGND 0.804f $ **FLOATING
C1462 a_23303_12559# VGND 0.524f $ **FLOATING
C1463 tdc0.w_ring_norsz[19] VGND 2.23f $ **FLOATING
C1464 net46 VGND 1.57f $ **FLOATING
C1465 tdc0.g_ring3[19].stg01_46.HI VGND 0.415f $ **FLOATING
C1466 tdc0.w_ring_int_norsz[2] VGND 0.897f $ **FLOATING
C1467 _090_ VGND 3.21f $ **FLOATING
C1468 a_21270_12809# VGND 0.191f $ **FLOATING
C1469 a_19977_12559# VGND 0.23f $ **FLOATING
C1470 net40 VGND 10.4f $ **FLOATING
C1471 a_21739_12559# VGND 0.524f $ **FLOATING
C1472 tdc0.w_ring_norsz[11] VGND 2.42f $ **FLOATING
C1473 a_21095_12559# VGND 0.847f $ **FLOATING
C1474 _083_ VGND 16.9f $ **FLOATING
C1475 tdc0.r_dly_store_ring[1] VGND 0.765f $ **FLOATING
C1476 a_20487_12925# VGND 0.609f $ **FLOATING
C1477 a_20655_12827# VGND 0.817f $ **FLOATING
C1478 a_20062_12925# VGND 0.626f $ **FLOATING
C1479 a_20230_12671# VGND 0.581f $ **FLOATING
C1480 a_19789_12559# VGND 1.43f $ **FLOATING
C1481 a_19623_12559# VGND 1.81f $ **FLOATING
C1482 tdc0.w_ring_buf[1] VGND 0.872f $ **FLOATING
C1483 a_17493_12559# VGND 0.23f $ **FLOATING
C1484 a_19347_12559# VGND 0.524f $ **FLOATING
C1485 a_18003_12925# VGND 0.609f $ **FLOATING
C1486 a_18171_12827# VGND 0.817f $ **FLOATING
C1487 a_17578_12925# VGND 0.626f $ **FLOATING
C1488 a_17746_12671# VGND 0.581f $ **FLOATING
C1489 a_17305_12559# VGND 1.43f $ **FLOATING
C1490 tdc0.w_ring_buf[9] VGND 1.11f $ **FLOATING
C1491 a_17139_12559# VGND 1.81f $ **FLOATING
C1492 net1 VGND 10.7f $ **FLOATING
C1493 a_16463_12533# VGND 1.2f $ **FLOATING
C1494 tdc0.w_ring_norsz[1] VGND 4.52f $ **FLOATING
C1495 tdc0.w_ring_int_norsz[17] VGND 5.97f $ **FLOATING
C1496 net45 VGND 1.6f $ **FLOATING
C1497 tdc0.g_ring3[18].stg01_45.HI VGND 0.415f $ **FLOATING
C1498 tdc0.w_ring_buf[13] VGND 1.03f $ **FLOATING
C1499 tdc0.w_ring_int_norsz[14] VGND 0.936f $ **FLOATING
C1500 _124_ VGND 1.38f $ **FLOATING
C1501 a_11601_12809# VGND 0.214f $ **FLOATING
C1502 a_11517_12809# VGND 0.167f $ **FLOATING
C1503 tdc0.w_ring_buf[14] VGND 0.968f $ **FLOATING
C1504 tdc0.g_ring3[31].stg01_58.HI VGND 0.415f $ **FLOATING
C1505 a_15483_12559# VGND 0.524f $ **FLOATING
C1506 tdc0.w_ring_norsz[17] VGND 2.41f $ **FLOATING
C1507 a_14703_12724# VGND 0.524f $ **FLOATING
C1508 a_14427_12724# VGND 0.524f $ **FLOATING
C1509 a_13735_12559# VGND 1.2f $ **FLOATING
C1510 tdc0.w_ring_norsz[13] VGND 2.73f $ **FLOATING
C1511 net38 VGND 13.9f $ **FLOATING
C1512 tdc0.w_ring_norsz[29] VGND 2.6f $ **FLOATING
C1513 tdc0.w_ring_int_norsz[30] VGND 0.722f $ **FLOATING
C1514 a_11435_12559# VGND 0.972f $ **FLOATING
C1515 tdc0.w_ring_norsz[14] VGND 4.07f $ **FLOATING
C1516 a_9643_12724# VGND 0.524f $ **FLOATING
C1517 a_8583_12559# VGND 0.524f $ **FLOATING
C1518 tdc0.w_ring_norsz[30] VGND 4.63f $ **FLOATING
C1519 net58 VGND 1.31f $ **FLOATING
C1520 tdc0.stg01_59.HI VGND 0.415f $ **FLOATING
C1521 a_6545_12559# VGND 0.23f $ **FLOATING
C1522 a_7055_12925# VGND 0.609f $ **FLOATING
C1523 a_7223_12827# VGND 0.817f $ **FLOATING
C1524 a_6630_12925# VGND 0.626f $ **FLOATING
C1525 a_6798_12671# VGND 0.581f $ **FLOATING
C1526 a_6357_12559# VGND 1.43f $ **FLOATING
C1527 a_6191_12559# VGND 1.81f $ **FLOATING
C1528 tdc0.w_ring_int_norsz[0] VGND 0.889f $ **FLOATING
C1529 net11 VGND 6.11f $ **FLOATING
C1530 a_3871_12925# VGND 0.168f $ **FLOATING
C1531 a_3668_12559# VGND 0.259f $ **FLOATING
C1532 tdc0.w_ring_norsz[31] VGND 3.19f $ **FLOATING
C1533 net59 VGND 0.931f $ **FLOATING
C1534 a_5271_12559# VGND 0.524f $ **FLOATING
C1535 tdc0.w_ring_norsz[0] VGND 1.87f $ **FLOATING
C1536 a_4328_12559# VGND 0.736f $ **FLOATING
C1537 a_4503_12533# VGND 0.971f $ **FLOATING
C1538 a_3763_12559# VGND 0.714f $ **FLOATING
C1539 _046_ VGND 1.7f $ **FLOATING
C1540 a_3981_12801# VGND 0.653f $ **FLOATING
C1541 a_3413_12559# VGND 1.57f $ **FLOATING
C1542 a_3247_12559# VGND 1.92f $ **FLOATING
C1543 _622_.X VGND 0.226f $ **FLOATING
C1544 a_2840_12533# VGND 0.648f $ **FLOATING
C1545 a_26513_13103# VGND 0.206f $ **FLOATING
C1546 _091_ VGND 0.828f $ **FLOATING
C1547 a_25221_13103# VGND 0.23f $ **FLOATING
C1548 tdc0.r_dly_store_ring[19] VGND 1f $ **FLOATING
C1549 a_23565_13103# VGND 0.23f $ **FLOATING
C1550 tdc0.r_dly_store_ring[11] VGND 1.16f $ **FLOATING
C1551 a_20341_13103# VGND 0.214f $ **FLOATING
C1552 a_20257_13103# VGND 0.167f $ **FLOATING
C1553 a_18877_13103# VGND 0.206f $ **FLOATING
C1554 a_22093_13103# VGND 0.23f $ **FLOATING
C1555 _088_ VGND 0.955f $ **FLOATING
C1556 _089_ VGND 1.54f $ **FLOATING
C1557 a_15105_13103# VGND 0.206f $ **FLOATING
C1558 a_16757_13103# VGND 0.23f $ **FLOATING
C1559 _116_ VGND 2.23f $ **FLOATING
C1560 a_13905_13103# VGND 0.23f $ **FLOATING
C1561 a_26431_13103# VGND 0.804f $ **FLOATING
C1562 tdc0.r_dly_store_ring[10] VGND 0.669f $ **FLOATING
C1563 a_25731_13103# VGND 0.609f $ **FLOATING
C1564 a_25899_13077# VGND 0.817f $ **FLOATING
C1565 a_25306_13103# VGND 0.626f $ **FLOATING
C1566 a_25474_13077# VGND 0.581f $ **FLOATING
C1567 a_25033_13109# VGND 1.43f $ **FLOATING
C1568 tdc0.w_ring_buf[10] VGND 1.05f $ **FLOATING
C1569 a_24867_13109# VGND 1.81f $ **FLOATING
C1570 a_24075_13103# VGND 0.609f $ **FLOATING
C1571 a_24243_13077# VGND 0.817f $ **FLOATING
C1572 a_23650_13103# VGND 0.626f $ **FLOATING
C1573 a_23818_13077# VGND 0.581f $ **FLOATING
C1574 a_23377_13109# VGND 1.43f $ **FLOATING
C1575 tdc0.w_ring_buf[19] VGND 0.961f $ **FLOATING
C1576 a_23211_13109# VGND 1.81f $ **FLOATING
C1577 a_22603_13103# VGND 0.609f $ **FLOATING
C1578 a_22771_13077# VGND 0.817f $ **FLOATING
C1579 a_22178_13103# VGND 0.626f $ **FLOATING
C1580 a_22346_13077# VGND 0.581f $ **FLOATING
C1581 a_21905_13109# VGND 1.43f $ **FLOATING
C1582 tdc0.w_ring_buf[11] VGND 1.01f $ **FLOATING
C1583 a_21739_13109# VGND 1.81f $ **FLOATING
C1584 a_20175_13103# VGND 0.972f $ **FLOATING
C1585 _087_ VGND 2.11f $ **FLOATING
C1586 a_18795_13103# VGND 0.804f $ **FLOATING
C1587 _067_ VGND 19.1f $ **FLOATING
C1588 tdc0.r_dly_store_ring[17] VGND 1.18f $ **FLOATING
C1589 _072_ VGND 18.3f $ **FLOATING
C1590 tdc0.r_dly_store_ring[9] VGND 0.915f $ **FLOATING
C1591 a_17267_13103# VGND 0.609f $ **FLOATING
C1592 a_17435_13077# VGND 0.817f $ **FLOATING
C1593 a_16842_13103# VGND 0.626f $ **FLOATING
C1594 a_17010_13077# VGND 0.581f $ **FLOATING
C1595 a_16569_13109# VGND 1.43f $ **FLOATING
C1596 tdc0.w_ring_buf[17] VGND 1.39f $ **FLOATING
C1597 a_16403_13109# VGND 1.81f $ **FLOATING
C1598 a_15023_13103# VGND 0.804f $ **FLOATING
C1599 tdc0.r_dly_store_ring[29] VGND 0.76f $ **FLOATING
C1600 a_14415_13103# VGND 0.609f $ **FLOATING
C1601 a_14583_13077# VGND 0.817f $ **FLOATING
C1602 a_13990_13103# VGND 0.626f $ **FLOATING
C1603 a_14158_13077# VGND 0.581f $ **FLOATING
C1604 a_13717_13109# VGND 1.43f $ **FLOATING
C1605 tdc0.w_ring_buf[29] VGND 1.34f $ **FLOATING
C1606 a_13551_13109# VGND 1.81f $ **FLOATING
C1607 tdc0.g_ring3[30].stg01_57.HI VGND 0.415f $ **FLOATING
C1608 net57 VGND 1.18f $ **FLOATING
C1609 a_12529_13103# VGND 0.206f $ **FLOATING
C1610 _110_ VGND 5.8f $ **FLOATING
C1611 tdc0.r_dly_store_ring[22] VGND 1.07f $ **FLOATING
C1612 a_10229_13103# VGND 0.206f $ **FLOATING
C1613 a_11329_13103# VGND 0.23f $ **FLOATING
C1614 _123_ VGND 1.1f $ **FLOATING
C1615 a_9029_13103# VGND 0.23f $ **FLOATING
C1616 tdc0.r_dly_store_ctr[13] VGND 3.57f $ **FLOATING
C1617 a_7557_13103# VGND 0.23f $ **FLOATING
C1618 a_12447_13103# VGND 0.804f $ **FLOATING
C1619 tdc0.r_dly_store_ctr[12] VGND 2.9f $ **FLOATING
C1620 a_11839_13103# VGND 0.609f $ **FLOATING
C1621 a_12007_13077# VGND 0.817f $ **FLOATING
C1622 a_11414_13103# VGND 0.626f $ **FLOATING
C1623 a_11582_13077# VGND 0.581f $ **FLOATING
C1624 a_11141_13109# VGND 1.43f $ **FLOATING
C1625 tdc0.w_ring_buf[22] VGND 1.22f $ **FLOATING
C1626 a_10975_13109# VGND 1.81f $ **FLOATING
C1627 a_10147_13103# VGND 0.804f $ **FLOATING
C1628 _069_ VGND 20.3f $ **FLOATING
C1629 tdc0.r_dly_store_ring[30] VGND 0.786f $ **FLOATING
C1630 a_9539_13103# VGND 0.609f $ **FLOATING
C1631 a_9707_13077# VGND 0.817f $ **FLOATING
C1632 a_9114_13103# VGND 0.626f $ **FLOATING
C1633 a_9282_13077# VGND 0.581f $ **FLOATING
C1634 a_8841_13109# VGND 1.43f $ **FLOATING
C1635 tdc0.w_ring_buf[30] VGND 1.03f $ **FLOATING
C1636 a_8675_13109# VGND 1.81f $ **FLOATING
C1637 a_8067_13103# VGND 0.609f $ **FLOATING
C1638 a_8235_13077# VGND 0.817f $ **FLOATING
C1639 a_7642_13103# VGND 0.626f $ **FLOATING
C1640 a_7810_13077# VGND 0.581f $ **FLOATING
C1641 a_7369_13109# VGND 1.43f $ **FLOATING
C1642 a_7203_13109# VGND 1.81f $ **FLOATING
C1643 tdc0.g_ring3[16].stg01_43.HI VGND 0.415f $ **FLOATING
C1644 net43 VGND 1.27f $ **FLOATING
C1645 tdc0.g_ring1[16].stg02_42.HI VGND 0.415f $ **FLOATING
C1646 net42 VGND 1.7f $ **FLOATING
C1647 tdc0.g_ring3[17].stg01_44.HI VGND 0.415f $ **FLOATING
C1648 net44 VGND 1.43f $ **FLOATING
C1649 _005_ VGND 1.39f $ **FLOATING
C1650 net21 VGND 9.82f $ **FLOATING
C1651 a_3799_13103# VGND 0.698f $ **FLOATING
C1652 tdc0.w_dly_stop[5] VGND 0.844f $ **FLOATING
C1653 net24 VGND 12.8f $ **FLOATING
C1654 a_3484_13077# VGND 0.648f $ **FLOATING
C1655 a_3155_13103# VGND 0.524f $ **FLOATING
C1656 a_2787_13103# VGND 0.524f $ **FLOATING
C1657 _104_ VGND 2.29f $ **FLOATING
C1658 a_24849_13897# VGND 0.214f $ **FLOATING
C1659 a_24765_13897# VGND 0.167f $ **FLOATING
C1660 a_22001_13647# VGND 0.23f $ **FLOATING
C1661 a_24683_13647# VGND 0.972f $ **FLOATING
C1662 _075_ VGND 21.6f $ **FLOATING
C1663 _077_ VGND 23f $ **FLOATING
C1664 tdc0.r_dly_store_ctr[11] VGND 1.33f $ **FLOATING
C1665 _103_ VGND 1.05f $ **FLOATING
C1666 a_22511_14013# VGND 0.609f $ **FLOATING
C1667 a_22679_13915# VGND 0.817f $ **FLOATING
C1668 a_22086_14013# VGND 0.626f $ **FLOATING
C1669 a_22254_13759# VGND 0.581f $ **FLOATING
C1670 a_21813_13647# VGND 1.43f $ **FLOATING
C1671 a_21647_13647# VGND 1.81f $ **FLOATING
C1672 a_21157_13647# VGND 0.23f $ **FLOATING
C1673 tdc0.r_dly_store_ctr[1] VGND 0.958f $ **FLOATING
C1674 tdc0.r_dly_store_ctr[9] VGND 0.849f $ **FLOATING
C1675 a_19057_13647# VGND 0.23f $ **FLOATING
C1676 a_20739_13647# VGND 0.581f $ **FLOATING
C1677 a_20810_13621# VGND 0.626f $ **FLOATING
C1678 a_20603_13621# VGND 1.81f $ **FLOATING
C1679 a_20610_13921# VGND 1.43f $ **FLOATING
C1680 a_20319_13621# VGND 0.609f $ **FLOATING
C1681 a_20223_13799# VGND 0.817f $ **FLOATING
C1682 a_19567_14013# VGND 0.609f $ **FLOATING
C1683 a_19735_13915# VGND 0.817f $ **FLOATING
C1684 a_19142_14013# VGND 0.626f $ **FLOATING
C1685 a_19310_13759# VGND 0.581f $ **FLOATING
C1686 a_18869_13647# VGND 1.43f $ **FLOATING
C1687 a_18703_13647# VGND 1.81f $ **FLOATING
C1688 a_18029_13647# VGND 0.23f $ **FLOATING
C1689 tdc0.r_dly_store_ctr[0] VGND 3.3f $ **FLOATING
C1690 a_15647_14013# VGND 0.168f $ **FLOATING
C1691 a_15444_13647# VGND 0.259f $ **FLOATING
C1692 a_17611_13647# VGND 0.581f $ **FLOATING
C1693 a_17682_13621# VGND 0.626f $ **FLOATING
C1694 a_17475_13621# VGND 1.81f $ **FLOATING
C1695 a_17482_13921# VGND 1.43f $ **FLOATING
C1696 a_17191_13621# VGND 0.609f $ **FLOATING
C1697 a_17095_13799# VGND 0.817f $ **FLOATING
C1698 a_16104_13647# VGND 0.736f $ **FLOATING
C1699 a_16279_13621# VGND 0.971f $ **FLOATING
C1700 a_15539_13647# VGND 0.714f $ **FLOATING
C1701 _043_ VGND 2.01f $ **FLOATING
C1702 a_15757_13889# VGND 0.653f $ **FLOATING
C1703 a_15189_13647# VGND 1.57f $ **FLOATING
C1704 a_15023_13647# VGND 1.92f $ **FLOATING
C1705 tdc0.r_dly_store_ctr[8] VGND 2.18f $ **FLOATING
C1706 a_13905_13647# VGND 0.23f $ **FLOATING
C1707 a_14415_14013# VGND 0.609f $ **FLOATING
C1708 a_14583_13915# VGND 0.817f $ **FLOATING
C1709 a_13990_14013# VGND 0.626f $ **FLOATING
C1710 a_14158_13759# VGND 0.581f $ **FLOATING
C1711 a_13717_13647# VGND 1.43f $ **FLOATING
C1712 a_13551_13647# VGND 1.81f $ **FLOATING
C1713 tdc0.r_dly_store_ctr[6] VGND 1.14f $ **FLOATING
C1714 a_10225_13647# VGND 0.23f $ **FLOATING
C1715 a_10735_14013# VGND 0.609f $ **FLOATING
C1716 a_10903_13915# VGND 0.817f $ **FLOATING
C1717 a_10310_14013# VGND 0.626f $ **FLOATING
C1718 a_10478_13759# VGND 0.581f $ **FLOATING
C1719 a_10037_13647# VGND 1.43f $ **FLOATING
C1720 a_9871_13647# VGND 1.81f $ **FLOATING
C1721 a_6739_13897# VGND 0.253f $ **FLOATING
C1722 tdc0.r_dly_store_ctr[14] VGND 2.55f $ **FLOATING
C1723 a_5349_13647# VGND 0.23f $ **FLOATING
C1724 a_6521_13621# VGND 0.55f $ **FLOATING
C1725 a_5859_14013# VGND 0.609f $ **FLOATING
C1726 a_6027_13915# VGND 0.817f $ **FLOATING
C1727 a_5434_14013# VGND 0.626f $ **FLOATING
C1728 a_5602_13759# VGND 0.581f $ **FLOATING
C1729 a_5161_13647# VGND 1.43f $ **FLOATING
C1730 a_4995_13647# VGND 1.81f $ **FLOATING
C1731 _161_ VGND 2.87f $ **FLOATING
C1732 _162_ VGND 0.883f $ **FLOATING
C1733 a_3789_13897# VGND 0.184f $ **FLOATING
C1734 a_4219_13621# VGND 0.729f $ **FLOATING
C1735 tdc0.r_ring_ctr[14] VGND 2.33f $ **FLOATING
C1736 a_3247_13647# VGND 0.648f $ **FLOATING
C1737 tdc0.w_dly_stop[4] VGND 0.871f $ **FLOATING
C1738 tdc0.w_dly_stop[2] VGND 0.834f $ **FLOATING
C1739 a_2879_13647# VGND 0.524f $ **FLOATING
C1740 tdc0.w_dly_stop[3] VGND 0.864f $ **FLOATING
C1741 a_2603_13647# VGND 0.524f $ **FLOATING
C1742 tdc0.w_dly_stop[1] VGND 0.683f $ **FLOATING
C1743 a_2327_13647# VGND 0.524f $ **FLOATING
C1744 tdc0.r_dly_store_ctr[2] VGND 1.19f $ **FLOATING
C1745 a_25221_14191# VGND 0.23f $ **FLOATING
C1746 tdc0.r_dly_store_ctr[10] VGND 1.76f $ **FLOATING
C1747 a_23749_14191# VGND 0.23f $ **FLOATING
C1748 a_18039_14191# VGND 0.168f $ **FLOATING
C1749 a_17836_14557# VGND 0.259f $ **FLOATING
C1750 net32 VGND 11.4f $ **FLOATING
C1751 a_15569_14511# VGND 0.171f $ **FLOATING
C1752 _002_ VGND 1.07f $ **FLOATING
C1753 tdc0.r_dly_store_ctr[5] VGND 2.12f $ **FLOATING
C1754 a_13629_14191# VGND 0.23f $ **FLOATING
C1755 tdc0.r_dly_store_ctr[4] VGND 0.992f $ **FLOATING
C1756 a_11697_14191# VGND 0.23f $ **FLOATING
C1757 tdc0.r_dly_store_ctr[7] VGND 2.34f $ **FLOATING
C1758 a_8569_14191# VGND 0.23f $ **FLOATING
C1759 a_6907_14191# VGND 0.168f $ **FLOATING
C1760 a_3689_14191# VGND 0.219f $ **FLOATING
C1761 a_6704_14557# VGND 0.259f $ **FLOATING
C1762 net2 VGND 2.19f $ **FLOATING
C1763 a_25731_14191# VGND 0.609f $ **FLOATING
C1764 a_25899_14165# VGND 0.817f $ **FLOATING
C1765 a_25306_14191# VGND 0.626f $ **FLOATING
C1766 a_25474_14165# VGND 0.581f $ **FLOATING
C1767 a_25033_14197# VGND 1.43f $ **FLOATING
C1768 a_24867_14197# VGND 1.81f $ **FLOATING
C1769 a_24259_14191# VGND 0.609f $ **FLOATING
C1770 a_24427_14165# VGND 0.817f $ **FLOATING
C1771 a_23834_14191# VGND 0.626f $ **FLOATING
C1772 a_24002_14165# VGND 0.581f $ **FLOATING
C1773 a_23561_14197# VGND 1.43f $ **FLOATING
C1774 a_23395_14197# VGND 1.81f $ **FLOATING
C1775 a_23080_14165# VGND 0.648f $ **FLOATING
C1776 a_18496_14569# VGND 0.736f $ **FLOATING
C1777 a_18671_14495# VGND 0.971f $ **FLOATING
C1778 a_17931_14569# VGND 0.714f $ **FLOATING
C1779 a_18149_14165# VGND 0.653f $ **FLOATING
C1780 a_17581_14197# VGND 1.57f $ **FLOATING
C1781 a_17415_14197# VGND 1.92f $ **FLOATING
C1782 a_17100_14165# VGND 0.648f $ **FLOATING
C1783 a_16127_14557# VGND 0.729f $ **FLOATING
C1784 tdc0.r_ring_ctr[11] VGND 4.51f $ **FLOATING
C1785 a_15351_14423# VGND 0.546f $ **FLOATING
C1786 a_14983_14165# VGND 0.698f $ **FLOATING
C1787 a_14139_14191# VGND 0.609f $ **FLOATING
C1788 a_14307_14165# VGND 0.817f $ **FLOATING
C1789 a_13714_14191# VGND 0.626f $ **FLOATING
C1790 a_13882_14165# VGND 0.581f $ **FLOATING
C1791 a_13441_14197# VGND 1.43f $ **FLOATING
C1792 a_13275_14197# VGND 1.81f $ **FLOATING
C1793 a_12207_14191# VGND 0.609f $ **FLOATING
C1794 a_12375_14165# VGND 0.817f $ **FLOATING
C1795 a_11782_14191# VGND 0.626f $ **FLOATING
C1796 a_11950_14165# VGND 0.581f $ **FLOATING
C1797 a_11509_14197# VGND 1.43f $ **FLOATING
C1798 a_11343_14197# VGND 1.81f $ **FLOATING
C1799 net29 VGND 12.5f $ **FLOATING
C1800 a_9924_14165# VGND 0.648f $ **FLOATING
C1801 a_9079_14191# VGND 0.609f $ **FLOATING
C1802 a_9247_14165# VGND 0.817f $ **FLOATING
C1803 a_8654_14191# VGND 0.626f $ **FLOATING
C1804 a_8822_14165# VGND 0.581f $ **FLOATING
C1805 a_8381_14197# VGND 1.43f $ **FLOATING
C1806 a_8215_14197# VGND 1.81f $ **FLOATING
C1807 net27 VGND 12.3f $ **FLOATING
C1808 a_7364_14569# VGND 0.736f $ **FLOATING
C1809 a_7539_14495# VGND 0.971f $ **FLOATING
C1810 a_6799_14569# VGND 0.714f $ **FLOATING
C1811 _045_ VGND 1.74f $ **FLOATING
C1812 a_7017_14165# VGND 0.653f $ **FLOATING
C1813 a_6449_14197# VGND 1.57f $ **FLOATING
C1814 a_6283_14197# VGND 1.92f $ **FLOATING
C1815 tdc0.r_ring_ctr[13] VGND 5.28f $ **FLOATING
C1816 net20 VGND 9.33f $ **FLOATING
C1817 a_3439_14191# VGND 0.684f $ **FLOATING
C1818 net28 VGND 12.3f $ **FLOATING
C1819 a_2932_14165# VGND 0.648f $ **FLOATING
C1820 a_2511_14191# VGND 0.698f $ **FLOATING
C1821 a_855_14191# VGND 0.524f $ **FLOATING
C1822 tdc0.r_dly_store_ctr[3] VGND 1.12f $ **FLOATING
C1823 a_24209_14735# VGND 0.23f $ **FLOATING
C1824 a_24719_15101# VGND 0.609f $ **FLOATING
C1825 a_24887_15003# VGND 0.817f $ **FLOATING
C1826 a_24294_15101# VGND 0.626f $ **FLOATING
C1827 a_24462_14847# VGND 0.581f $ **FLOATING
C1828 a_24021_14735# VGND 1.43f $ **FLOATING
C1829 a_23855_14735# VGND 1.81f $ **FLOATING
C1830 net35 VGND 10.2f $ **FLOATING
C1831 a_22271_15101# VGND 0.168f $ **FLOATING
C1832 a_22068_14735# VGND 0.259f $ **FLOATING
C1833 a_22728_14735# VGND 0.736f $ **FLOATING
C1834 a_22903_14709# VGND 0.971f $ **FLOATING
C1835 a_22163_14735# VGND 0.714f $ **FLOATING
C1836 _034_ VGND 1.61f $ **FLOATING
C1837 a_22381_14977# VGND 0.653f $ **FLOATING
C1838 a_21813_14735# VGND 1.57f $ **FLOATING
C1839 a_21647_14735# VGND 1.92f $ **FLOATING
C1840 _008_ VGND 1.15f $ **FLOATING
C1841 a_19715_14985# VGND 0.238f $ **FLOATING
C1842 _140_ VGND 1.2f $ **FLOATING
C1843 a_20727_14735# VGND 0.619f $ **FLOATING
C1844 a_20083_14735# VGND 0.729f $ **FLOATING
C1845 tdc0.r_ring_ctr[2] VGND 4.12f $ **FLOATING
C1846 a_19255_14735# VGND 0.648f $ **FLOATING
C1847 net23 VGND 9.72f $ **FLOATING
C1848 _042_ VGND 1.61f $ **FLOATING
C1849 net33 VGND 10.8f $ **FLOATING
C1850 _001_ VGND 1.45f $ **FLOATING
C1851 a_16845_14985# VGND 0.219f $ **FLOATING
C1852 _155_ VGND 0.931f $ **FLOATING
C1853 a_12243_15101# VGND 0.168f $ **FLOATING
C1854 a_12040_14735# VGND 0.259f $ **FLOATING
C1855 a_18703_14735# VGND 0.988f $ **FLOATING
C1856 net22 VGND 8.14f $ **FLOATING
C1857 a_17283_14709# VGND 0.698f $ **FLOATING
C1858 a_16595_14985# VGND 0.684f $ **FLOATING
C1859 _154_ VGND 1.39f $ **FLOATING
C1860 tdc0.r_ring_ctr[10] VGND 5.78f $ **FLOATING
C1861 a_15627_14709# VGND 0.729f $ **FLOATING
C1862 a_15115_14735# VGND 0.619f $ **FLOATING
C1863 a_12700_14735# VGND 0.736f $ **FLOATING
C1864 a_12875_14709# VGND 0.971f $ **FLOATING
C1865 a_12135_14735# VGND 0.714f $ **FLOATING
C1866 _037_ VGND 1.64f $ **FLOATING
C1867 a_12353_14977# VGND 0.653f $ **FLOATING
C1868 a_11785_14735# VGND 1.57f $ **FLOATING
C1869 a_11619_14735# VGND 1.92f $ **FLOATING
C1870 _158_ VGND 5.41f $ **FLOATING
C1871 a_6191_14735# VGND 0.171f $ **FLOATING
C1872 _004_ VGND 1.09f $ **FLOATING
C1873 tdc0.r_ring_ctr[12] VGND 6.04f $ **FLOATING
C1874 a_4423_15101# VGND 0.168f $ **FLOATING
C1875 a_4220_14735# VGND 0.259f $ **FLOATING
C1876 a_11219_14887# VGND 0.56f $ **FLOATING
C1877 a_10699_14735# VGND 0.698f $ **FLOATING
C1878 _151_ VGND 0.688f $ **FLOATING
C1879 a_10239_14735# VGND 0.619f $ **FLOATING
C1880 _150_ VGND 1.47f $ **FLOATING
C1881 _156_ VGND 4.45f $ **FLOATING
C1882 a_9647_14709# VGND 0.729f $ **FLOATING
C1883 a_9167_14763# VGND 0.56f $ **FLOATING
C1884 a_6364_14985# VGND 0.546f $ **FLOATING
C1885 _160_ VGND 1.01f $ **FLOATING
C1886 _159_ VGND 0.945f $ **FLOATING
C1887 _157_ VGND 5.29f $ **FLOATING
C1888 a_4880_14735# VGND 0.736f $ **FLOATING
C1889 a_5055_14709# VGND 1.13f $ **FLOATING
C1890 a_4315_14735# VGND 0.714f $ **FLOATING
C1891 _044_ VGND 1.66f $ **FLOATING
C1892 a_4533_14977# VGND 0.653f $ **FLOATING
C1893 a_3965_14735# VGND 1.57f $ **FLOATING
C1894 _003_ VGND 1.26f $ **FLOATING
C1895 a_3799_14735# VGND 1.92f $ **FLOATING
C1896 net36 VGND 14.4f $ **FLOATING
C1897 a_22455_15279# VGND 0.168f $ **FLOATING
C1898 a_19973_15279# VGND 0.219f $ **FLOATING
C1899 a_11343_15279# VGND 0.238f $ **FLOATING
C1900 a_22252_15645# VGND 0.259f $ **FLOATING
C1901 _011_ VGND 1.25f $ **FLOATING
C1902 a_8912_15599# VGND 0.205f $ **FLOATING
C1903 a_7275_15279# VGND 0.168f $ **FLOATING
C1904 a_7072_15645# VGND 0.259f $ **FLOATING
C1905 a_23671_15287# VGND 0.648f $ **FLOATING
C1906 net37 VGND 15.7f $ **FLOATING
C1907 a_22912_15657# VGND 0.736f $ **FLOATING
C1908 a_23087_15583# VGND 0.971f $ **FLOATING
C1909 a_22347_15657# VGND 0.714f $ **FLOATING
C1910 a_22565_15253# VGND 0.653f $ **FLOATING
C1911 a_21997_15285# VGND 1.57f $ **FLOATING
C1912 _009_ VGND 1.22f $ **FLOATING
C1913 a_21831_15285# VGND 1.92f $ **FLOATING
C1914 _144_ VGND 0.832f $ **FLOATING
C1915 _141_ VGND 1.31f $ **FLOATING
C1916 tdc0.r_ring_ctr[3] VGND 3.77f $ **FLOATING
C1917 _142_ VGND 0.846f $ **FLOATING
C1918 a_20503_15253# VGND 0.698f $ **FLOATING
C1919 a_19723_15279# VGND 0.684f $ **FLOATING
C1920 _147_ VGND 0.744f $ **FLOATING
C1921 tdc0.r_ring_ctr[5] VGND 2.87f $ **FLOATING
C1922 a_10363_15617# VGND 0.56f $ **FLOATING
C1923 _145_ VGND 3.04f $ **FLOATING
C1924 a_9551_15511# VGND 0.619f $ **FLOATING
C1925 tdc0.r_ring_ctr[7] VGND 2.66f $ **FLOATING
C1926 a_8686_15395# VGND 0.443f $ **FLOATING
C1927 a_8543_15253# VGND 0.65f $ **FLOATING
C1928 a_7732_15657# VGND 0.736f $ **FLOATING
C1929 a_7907_15583# VGND 0.971f $ **FLOATING
C1930 a_7167_15657# VGND 0.714f $ **FLOATING
C1931 _039_ VGND 1.69f $ **FLOATING
C1932 a_7385_15253# VGND 0.653f $ **FLOATING
C1933 a_6817_15285# VGND 1.57f $ **FLOATING
C1934 _013_ VGND 1.49f $ **FLOATING
C1935 a_6651_15285# VGND 1.92f $ **FLOATING
C1936 _035_ VGND 1.61f $ **FLOATING
C1937 tdc0.r_ring_ctr[1] VGND 5.55f $ **FLOATING
C1938 a_21259_16189# VGND 0.168f $ **FLOATING
C1939 a_21056_15823# VGND 0.259f $ **FLOATING
C1940 a_21716_15823# VGND 0.736f $ **FLOATING
C1941 a_21891_15797# VGND 0.971f $ **FLOATING
C1942 a_21151_15823# VGND 0.714f $ **FLOATING
C1943 a_21369_16065# VGND 0.653f $ **FLOATING
C1944 a_20801_15823# VGND 1.57f $ **FLOATING
C1945 _007_ VGND 1.52f $ **FLOATING
C1946 a_20635_15823# VGND 1.92f $ **FLOATING
C1947 tdc0.r_ring_ctr[0] VGND 5.76f $ **FLOATING
C1948 a_19327_16189# VGND 0.168f $ **FLOATING
C1949 a_19124_15823# VGND 0.259f $ **FLOATING
C1950 a_19784_15823# VGND 0.736f $ **FLOATING
C1951 a_19959_15797# VGND 1.13f $ **FLOATING
C1952 a_19219_15823# VGND 0.714f $ **FLOATING
C1953 _032_ VGND 1.73f $ **FLOATING
C1954 a_19437_16065# VGND 0.653f $ **FLOATING
C1955 a_18869_15823# VGND 1.57f $ **FLOATING
C1956 _000_ VGND 1.37f $ **FLOATING
C1957 a_18703_15823# VGND 1.92f $ **FLOATING
C1958 a_15925_15823# VGND 0.211f $ **FLOATING
C1959 a_16935_16189# VGND 0.168f $ **FLOATING
C1960 a_16732_15823# VGND 0.259f $ **FLOATING
C1961 a_17392_15823# VGND 0.736f $ **FLOATING
C1962 a_17567_15797# VGND 0.971f $ **FLOATING
C1963 a_16827_15823# VGND 0.714f $ **FLOATING
C1964 _041_ VGND 1.6f $ **FLOATING
C1965 a_17045_16065# VGND 0.653f $ **FLOATING
C1966 a_16477_15823# VGND 1.57f $ **FLOATING
C1967 a_16311_15823# VGND 1.92f $ **FLOATING
C1968 _015_ VGND 1.05f $ **FLOATING
C1969 a_14267_16189# VGND 0.168f $ **FLOATING
C1970 a_14064_15823# VGND 0.259f $ **FLOATING
C1971 a_15687_15823# VGND 0.706f $ **FLOATING
C1972 tdc0.r_ring_ctr[9] VGND 6.91f $ **FLOATING
C1973 _153_ VGND 1.3f $ **FLOATING
C1974 a_14724_15823# VGND 0.736f $ **FLOATING
C1975 a_14899_15797# VGND 1.13f $ **FLOATING
C1976 a_14159_15823# VGND 0.714f $ **FLOATING
C1977 _040_ VGND 1.66f $ **FLOATING
C1978 a_14377_16065# VGND 0.653f $ **FLOATING
C1979 a_13809_15823# VGND 1.57f $ **FLOATING
C1980 a_13643_15823# VGND 1.92f $ **FLOATING
C1981 net10 VGND 9.34f $ **FLOATING
C1982 _014_ VGND 1.15f $ **FLOATING
C1983 a_13073_16073# VGND 0.219f $ **FLOATING
C1984 a_11049_16073# VGND 0.219f $ **FLOATING
C1985 a_12823_16073# VGND 0.684f $ **FLOATING
C1986 tdc0.r_ring_ctr[8] VGND 6.72f $ **FLOATING
C1987 _152_ VGND 7.37f $ **FLOATING
C1988 a_10799_16073# VGND 0.684f $ **FLOATING
C1989 _143_ VGND 9.35f $ **FLOATING
C1990 _146_ VGND 1.7f $ **FLOATING
C1991 a_9690_16189# VGND 0.259f $ **FLOATING
C1992 a_9272_16189# VGND 0.168f $ **FLOATING
C1993 tdc0.r_ring_ctr[6] VGND 4.5f $ **FLOATING
C1994 a_9058_16189# VGND 0.653f $ **FLOATING
C1995 a_9127_16060# VGND 0.714f $ **FLOATING
C1996 a_8971_15965# VGND 1.92f $ **FLOATING
C1997 a_8932_16091# VGND 1.57f $ **FLOATING
C1998 a_8654_16075# VGND 0.736f $ **FLOATING
C1999 a_8451_15797# VGND 0.971f $ **FLOATING
C2000 _033_ VGND 1.69f $ **FLOATING
C2001 tdc0.r_ring_ctr[4] VGND 3.74f $ **FLOATING
C2002 a_11967_16367# VGND 0.168f $ **FLOATING
C2003 a_11764_16733# VGND 0.259f $ **FLOATING
C2004 _012_ VGND 1.15f $ **FLOATING
C2005 _038_ VGND 1.69f $ **FLOATING
C2006 a_18059_16375# VGND 0.648f $ **FLOATING
C2007 tdc0.w_ring_buf[0] VGND 4.71f $ **FLOATING
C2008 a_12424_16745# VGND 0.736f $ **FLOATING
C2009 a_12599_16671# VGND 0.971f $ **FLOATING
C2010 a_11859_16745# VGND 0.714f $ **FLOATING
C2011 _036_ VGND 1.74f $ **FLOATING
C2012 a_12077_16341# VGND 0.653f $ **FLOATING
C2013 a_11509_16373# VGND 1.57f $ **FLOATING
C2014 _010_ VGND 1.28f $ **FLOATING
C2015 a_11343_16373# VGND 1.92f $ **FLOATING
C2016 net9 VGND 16f $ **FLOATING
C2017 _149_ VGND 1.12f $ **FLOATING
C2018 _148_ VGND 1.87f $ **FLOATING
C2019 _195_ VGND 15.8f $ **FLOATING
C2020 tt_um_hpretl_tt06_tdc_v2_91.HI VGND 0.415f $ **FLOATING
C2021 tt_um_hpretl_tt06_tdc_v2_82.HI VGND 0.415f $ **FLOATING
C2022 tt_um_hpretl_tt06_tdc_v2_87.HI VGND 0.415f $ **FLOATING
C2023 tt_um_hpretl_tt06_tdc_v2_83.HI VGND 0.415f $ **FLOATING
C2024 tt_um_hpretl_tt06_tdc_v2_78.HI VGND 0.415f $ **FLOATING
C2025 tt_um_hpretl_tt06_tdc_v2_79.HI VGND 0.415f $ **FLOATING
C2026 tt_um_hpretl_tt06_tdc_v2_80.HI VGND 0.415f $ **FLOATING
C2027 tt_um_hpretl_tt06_tdc_v2_93.HI VGND 0.415f $ **FLOATING
C2028 tt_um_hpretl_tt06_tdc_v2_81.HI VGND 0.415f $ **FLOATING
C2029 tt_um_hpretl_tt06_tdc_v2_89.HI VGND 0.415f $ **FLOATING
C2030 tt_um_hpretl_tt06_tdc_v2_85.HI VGND 0.415f $ **FLOATING
C2031 tt_um_hpretl_tt06_tdc_v2_88.HI VGND 0.415f $ **FLOATING
C2032 tt_um_hpretl_tt06_tdc_v2_86.HI VGND 0.415f $ **FLOATING
.ends
