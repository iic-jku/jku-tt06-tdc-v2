magic
tech sky130A
magscale 1 2
timestamp 1711104299
<< viali >>
rect 13829 18785 13863 18819
rect 13645 18581 13679 18615
rect 17509 13957 17543 13991
rect 19717 13957 19751 13991
rect 15209 13821 15243 13855
rect 17601 13821 17635 13855
rect 17969 13821 18003 13855
rect 18153 13821 18187 13855
rect 18245 13821 18279 13855
rect 18889 13821 18923 13855
rect 19257 13821 19291 13855
rect 19625 13821 19659 13855
rect 20085 13821 20119 13855
rect 18337 13753 18371 13787
rect 18521 13753 18555 13787
rect 15301 13685 15335 13719
rect 18061 13685 18095 13719
rect 18429 13685 18463 13719
rect 19901 13685 19935 13719
rect 16926 13413 16960 13447
rect 18429 13413 18463 13447
rect 20186 13413 20220 13447
rect 15577 13345 15611 13379
rect 18337 13345 18371 13379
rect 18613 13345 18647 13379
rect 14933 13277 14967 13311
rect 16681 13277 16715 13311
rect 18797 13277 18831 13311
rect 20453 13277 20487 13311
rect 15301 13209 15335 13243
rect 15393 13209 15427 13243
rect 15761 13141 15795 13175
rect 18061 13141 18095 13175
rect 19073 13141 19107 13175
rect 19993 12937 20027 12971
rect 21833 12937 21867 12971
rect 15301 12869 15335 12903
rect 16681 12801 16715 12835
rect 13369 12733 13403 12767
rect 13553 12733 13587 12767
rect 14013 12733 14047 12767
rect 14381 12733 14415 12767
rect 14657 12733 14691 12767
rect 16957 12733 16991 12767
rect 20545 12733 20579 12767
rect 14565 12665 14599 12699
rect 16589 12665 16623 12699
rect 18705 12665 18739 12699
rect 13185 12597 13219 12631
rect 13737 12597 13771 12631
rect 13921 12597 13955 12631
rect 18061 12597 18095 12631
rect 18889 12393 18923 12427
rect 20821 12393 20855 12427
rect 21649 12393 21683 12427
rect 22201 12393 22235 12427
rect 12633 12325 12667 12359
rect 17601 12325 17635 12359
rect 21281 12325 21315 12359
rect 21465 12325 21499 12359
rect 21925 12325 21959 12359
rect 10977 12257 11011 12291
rect 11713 12257 11747 12291
rect 11989 12257 12023 12291
rect 12265 12257 12299 12291
rect 12725 12257 12759 12291
rect 13001 12257 13035 12291
rect 13369 12257 13403 12291
rect 13553 12257 13587 12291
rect 15669 12257 15703 12291
rect 15945 12257 15979 12291
rect 19697 12257 19731 12291
rect 20913 12257 20947 12291
rect 19441 12189 19475 12223
rect 12081 12121 12115 12155
rect 12449 12121 12483 12155
rect 21005 12121 21039 12155
rect 11069 12053 11103 12087
rect 11805 12053 11839 12087
rect 12909 12053 12943 12087
rect 13645 12053 13679 12087
rect 14013 12053 14047 12087
rect 14565 12053 14599 12087
rect 21465 12053 21499 12087
rect 11069 11849 11103 11883
rect 11161 11849 11195 11883
rect 11897 11849 11931 11883
rect 12633 11849 12667 11883
rect 13093 11849 13127 11883
rect 14473 11849 14507 11883
rect 16773 11849 16807 11883
rect 10425 11781 10459 11815
rect 13829 11781 13863 11815
rect 16313 11781 16347 11815
rect 12081 11713 12115 11747
rect 16405 11713 16439 11747
rect 18797 11713 18831 11747
rect 18889 11713 18923 11747
rect 24225 11713 24259 11747
rect 10241 11645 10275 11679
rect 10333 11645 10367 11679
rect 10609 11645 10643 11679
rect 10701 11645 10735 11679
rect 10885 11645 10919 11679
rect 11063 11645 11097 11679
rect 11167 11645 11201 11679
rect 11345 11645 11379 11679
rect 11437 11645 11471 11679
rect 11621 11645 11655 11679
rect 11713 11645 11747 11679
rect 11989 11645 12023 11679
rect 12449 11645 12483 11679
rect 12633 11645 12667 11679
rect 12725 11645 12759 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 15761 11645 15795 11679
rect 15853 11645 15887 11679
rect 16037 11645 16071 11679
rect 18245 11645 18279 11679
rect 18337 11645 18371 11679
rect 18705 11645 18739 11679
rect 19073 11645 19107 11679
rect 23949 11645 23983 11679
rect 11529 11577 11563 11611
rect 13185 11577 13219 11611
rect 13369 11577 13403 11611
rect 19349 11577 19383 11611
rect 21097 11577 21131 11611
rect 21189 11577 21223 11611
rect 22937 11577 22971 11611
rect 10149 11509 10183 11543
rect 12357 11509 12391 11543
rect 18429 11509 18463 11543
rect 9597 11305 9631 11339
rect 9873 11305 9907 11339
rect 11437 11305 11471 11339
rect 14289 11305 14323 11339
rect 18981 11305 19015 11339
rect 23489 11305 23523 11339
rect 12725 11237 12759 11271
rect 16129 11237 16163 11271
rect 18889 11237 18923 11271
rect 9505 11169 9539 11203
rect 9689 11169 9723 11203
rect 9781 11169 9815 11203
rect 9965 11169 9999 11203
rect 10057 11169 10091 11203
rect 10333 11169 10367 11203
rect 10609 11169 10643 11203
rect 13369 11169 13403 11203
rect 14197 11169 14231 11203
rect 14821 11169 14855 11203
rect 16221 11169 16255 11203
rect 16957 11169 16991 11203
rect 19349 11169 19383 11203
rect 21281 11169 21315 11203
rect 23213 11169 23247 11203
rect 23673 11169 23707 11203
rect 14565 11101 14599 11135
rect 18705 11101 18739 11135
rect 23029 11101 23063 11135
rect 10701 11033 10735 11067
rect 13185 11033 13219 11067
rect 20637 11033 20671 11067
rect 23765 11033 23799 11067
rect 10149 10965 10183 10999
rect 10425 10965 10459 10999
rect 15945 10965 15979 10999
rect 9689 10761 9723 10795
rect 10425 10761 10459 10795
rect 13645 10761 13679 10795
rect 23397 10761 23431 10795
rect 23581 10761 23615 10795
rect 9413 10693 9447 10727
rect 13369 10625 13403 10659
rect 14473 10625 14507 10659
rect 22017 10625 22051 10659
rect 24225 10625 24259 10659
rect 9321 10557 9355 10591
rect 9413 10557 9447 10591
rect 9573 10557 9607 10591
rect 9689 10557 9723 10591
rect 9873 10557 9907 10591
rect 9965 10557 9999 10591
rect 10057 10557 10091 10591
rect 10241 10557 10275 10591
rect 10425 10557 10459 10591
rect 10517 10557 10551 10591
rect 10793 10557 10827 10591
rect 11253 10557 11287 10591
rect 11345 10557 11379 10591
rect 11529 10557 11563 10591
rect 11897 10557 11931 10591
rect 13553 10557 13587 10591
rect 14657 10557 14691 10591
rect 20545 10557 20579 10591
rect 23489 10557 23523 10591
rect 23857 10557 23891 10591
rect 24317 10557 24351 10591
rect 24409 10557 24443 10591
rect 11437 10489 11471 10523
rect 13102 10489 13136 10523
rect 14933 10489 14967 10523
rect 16773 10489 16807 10523
rect 18705 10489 18739 10523
rect 20453 10489 20487 10523
rect 20812 10489 20846 10523
rect 22284 10489 22318 10523
rect 23949 10489 23983 10523
rect 9229 10421 9263 10455
rect 10609 10421 10643 10455
rect 10885 10421 10919 10455
rect 11161 10421 11195 10455
rect 11713 10421 11747 10455
rect 11989 10421 12023 10455
rect 16221 10421 16255 10455
rect 18061 10421 18095 10455
rect 21925 10421 21959 10455
rect 24501 10421 24535 10455
rect 9321 10217 9355 10251
rect 9597 10217 9631 10251
rect 10149 10217 10183 10251
rect 10701 10217 10735 10251
rect 11253 10217 11287 10251
rect 15485 10217 15519 10251
rect 16497 10217 16531 10251
rect 17141 10217 17175 10251
rect 18981 10217 19015 10251
rect 9873 10149 9907 10183
rect 11529 10149 11563 10183
rect 14105 10149 14139 10183
rect 18429 10149 18463 10183
rect 20269 10149 20303 10183
rect 8953 10081 8987 10115
rect 9137 10081 9171 10115
rect 9229 10081 9263 10115
rect 9413 10081 9447 10115
rect 9505 10081 9539 10115
rect 9689 10081 9723 10115
rect 9781 10081 9815 10115
rect 9965 10081 9999 10115
rect 10057 10081 10091 10115
rect 10241 10081 10275 10115
rect 10333 10081 10367 10115
rect 10425 10081 10459 10115
rect 10609 10081 10643 10115
rect 10793 10081 10827 10115
rect 11161 10081 11195 10115
rect 11345 10081 11379 10115
rect 11437 10081 11471 10115
rect 11889 10079 11923 10113
rect 12265 10081 12299 10115
rect 14197 10081 14231 10115
rect 16221 10081 16255 10115
rect 20453 10081 20487 10115
rect 21097 10081 21131 10115
rect 21281 10081 21315 10115
rect 23121 10081 23155 10115
rect 24961 10081 24995 10115
rect 12357 10013 12391 10047
rect 21005 10013 21039 10047
rect 24869 10013 24903 10047
rect 9137 9945 9171 9979
rect 20729 9945 20763 9979
rect 11805 9877 11839 9911
rect 22753 9877 22787 9911
rect 25053 9877 25087 9911
rect 10241 9673 10275 9707
rect 23213 9673 23247 9707
rect 23857 9673 23891 9707
rect 10793 9605 10827 9639
rect 15577 9605 15611 9639
rect 19165 9605 19199 9639
rect 21005 9605 21039 9639
rect 9597 9469 9631 9503
rect 9873 9469 9907 9503
rect 10149 9469 10183 9503
rect 10609 9469 10643 9503
rect 10701 9469 10735 9503
rect 11069 9469 11103 9503
rect 11161 9469 11195 9503
rect 11529 9469 11563 9503
rect 13645 9469 13679 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 22293 9469 22327 9503
rect 23673 9469 23707 9503
rect 25237 9469 25271 9503
rect 25513 9469 25547 9503
rect 25605 9469 25639 9503
rect 25881 9469 25915 9503
rect 13369 9401 13403 9435
rect 13890 9401 13924 9435
rect 17386 9401 17420 9435
rect 20453 9401 20487 9435
rect 22477 9401 22511 9435
rect 23305 9401 23339 9435
rect 24992 9401 25026 9435
rect 25973 9401 26007 9435
rect 9781 9333 9815 9367
rect 10057 9333 10091 9367
rect 10425 9333 10459 9367
rect 11345 9333 11379 9367
rect 11897 9333 11931 9367
rect 15025 9333 15059 9367
rect 18521 9333 18555 9367
rect 22753 9333 22787 9367
rect 23581 9333 23615 9367
rect 25421 9333 25455 9367
rect 25697 9333 25731 9367
rect 22569 9129 22603 9163
rect 25329 9129 25363 9163
rect 10149 9061 10183 9095
rect 12173 9061 12207 9095
rect 14197 9061 14231 9095
rect 16497 9061 16531 9095
rect 21281 9061 21315 9095
rect 10057 8993 10091 9027
rect 10241 8993 10275 9027
rect 10425 8993 10459 9027
rect 10517 8993 10551 9027
rect 10793 8993 10827 9027
rect 11161 8993 11195 9027
rect 11253 8993 11287 9027
rect 11437 8993 11471 9027
rect 11621 8993 11655 9027
rect 11713 8993 11747 9027
rect 12541 8993 12575 9027
rect 14105 8993 14139 9027
rect 16129 8993 16163 9027
rect 18705 8993 18739 9027
rect 18797 8993 18831 9027
rect 20729 8993 20763 9027
rect 23121 8993 23155 9027
rect 23489 8993 23523 9027
rect 25329 8993 25363 9027
rect 25513 8993 25547 9027
rect 16221 8925 16255 8959
rect 11345 8857 11379 8891
rect 17233 8857 17267 8891
rect 10701 8789 10735 8823
rect 11069 8789 11103 8823
rect 12081 8789 12115 8823
rect 15669 8789 15703 8823
rect 16773 8789 16807 8823
rect 20085 8789 20119 8823
rect 21005 8789 21039 8823
rect 24777 8789 24811 8823
rect 10241 8585 10275 8619
rect 11897 8585 11931 8619
rect 13645 8585 13679 8619
rect 13829 8585 13863 8619
rect 16589 8585 16623 8619
rect 18521 8585 18555 8619
rect 21833 8585 21867 8619
rect 22661 8585 22695 8619
rect 23029 8585 23063 8619
rect 19165 8517 19199 8551
rect 23397 8517 23431 8551
rect 9413 8381 9447 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 11529 8381 11563 8415
rect 13737 8381 13771 8415
rect 15209 8381 15243 8415
rect 17141 8381 17175 8415
rect 20545 8381 20579 8415
rect 23213 8381 23247 8415
rect 23581 8381 23615 8415
rect 23857 8381 23891 8415
rect 25329 8381 25363 8415
rect 25605 8381 25639 8415
rect 9321 8313 9355 8347
rect 13369 8313 13403 8347
rect 14942 8313 14976 8347
rect 15301 8313 15335 8347
rect 17408 8313 17442 8347
rect 20453 8313 20487 8347
rect 22753 8313 22787 8347
rect 24102 8313 24136 8347
rect 9689 8245 9723 8279
rect 25237 8245 25271 8279
rect 25421 8245 25455 8279
rect 25697 8245 25731 8279
rect 10149 8041 10183 8075
rect 13645 8041 13679 8075
rect 15669 8041 15703 8075
rect 16957 8041 16991 8075
rect 18521 8041 18555 8075
rect 20361 8041 20395 8075
rect 22753 8041 22787 8075
rect 23121 7973 23155 8007
rect 10241 7905 10275 7939
rect 10333 7905 10367 7939
rect 10517 7905 10551 7939
rect 10701 7905 10735 7939
rect 10793 7905 10827 7939
rect 11253 7905 11287 7939
rect 11529 7905 11563 7939
rect 11897 7905 11931 7939
rect 11989 7905 12023 7939
rect 12357 7905 12391 7939
rect 14197 7905 14231 7939
rect 16221 7905 16255 7939
rect 17141 7905 17175 7939
rect 17233 7905 17267 7939
rect 19073 7905 19107 7939
rect 20913 7905 20947 7939
rect 21281 7905 21315 7939
rect 11161 7837 11195 7871
rect 11437 7837 11471 7871
rect 11713 7769 11747 7803
rect 10425 7701 10459 7735
rect 12173 7701 12207 7735
rect 16497 7701 16531 7735
rect 21005 7701 21039 7735
rect 24409 7701 24443 7735
rect 15853 7497 15887 7531
rect 19901 7497 19935 7531
rect 20729 7429 20763 7463
rect 23489 7361 23523 7395
rect 13645 7293 13679 7327
rect 14565 7293 14599 7327
rect 16405 7293 16439 7327
rect 18521 7293 18555 7327
rect 20085 7293 20119 7327
rect 11529 7225 11563 7259
rect 11805 7225 11839 7259
rect 13369 7225 13403 7259
rect 14105 7225 14139 7259
rect 18797 7225 18831 7259
rect 19165 7225 19199 7259
rect 19349 7225 19383 7259
rect 19717 7225 19751 7259
rect 22017 7225 22051 7259
rect 23222 7225 23256 7259
rect 10241 7157 10275 7191
rect 13829 7157 13863 7191
rect 14197 7157 14231 7191
rect 17693 7157 17727 7191
rect 22109 7157 22143 7191
rect 13645 6953 13679 6987
rect 17417 6953 17451 6987
rect 22385 6953 22419 6987
rect 23029 6953 23063 6987
rect 22201 6885 22235 6919
rect 11253 6817 11287 6851
rect 11437 6817 11471 6851
rect 11713 6817 11747 6851
rect 12173 6817 12207 6851
rect 12357 6817 12391 6851
rect 14197 6817 14231 6851
rect 16129 6817 16163 6851
rect 17969 6817 18003 6851
rect 18225 6817 18259 6851
rect 19441 6817 19475 6851
rect 19984 6817 20018 6851
rect 21373 6817 21407 6851
rect 21741 6817 21775 6851
rect 22385 6817 22419 6851
rect 22569 6817 22603 6851
rect 22661 6817 22695 6851
rect 23121 6817 23155 6851
rect 11621 6749 11655 6783
rect 19717 6749 19751 6783
rect 11345 6681 11379 6715
rect 19349 6681 19383 6715
rect 21097 6681 21131 6715
rect 12081 6613 12115 6647
rect 15669 6613 15703 6647
rect 19533 6613 19567 6647
rect 21925 6613 21959 6647
rect 22753 6613 22787 6647
rect 11989 6409 12023 6443
rect 17141 6409 17175 6443
rect 18797 6409 18831 6443
rect 21833 6409 21867 6443
rect 22109 6409 22143 6443
rect 14105 6341 14139 6375
rect 17325 6341 17359 6375
rect 22385 6341 22419 6375
rect 13369 6205 13403 6239
rect 15393 6205 15427 6239
rect 15485 6205 15519 6239
rect 15761 6205 15795 6239
rect 17509 6205 17543 6239
rect 17785 6205 17819 6239
rect 18337 6205 18371 6239
rect 18705 6205 18739 6239
rect 19441 6205 19475 6239
rect 19809 6205 19843 6239
rect 21741 6205 21775 6239
rect 22017 6207 22051 6241
rect 22201 6205 22235 6239
rect 22293 6205 22327 6239
rect 13102 6137 13136 6171
rect 16028 6137 16062 6171
rect 19901 6137 19935 6171
rect 15577 6069 15611 6103
rect 17693 6069 17727 6103
rect 18153 6069 18187 6103
rect 19257 6069 19291 6103
rect 19625 6069 19659 6103
rect 21189 6069 21223 6103
rect 12357 5865 12391 5899
rect 12909 5865 12943 5899
rect 19625 5865 19659 5899
rect 19993 5865 20027 5899
rect 21649 5865 21683 5899
rect 15761 5797 15795 5831
rect 17233 5797 17267 5831
rect 18981 5797 19015 5831
rect 12449 5729 12483 5763
rect 12817 5729 12851 5763
rect 13277 5729 13311 5763
rect 13921 5729 13955 5763
rect 16221 5729 16255 5763
rect 16681 5729 16715 5763
rect 19073 5729 19107 5763
rect 19165 5729 19199 5763
rect 19349 5729 19383 5763
rect 19533 5729 19567 5763
rect 19625 5729 19659 5763
rect 19809 5729 19843 5763
rect 20085 5729 20119 5763
rect 20177 5729 20211 5763
rect 20637 5729 20671 5763
rect 20729 5729 20763 5763
rect 20821 5729 20855 5763
rect 21465 5729 21499 5763
rect 21741 5729 21775 5763
rect 13369 5661 13403 5695
rect 19441 5661 19475 5695
rect 21373 5593 21407 5627
rect 13737 5525 13771 5559
rect 14473 5525 14507 5559
rect 16313 5525 16347 5559
rect 16865 5525 16899 5559
rect 20269 5525 20303 5559
rect 20545 5525 20579 5559
rect 14105 5321 14139 5355
rect 16129 5321 16163 5355
rect 16589 5321 16623 5355
rect 18061 5321 18095 5355
rect 18337 5321 18371 5355
rect 18981 5321 19015 5355
rect 22017 5321 22051 5355
rect 15945 5253 15979 5287
rect 14565 5185 14599 5219
rect 17785 5185 17819 5219
rect 14197 5117 14231 5151
rect 14473 5117 14507 5151
rect 14821 5117 14855 5151
rect 16037 5117 16071 5151
rect 16497 5117 16531 5151
rect 16681 5117 16715 5151
rect 17601 5117 17635 5151
rect 17693 5117 17727 5151
rect 17969 5117 18003 5151
rect 18153 5117 18187 5151
rect 18429 5117 18463 5151
rect 20453 5117 20487 5151
rect 20545 5117 20579 5151
rect 17509 5049 17543 5083
rect 14381 4981 14415 5015
rect 15485 4777 15519 4811
rect 18061 4777 18095 4811
rect 18705 4777 18739 4811
rect 14105 4641 14139 4675
rect 14372 4641 14406 4675
rect 18153 4641 18187 4675
rect 18521 4641 18555 4675
rect 18705 4641 18739 4675
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 13538 18912 13544 18964
rect 13596 18912 13602 18964
rect 13556 18816 13584 18912
rect 13817 18819 13875 18825
rect 13817 18816 13829 18819
rect 13556 18788 13829 18816
rect 13817 18785 13829 18788
rect 13863 18785 13875 18819
rect 13817 18779 13875 18785
rect 13446 18572 13452 18624
rect 13504 18612 13510 18624
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 13504 18584 13645 18612
rect 13504 18572 13510 18584
rect 13633 18581 13645 18584
rect 13679 18581 13691 18615
rect 13633 18575 13691 18581
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 18690 15988 18696 16040
rect 18748 16028 18754 16040
rect 20806 16028 20812 16040
rect 18748 16000 20812 16028
rect 18748 15988 18754 16000
rect 20806 15988 20812 16000
rect 20864 15988 20870 16040
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 19978 15376 19984 15428
rect 20036 15416 20042 15428
rect 22186 15416 22192 15428
rect 20036 15388 22192 15416
rect 20036 15376 20042 15388
rect 22186 15376 22192 15388
rect 22244 15376 22250 15428
rect 20622 15308 20628 15360
rect 20680 15348 20686 15360
rect 24210 15348 24216 15360
rect 20680 15320 24216 15348
rect 20680 15308 20686 15320
rect 24210 15308 24216 15320
rect 24268 15308 24274 15360
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 23842 14328 23848 14340
rect 22066 14300 23848 14328
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 22066 14260 22094 14300
rect 23842 14288 23848 14300
rect 23900 14288 23906 14340
rect 18196 14232 22094 14260
rect 18196 14220 18202 14232
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 17420 14028 19656 14056
rect 15194 13812 15200 13864
rect 15252 13812 15258 13864
rect 17420 13852 17448 14028
rect 17497 13991 17555 13997
rect 17497 13957 17509 13991
rect 17543 13988 17555 13991
rect 18414 13988 18420 14000
rect 17543 13960 18420 13988
rect 17543 13957 17555 13960
rect 17497 13951 17555 13957
rect 18414 13948 18420 13960
rect 18472 13948 18478 14000
rect 19518 13920 19524 13932
rect 18064 13892 19524 13920
rect 17589 13855 17647 13861
rect 17589 13852 17601 13855
rect 17420 13824 17601 13852
rect 17589 13821 17601 13824
rect 17635 13821 17647 13855
rect 17589 13815 17647 13821
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18064 13852 18092 13892
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 18003 13824 18092 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18138 13812 18144 13864
rect 18196 13812 18202 13864
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18233 13815 18291 13821
rect 18340 13824 18889 13852
rect 18248 13784 18276 13815
rect 18340 13796 18368 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19334 13852 19340 13864
rect 19291 13824 19340 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19628 13861 19656 14028
rect 19705 13991 19763 13997
rect 19705 13957 19717 13991
rect 19751 13988 19763 13991
rect 20714 13988 20720 14000
rect 19751 13960 20720 13988
rect 19751 13957 19763 13960
rect 19705 13951 19763 13957
rect 20714 13948 20720 13960
rect 20772 13948 20778 14000
rect 21450 13920 21456 13932
rect 19700 13892 21456 13920
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19444 13824 19625 13852
rect 19444 13796 19472 13824
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 18156 13756 18276 13784
rect 18156 13728 18184 13756
rect 18322 13744 18328 13796
rect 18380 13744 18386 13796
rect 18509 13787 18567 13793
rect 18509 13753 18521 13787
rect 18555 13784 18567 13787
rect 18598 13784 18604 13796
rect 18555 13756 18604 13784
rect 18555 13753 18567 13756
rect 18509 13747 18567 13753
rect 18598 13744 18604 13756
rect 18656 13744 18662 13796
rect 19426 13744 19432 13796
rect 19484 13744 19490 13796
rect 15286 13676 15292 13728
rect 15344 13676 15350 13728
rect 18046 13676 18052 13728
rect 18104 13676 18110 13728
rect 18138 13676 18144 13728
rect 18196 13676 18202 13728
rect 18417 13719 18475 13725
rect 18417 13685 18429 13719
rect 18463 13716 18475 13719
rect 19700 13716 19728 13892
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 21634 13852 21640 13864
rect 20119 13824 21640 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 21634 13812 21640 13824
rect 21692 13812 21698 13864
rect 18463 13688 19728 13716
rect 18463 13685 18475 13688
rect 18417 13679 18475 13685
rect 19886 13676 19892 13728
rect 19944 13676 19950 13728
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 16914 13447 16972 13453
rect 16914 13444 16926 13447
rect 14936 13416 16926 13444
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 14936 13317 14964 13416
rect 16914 13413 16926 13416
rect 16960 13444 16972 13447
rect 18138 13444 18144 13456
rect 16960 13416 18144 13444
rect 16960 13413 16972 13416
rect 16914 13407 16972 13413
rect 18138 13404 18144 13416
rect 18196 13444 18202 13456
rect 18417 13447 18475 13453
rect 18417 13444 18429 13447
rect 18196 13416 18429 13444
rect 18196 13404 18202 13416
rect 18417 13413 18429 13416
rect 18463 13444 18475 13447
rect 18690 13444 18696 13456
rect 18463 13416 18696 13444
rect 18463 13413 18475 13416
rect 18417 13407 18475 13413
rect 18690 13404 18696 13416
rect 18748 13404 18754 13456
rect 19886 13404 19892 13456
rect 19944 13444 19950 13456
rect 20174 13447 20232 13453
rect 20174 13444 20186 13447
rect 19944 13416 20186 13444
rect 19944 13404 19950 13416
rect 20174 13413 20186 13416
rect 20220 13413 20232 13447
rect 20174 13407 20232 13413
rect 15565 13379 15623 13385
rect 15565 13376 15577 13379
rect 15396 13348 15577 13376
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14700 13280 14933 13308
rect 14700 13268 14706 13280
rect 14921 13277 14933 13280
rect 14967 13277 14979 13311
rect 14921 13271 14979 13277
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 15396 13249 15424 13348
rect 15565 13345 15577 13348
rect 15611 13345 15623 13379
rect 18322 13376 18328 13388
rect 15565 13339 15623 13345
rect 17972 13348 18328 13376
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 17972 13252 18000 13348
rect 18322 13336 18328 13348
rect 18380 13336 18386 13388
rect 18598 13336 18604 13388
rect 18656 13336 18662 13388
rect 20622 13376 20628 13388
rect 18800 13348 20628 13376
rect 15381 13243 15439 13249
rect 15381 13209 15393 13243
rect 15427 13209 15439 13243
rect 15381 13203 15439 13209
rect 17954 13200 17960 13252
rect 18012 13200 18018 13252
rect 18616 13240 18644 13336
rect 18800 13317 18828 13348
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13308 20499 13311
rect 20487 13280 21864 13308
rect 20487 13277 20499 13280
rect 20441 13271 20499 13277
rect 18616 13212 19104 13240
rect 15746 13132 15752 13184
rect 15804 13132 15810 13184
rect 18049 13175 18107 13181
rect 18049 13141 18061 13175
rect 18095 13172 18107 13175
rect 18506 13172 18512 13184
rect 18095 13144 18512 13172
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 19076 13181 19104 13212
rect 21836 13184 21864 13280
rect 19061 13175 19119 13181
rect 19061 13141 19073 13175
rect 19107 13172 19119 13175
rect 19242 13172 19248 13184
rect 19107 13144 19248 13172
rect 19107 13141 19119 13144
rect 19061 13135 19119 13141
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 21818 13132 21824 13184
rect 21876 13132 21882 13184
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 19981 12971 20039 12977
rect 19981 12968 19993 12971
rect 19484 12940 19993 12968
rect 19484 12928 19490 12940
rect 19981 12937 19993 12940
rect 20027 12937 20039 12971
rect 19981 12931 20039 12937
rect 21818 12928 21824 12980
rect 21876 12928 21882 12980
rect 15289 12903 15347 12909
rect 15289 12869 15301 12903
rect 15335 12869 15347 12903
rect 15289 12863 15347 12869
rect 14458 12832 14464 12844
rect 14016 12804 14464 12832
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12764 13415 12767
rect 13446 12764 13452 12776
rect 13403 12736 13452 12764
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 14016 12773 14044 12804
rect 14458 12792 14464 12804
rect 14516 12832 14522 12844
rect 15194 12832 15200 12844
rect 14516 12804 15200 12832
rect 14516 12792 14522 12804
rect 14001 12767 14059 12773
rect 14001 12733 14013 12767
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14660 12773 14688 12804
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15304 12832 15332 12863
rect 16206 12832 16212 12844
rect 15304 12804 16212 12832
rect 16206 12792 16212 12804
rect 16264 12832 16270 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16264 12804 16681 12832
rect 16264 12792 16270 12804
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 18874 12832 18880 12844
rect 16669 12795 16727 12801
rect 16868 12804 18880 12832
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14240 12736 14381 12764
rect 14240 12724 14246 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12733 14703 12767
rect 16868 12764 16896 12804
rect 18874 12792 18880 12804
rect 18932 12832 18938 12844
rect 18932 12804 20576 12832
rect 18932 12792 18938 12804
rect 14645 12727 14703 12733
rect 16592 12736 16896 12764
rect 12342 12656 12348 12708
rect 12400 12696 12406 12708
rect 16592 12705 16620 12736
rect 16942 12724 16948 12776
rect 17000 12724 17006 12776
rect 20548 12773 20576 12804
rect 20533 12767 20591 12773
rect 20533 12733 20545 12767
rect 20579 12733 20591 12767
rect 20533 12727 20591 12733
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 12400 12668 14565 12696
rect 12400 12656 12406 12668
rect 14553 12665 14565 12668
rect 14599 12665 14611 12699
rect 14553 12659 14611 12665
rect 16577 12699 16635 12705
rect 16577 12665 16589 12699
rect 16623 12665 16635 12699
rect 16577 12659 16635 12665
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 18693 12699 18751 12705
rect 18693 12696 18705 12699
rect 17736 12668 18705 12696
rect 17736 12656 17742 12668
rect 18693 12665 18705 12668
rect 18739 12665 18751 12699
rect 18693 12659 18751 12665
rect 13170 12588 13176 12640
rect 13228 12588 13234 12640
rect 13725 12631 13783 12637
rect 13725 12597 13737 12631
rect 13771 12628 13783 12631
rect 13814 12628 13820 12640
rect 13771 12600 13820 12628
rect 13771 12597 13783 12600
rect 13725 12591 13783 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 13906 12588 13912 12640
rect 13964 12588 13970 12640
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18049 12631 18107 12637
rect 18049 12628 18061 12631
rect 18012 12600 18061 12628
rect 18012 12588 18018 12600
rect 18049 12597 18061 12600
rect 18095 12597 18107 12631
rect 18049 12591 18107 12597
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 13630 12384 13636 12436
rect 13688 12384 13694 12436
rect 13832 12396 16574 12424
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 12621 12359 12679 12365
rect 12621 12356 12633 12359
rect 11572 12328 12633 12356
rect 11572 12316 11578 12328
rect 12621 12325 12633 12328
rect 12667 12325 12679 12359
rect 12621 12319 12679 12325
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 9640 12260 10977 12288
rect 9640 12248 9646 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11112 12260 11713 12288
rect 11112 12248 11118 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 12434 12288 12440 12300
rect 12299 12260 12440 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11992 12220 12020 12251
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 12710 12248 12716 12300
rect 12768 12248 12774 12300
rect 12989 12291 13047 12297
rect 12989 12257 13001 12291
rect 13035 12257 13047 12291
rect 12989 12251 13047 12257
rect 11296 12192 12020 12220
rect 13004 12220 13032 12251
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 13320 12260 13369 12288
rect 13320 12248 13326 12260
rect 13357 12257 13369 12260
rect 13403 12288 13415 12291
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 13403 12260 13553 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 13541 12257 13553 12260
rect 13587 12288 13599 12291
rect 13648 12288 13676 12384
rect 13832 12368 13860 12396
rect 13814 12316 13820 12368
rect 13872 12316 13878 12368
rect 16546 12356 16574 12396
rect 18874 12384 18880 12436
rect 18932 12384 18938 12436
rect 20809 12427 20867 12433
rect 20809 12393 20821 12427
rect 20855 12424 20867 12427
rect 20855 12396 21588 12424
rect 20855 12393 20867 12396
rect 20809 12387 20867 12393
rect 17589 12359 17647 12365
rect 17589 12356 17601 12359
rect 16546 12328 17601 12356
rect 17589 12325 17601 12328
rect 17635 12325 17647 12359
rect 17589 12319 17647 12325
rect 18782 12316 18788 12368
rect 18840 12356 18846 12368
rect 18840 12328 19840 12356
rect 18840 12316 18846 12328
rect 13587 12260 13676 12288
rect 13587 12257 13599 12260
rect 13541 12251 13599 12257
rect 15654 12248 15660 12300
rect 15712 12248 15718 12300
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16206 12288 16212 12300
rect 15979 12260 16212 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 19058 12248 19064 12300
rect 19116 12288 19122 12300
rect 19685 12291 19743 12297
rect 19685 12288 19697 12291
rect 19116 12260 19697 12288
rect 19116 12248 19122 12260
rect 19685 12257 19697 12260
rect 19731 12257 19743 12291
rect 19812 12288 19840 12328
rect 20714 12316 20720 12368
rect 20772 12356 20778 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 20772 12328 21281 12356
rect 20772 12316 20778 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 21450 12316 21456 12368
rect 21508 12316 21514 12368
rect 21560 12356 21588 12396
rect 21634 12384 21640 12436
rect 21692 12384 21698 12436
rect 22186 12384 22192 12436
rect 22244 12384 22250 12436
rect 21913 12359 21971 12365
rect 21913 12356 21925 12359
rect 21560 12328 21925 12356
rect 21913 12325 21925 12328
rect 21959 12325 21971 12359
rect 21913 12319 21971 12325
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 19812 12260 20913 12288
rect 19685 12251 19743 12257
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 19429 12223 19487 12229
rect 13004 12192 13860 12220
rect 11296 12180 11302 12192
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 12069 12155 12127 12161
rect 12069 12152 12081 12155
rect 11664 12124 12081 12152
rect 11664 12112 11670 12124
rect 12069 12121 12081 12124
rect 12115 12121 12127 12155
rect 12069 12115 12127 12121
rect 12437 12155 12495 12161
rect 12437 12121 12449 12155
rect 12483 12152 12495 12155
rect 12483 12124 13676 12152
rect 12483 12121 12495 12124
rect 12437 12115 12495 12121
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10008 12056 11069 12084
rect 10008 12044 10014 12056
rect 11057 12053 11069 12056
rect 11103 12053 11115 12087
rect 11057 12047 11115 12053
rect 11790 12044 11796 12096
rect 11848 12044 11854 12096
rect 12894 12044 12900 12096
rect 12952 12044 12958 12096
rect 13648 12093 13676 12124
rect 13832 12096 13860 12192
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 13633 12087 13691 12093
rect 13633 12053 13645 12087
rect 13679 12053 13691 12087
rect 13633 12047 13691 12053
rect 13814 12044 13820 12096
rect 13872 12044 13878 12096
rect 13998 12044 14004 12096
rect 14056 12044 14062 12096
rect 14553 12087 14611 12093
rect 14553 12053 14565 12087
rect 14599 12084 14611 12087
rect 14642 12084 14648 12096
rect 14599 12056 14648 12084
rect 14599 12053 14611 12056
rect 14553 12047 14611 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 19444 12084 19472 12183
rect 20530 12112 20536 12164
rect 20588 12152 20594 12164
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 20588 12124 21005 12152
rect 20588 12112 20594 12124
rect 20993 12121 21005 12124
rect 21039 12121 21051 12155
rect 20993 12115 21051 12121
rect 20346 12084 20352 12096
rect 19444 12056 20352 12084
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 20622 12044 20628 12096
rect 20680 12084 20686 12096
rect 21453 12087 21511 12093
rect 21453 12084 21465 12087
rect 20680 12056 21465 12084
rect 20680 12044 20686 12056
rect 21453 12053 21465 12056
rect 21499 12053 21511 12087
rect 21453 12047 21511 12053
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 11054 11840 11060 11892
rect 11112 11840 11118 11892
rect 11149 11883 11207 11889
rect 11149 11849 11161 11883
rect 11195 11880 11207 11883
rect 11238 11880 11244 11892
rect 11195 11852 11244 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11790 11840 11796 11892
rect 11848 11840 11854 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 12434 11880 12440 11892
rect 11931 11852 12440 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 12710 11880 12716 11892
rect 12667 11852 12716 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 13538 11880 13544 11892
rect 13127 11852 13544 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 14458 11880 14464 11892
rect 14148 11852 14464 11880
rect 14148 11840 14154 11852
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16761 11883 16819 11889
rect 16761 11880 16773 11883
rect 15804 11852 16773 11880
rect 15804 11840 15810 11852
rect 16761 11849 16773 11852
rect 16807 11880 16819 11883
rect 17678 11880 17684 11892
rect 16807 11852 17684 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 18690 11840 18696 11892
rect 18748 11840 18754 11892
rect 9674 11772 9680 11824
rect 9732 11812 9738 11824
rect 10413 11815 10471 11821
rect 10413 11812 10425 11815
rect 9732 11784 10425 11812
rect 9732 11772 9738 11784
rect 10413 11781 10425 11784
rect 10459 11781 10471 11815
rect 10413 11775 10471 11781
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 11808 11744 11836 11840
rect 13170 11812 13176 11824
rect 9824 11716 10364 11744
rect 9824 11704 9830 11716
rect 10226 11636 10232 11688
rect 10284 11636 10290 11688
rect 10336 11685 10364 11716
rect 11348 11716 11836 11744
rect 11900 11784 13176 11812
rect 11348 11685 11376 11716
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 10735 11648 10885 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 11051 11679 11109 11685
rect 11051 11645 11063 11679
rect 11097 11678 11109 11679
rect 11155 11679 11213 11685
rect 11155 11678 11167 11679
rect 11097 11650 11167 11678
rect 11097 11645 11109 11650
rect 11051 11639 11109 11645
rect 11155 11645 11167 11650
rect 11201 11676 11213 11679
rect 11333 11679 11391 11685
rect 11201 11648 11284 11676
rect 11201 11645 11213 11648
rect 11155 11639 11213 11645
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10612 11608 10640 11639
rect 9916 11580 10640 11608
rect 11256 11608 11284 11648
rect 11333 11645 11345 11679
rect 11379 11645 11391 11679
rect 11333 11639 11391 11645
rect 11422 11636 11428 11688
rect 11480 11636 11486 11688
rect 11606 11636 11612 11688
rect 11664 11636 11670 11688
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11676 11759 11679
rect 11900 11676 11928 11784
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 13814 11772 13820 11824
rect 13872 11772 13878 11824
rect 14642 11772 14648 11824
rect 14700 11812 14706 11824
rect 16301 11815 16359 11821
rect 14700 11784 15976 11812
rect 14700 11772 14706 11784
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11744 12127 11747
rect 12115 11716 12664 11744
rect 12115 11713 12127 11716
rect 12069 11707 12127 11713
rect 11747 11648 11928 11676
rect 11977 11679 12035 11685
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 11977 11645 11989 11679
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11672 12495 11679
rect 12526 11672 12532 11688
rect 12483 11645 12532 11672
rect 12437 11644 12532 11645
rect 12437 11639 12495 11644
rect 11440 11608 11468 11636
rect 11256 11580 11468 11608
rect 11517 11611 11575 11617
rect 9916 11568 9922 11580
rect 11517 11577 11529 11611
rect 11563 11608 11575 11611
rect 11992 11608 12020 11639
rect 12526 11636 12532 11644
rect 12584 11636 12590 11688
rect 12636 11685 12664 11716
rect 12728 11716 13676 11744
rect 12728 11685 12756 11716
rect 13648 11688 13676 11716
rect 13832 11716 14228 11744
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 12713 11679 12771 11685
rect 12713 11645 12725 11679
rect 12759 11645 12771 11679
rect 12713 11639 12771 11645
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 13630 11636 13636 11688
rect 13688 11636 13694 11688
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 13832 11676 13860 11716
rect 14200 11688 14228 11716
rect 13771 11648 13860 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 13906 11636 13912 11688
rect 13964 11636 13970 11688
rect 14182 11636 14188 11688
rect 14240 11636 14246 11688
rect 15746 11636 15752 11688
rect 15804 11636 15810 11688
rect 15841 11679 15899 11685
rect 15841 11645 15853 11679
rect 15887 11645 15899 11679
rect 15948 11676 15976 11784
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 16942 11812 16948 11824
rect 16347 11784 16948 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 18708 11812 18736 11840
rect 18708 11784 18920 11812
rect 18892 11753 18920 11784
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11744 16451 11747
rect 18785 11747 18843 11753
rect 18785 11744 18797 11747
rect 16439 11716 18797 11744
rect 16439 11713 16451 11716
rect 16393 11707 16451 11713
rect 18785 11713 18797 11716
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11713 18935 11747
rect 18877 11707 18935 11713
rect 24210 11704 24216 11756
rect 24268 11704 24274 11756
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 15948 11648 16037 11676
rect 15841 11639 15899 11645
rect 16025 11645 16037 11648
rect 16071 11645 16083 11679
rect 17954 11676 17960 11688
rect 16025 11639 16083 11645
rect 16546 11648 17960 11676
rect 11563 11580 12020 11608
rect 13173 11611 13231 11617
rect 11563 11577 11575 11580
rect 11517 11571 11575 11577
rect 13173 11577 13185 11611
rect 13219 11608 13231 11611
rect 13262 11608 13268 11620
rect 13219 11580 13268 11608
rect 13219 11577 13231 11580
rect 13173 11571 13231 11577
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 13357 11611 13415 11617
rect 13357 11577 13369 11611
rect 13403 11608 13415 11611
rect 13924 11608 13952 11636
rect 13403 11580 13952 11608
rect 14200 11608 14228 11636
rect 15010 11608 15016 11620
rect 14200 11580 15016 11608
rect 13403 11577 13415 11580
rect 13357 11571 13415 11577
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 15856 11608 15884 11639
rect 16546 11608 16574 11648
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 18104 11648 18245 11676
rect 18104 11636 18110 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 18322 11636 18328 11688
rect 18380 11636 18386 11688
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18472 11648 18705 11676
rect 18472 11636 18478 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 19058 11636 19064 11688
rect 19116 11636 19122 11688
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 22278 11676 22284 11688
rect 19300 11648 22284 11676
rect 19300 11636 19306 11648
rect 22278 11636 22284 11648
rect 22336 11676 22342 11688
rect 23937 11679 23995 11685
rect 23937 11676 23949 11679
rect 22336 11648 23949 11676
rect 22336 11636 22342 11648
rect 23937 11645 23949 11648
rect 23983 11645 23995 11679
rect 23937 11639 23995 11645
rect 15856 11580 16574 11608
rect 17972 11608 18000 11636
rect 19076 11608 19104 11636
rect 17972 11580 19104 11608
rect 19337 11611 19395 11617
rect 19337 11577 19349 11611
rect 19383 11608 19395 11611
rect 19426 11608 19432 11620
rect 19383 11580 19432 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 19426 11568 19432 11580
rect 19484 11568 19490 11620
rect 21082 11568 21088 11620
rect 21140 11568 21146 11620
rect 21174 11568 21180 11620
rect 21232 11568 21238 11620
rect 22925 11611 22983 11617
rect 22925 11577 22937 11611
rect 22971 11608 22983 11611
rect 24026 11608 24032 11620
rect 22971 11580 24032 11608
rect 22971 11577 22983 11580
rect 22925 11571 22983 11577
rect 24026 11568 24032 11580
rect 24084 11568 24090 11620
rect 10134 11500 10140 11552
rect 10192 11500 10198 11552
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 12345 11543 12403 11549
rect 12345 11540 12357 11543
rect 12308 11512 12357 11540
rect 12308 11500 12314 11512
rect 12345 11509 12357 11512
rect 12391 11509 12403 11543
rect 12345 11503 12403 11509
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 14090 11540 14096 11552
rect 12584 11512 14096 11540
rect 12584 11500 12590 11512
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 16666 11540 16672 11552
rect 14608 11512 16672 11540
rect 14608 11500 14614 11512
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 18417 11543 18475 11549
rect 18417 11540 18429 11543
rect 17184 11512 18429 11540
rect 17184 11500 17190 11512
rect 18417 11509 18429 11512
rect 18463 11509 18475 11543
rect 18417 11503 18475 11509
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 9582 11296 9588 11348
rect 9640 11296 9646 11348
rect 9858 11296 9864 11348
rect 9916 11296 9922 11348
rect 10134 11296 10140 11348
rect 10192 11296 10198 11348
rect 11422 11296 11428 11348
rect 11480 11296 11486 11348
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 13538 11336 13544 11348
rect 12308 11308 13544 11336
rect 12308 11296 12314 11308
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 13688 11308 14289 11336
rect 13688 11296 13694 11308
rect 14277 11305 14289 11308
rect 14323 11336 14335 11339
rect 14323 11308 14964 11336
rect 14323 11305 14335 11308
rect 14277 11299 14335 11305
rect 10152 11268 10180 11296
rect 9692 11240 10180 11268
rect 12713 11271 12771 11277
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 9692 11209 9720 11240
rect 12713 11237 12725 11271
rect 12759 11268 12771 11271
rect 14458 11268 14464 11280
rect 12759 11240 14464 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 14936 11268 14964 11308
rect 15010 11296 15016 11348
rect 15068 11336 15074 11348
rect 15068 11308 15608 11336
rect 15068 11296 15074 11308
rect 15580 11268 15608 11308
rect 16390 11296 16396 11348
rect 16448 11336 16454 11348
rect 18322 11336 18328 11348
rect 16448 11308 18328 11336
rect 16448 11296 16454 11308
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 18969 11339 19027 11345
rect 18969 11336 18981 11339
rect 18432 11308 18981 11336
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 14936 11240 15056 11268
rect 15580 11240 16129 11268
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 9456 11172 9505 11200
rect 9456 11160 9462 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 9508 11132 9536 11163
rect 9784 11132 9812 11163
rect 9950 11160 9956 11212
rect 10008 11160 10014 11212
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10410 11200 10416 11212
rect 10367 11172 10416 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 13906 11200 13912 11212
rect 13403 11172 13912 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 9508 11104 9812 11132
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10612 11132 10640 11163
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 14056 11172 14197 11200
rect 14056 11160 14062 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14185 11163 14243 11169
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 14809 11203 14867 11209
rect 14809 11200 14821 11203
rect 14332 11172 14821 11200
rect 14332 11160 14338 11172
rect 14809 11169 14821 11172
rect 14855 11169 14867 11203
rect 15028 11200 15056 11240
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 16117 11231 16175 11237
rect 18138 11228 18144 11280
rect 18196 11268 18202 11280
rect 18432 11268 18460 11308
rect 18969 11305 18981 11308
rect 19015 11305 19027 11339
rect 18969 11299 19027 11305
rect 23477 11339 23535 11345
rect 23477 11305 23489 11339
rect 23523 11336 23535 11339
rect 28258 11336 28264 11348
rect 23523 11308 28264 11336
rect 23523 11305 23535 11308
rect 23477 11299 23535 11305
rect 28258 11296 28264 11308
rect 28316 11296 28322 11348
rect 18196 11240 18460 11268
rect 18196 11228 18202 11240
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 18877 11271 18935 11277
rect 18877 11268 18889 11271
rect 18564 11240 18889 11268
rect 18564 11228 18570 11240
rect 18877 11237 18889 11240
rect 18923 11237 18935 11271
rect 18877 11231 18935 11237
rect 22020 11240 23704 11268
rect 22020 11212 22048 11240
rect 16209 11203 16267 11209
rect 16209 11200 16221 11203
rect 15028 11172 16221 11200
rect 14809 11163 14867 11169
rect 16209 11169 16221 11172
rect 16255 11169 16267 11203
rect 16209 11163 16267 11169
rect 16945 11203 17003 11209
rect 16945 11169 16957 11203
rect 16991 11200 17003 11203
rect 17494 11200 17500 11212
rect 16991 11172 17500 11200
rect 16991 11169 17003 11172
rect 16945 11163 17003 11169
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 19334 11160 19340 11212
rect 19392 11160 19398 11212
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 20640 11172 21281 11200
rect 14366 11132 14372 11144
rect 9916 11104 10640 11132
rect 13188 11104 14372 11132
rect 9916 11092 9922 11104
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 13188 11073 13216 11104
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 14550 11092 14556 11144
rect 14608 11092 14614 11144
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 10689 11067 10747 11073
rect 10689 11064 10701 11067
rect 9732 11036 10701 11064
rect 9732 11024 9738 11036
rect 10689 11033 10701 11036
rect 10735 11033 10747 11067
rect 10689 11027 10747 11033
rect 13173 11067 13231 11073
rect 13173 11033 13185 11067
rect 13219 11033 13231 11067
rect 14568 11064 14596 11092
rect 20640 11073 20668 11172
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 22002 11160 22008 11212
rect 22060 11160 22066 11212
rect 23198 11160 23204 11212
rect 23256 11160 23262 11212
rect 23676 11209 23704 11240
rect 23661 11203 23719 11209
rect 23661 11169 23673 11203
rect 23707 11169 23719 11203
rect 23661 11163 23719 11169
rect 23017 11135 23075 11141
rect 23017 11101 23029 11135
rect 23063 11132 23075 11135
rect 23566 11132 23572 11144
rect 23063 11104 23572 11132
rect 23063 11101 23075 11104
rect 23017 11095 23075 11101
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 13173 11027 13231 11033
rect 13740 11036 14596 11064
rect 20625 11067 20683 11073
rect 10134 10956 10140 11008
rect 10192 10956 10198 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10376 10968 10425 10996
rect 10376 10956 10382 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10413 10959 10471 10965
rect 11330 10956 11336 11008
rect 11388 10996 11394 11008
rect 12894 10996 12900 11008
rect 11388 10968 12900 10996
rect 11388 10956 11394 10968
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 13740 10996 13768 11036
rect 20625 11033 20637 11067
rect 20671 11033 20683 11067
rect 20625 11027 20683 11033
rect 23753 11067 23811 11073
rect 23753 11033 23765 11067
rect 23799 11064 23811 11067
rect 25314 11064 25320 11076
rect 23799 11036 25320 11064
rect 23799 11033 23811 11036
rect 23753 11027 23811 11033
rect 13688 10968 13768 10996
rect 15933 10999 15991 11005
rect 13688 10956 13694 10968
rect 15933 10965 15945 10999
rect 15979 10996 15991 10999
rect 16114 10996 16120 11008
rect 15979 10968 16120 10996
rect 15979 10965 15991 10968
rect 15933 10959 15991 10965
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 20070 10956 20076 11008
rect 20128 10996 20134 11008
rect 20640 10996 20668 11027
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 20128 10968 20668 10996
rect 20128 10956 20134 10968
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 9677 10795 9735 10801
rect 9677 10761 9689 10795
rect 9723 10792 9735 10795
rect 9766 10792 9772 10804
rect 9723 10764 9772 10792
rect 9723 10761 9735 10764
rect 9677 10755 9735 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10284 10764 10425 10792
rect 10284 10752 10290 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 11422 10752 11428 10804
rect 11480 10752 11486 10804
rect 13633 10795 13691 10801
rect 13633 10761 13645 10795
rect 13679 10792 13691 10795
rect 14274 10792 14280 10804
rect 13679 10764 14280 10792
rect 13679 10761 13691 10764
rect 13633 10755 13691 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 20548 10764 22048 10792
rect 9401 10727 9459 10733
rect 9401 10693 9413 10727
rect 9447 10693 9459 10727
rect 11440 10724 11468 10752
rect 9401 10687 9459 10693
rect 10612 10696 11468 10724
rect 9416 10656 9444 10687
rect 10612 10656 10640 10696
rect 14090 10684 14096 10736
rect 14148 10684 14154 10736
rect 9416 10628 9996 10656
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 9582 10597 9588 10600
rect 9561 10591 9588 10597
rect 9561 10557 9573 10591
rect 9561 10551 9588 10557
rect 9582 10548 9588 10551
rect 9640 10548 9646 10600
rect 9968 10597 9996 10628
rect 10428 10628 10640 10656
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10557 9735 10591
rect 9677 10551 9735 10557
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 10091 10560 10241 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 10229 10557 10241 10560
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 9214 10412 9220 10464
rect 9272 10412 9278 10464
rect 9416 10452 9444 10548
rect 9692 10452 9720 10551
rect 9876 10520 9904 10551
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 10428 10597 10456 10628
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 12250 10656 12256 10668
rect 10744 10628 12256 10656
rect 10744 10616 10750 10628
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 10336 10520 10364 10548
rect 9876 10492 10364 10520
rect 9766 10452 9772 10464
rect 9416 10424 9772 10452
rect 9766 10412 9772 10424
rect 9824 10452 9830 10464
rect 10428 10452 10456 10551
rect 10502 10548 10508 10600
rect 10560 10548 10566 10600
rect 10778 10548 10784 10600
rect 10836 10548 10842 10600
rect 11348 10597 11376 10628
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 13630 10656 13636 10668
rect 13403 10628 13636 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10557 11391 10591
rect 11333 10551 11391 10557
rect 11256 10520 11284 10551
rect 11514 10548 11520 10600
rect 11572 10548 11578 10600
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10588 11943 10591
rect 12342 10588 12348 10600
rect 11931 10560 12348 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 14108 10588 14136 10684
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 15378 10656 15384 10668
rect 14507 10628 15384 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 13587 10560 14136 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 14642 10548 14648 10600
rect 14700 10548 14706 10600
rect 14826 10548 14832 10600
rect 14884 10548 14890 10600
rect 20346 10548 20352 10600
rect 20404 10588 20410 10600
rect 20548 10597 20576 10764
rect 22020 10665 22048 10764
rect 23198 10752 23204 10804
rect 23256 10792 23262 10804
rect 23385 10795 23443 10801
rect 23385 10792 23397 10795
rect 23256 10764 23397 10792
rect 23256 10752 23262 10764
rect 23385 10761 23397 10764
rect 23431 10761 23443 10795
rect 23385 10755 23443 10761
rect 23569 10795 23627 10801
rect 23569 10761 23581 10795
rect 23615 10792 23627 10795
rect 23842 10792 23848 10804
rect 23615 10764 23848 10792
rect 23615 10761 23627 10764
rect 23569 10755 23627 10761
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 24026 10684 24032 10736
rect 24084 10724 24090 10736
rect 24084 10696 24440 10724
rect 24084 10684 24090 10696
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 23290 10616 23296 10668
rect 23348 10656 23354 10668
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23348 10628 24225 10656
rect 23348 10616 23354 10628
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 24412 10600 24440 10696
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 20404 10560 20545 10588
rect 20404 10548 20410 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 20533 10551 20591 10557
rect 21082 10548 21088 10600
rect 21140 10588 21146 10600
rect 23477 10591 23535 10597
rect 21928 10588 22094 10590
rect 23477 10588 23489 10591
rect 21140 10562 23489 10588
rect 21140 10560 21956 10562
rect 22066 10560 23489 10562
rect 21140 10548 21146 10560
rect 23477 10557 23489 10560
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 23566 10548 23572 10600
rect 23624 10588 23630 10600
rect 23845 10591 23903 10597
rect 23845 10588 23857 10591
rect 23624 10560 23857 10588
rect 23624 10548 23630 10560
rect 23845 10557 23857 10560
rect 23891 10557 23903 10591
rect 23845 10551 23903 10557
rect 24302 10548 24308 10600
rect 24360 10548 24366 10600
rect 24394 10548 24400 10600
rect 24452 10548 24458 10600
rect 11425 10523 11483 10529
rect 11425 10520 11437 10523
rect 11256 10492 11437 10520
rect 11425 10489 11437 10492
rect 11471 10489 11483 10523
rect 11425 10483 11483 10489
rect 11716 10492 13032 10520
rect 9824 10424 10456 10452
rect 9824 10412 9830 10424
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 10870 10412 10876 10464
rect 10928 10412 10934 10464
rect 11146 10412 11152 10464
rect 11204 10412 11210 10464
rect 11716 10461 11744 10492
rect 11701 10455 11759 10461
rect 11701 10421 11713 10455
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 11977 10455 12035 10461
rect 11977 10421 11989 10455
rect 12023 10452 12035 10455
rect 12342 10452 12348 10464
rect 12023 10424 12348 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12342 10412 12348 10424
rect 12400 10412 12406 10464
rect 13004 10452 13032 10492
rect 13078 10480 13084 10532
rect 13136 10529 13142 10532
rect 13136 10483 13148 10529
rect 13136 10480 13142 10483
rect 14844 10452 14872 10548
rect 14921 10523 14979 10529
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 15654 10520 15660 10532
rect 14967 10492 15660 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 16298 10480 16304 10532
rect 16356 10520 16362 10532
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 16356 10492 16773 10520
rect 16356 10480 16362 10492
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 16761 10483 16819 10489
rect 18414 10480 18420 10532
rect 18472 10520 18478 10532
rect 18693 10523 18751 10529
rect 18693 10520 18705 10523
rect 18472 10492 18705 10520
rect 18472 10480 18478 10492
rect 18693 10489 18705 10492
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 20438 10480 20444 10532
rect 20496 10480 20502 10532
rect 22278 10529 22284 10532
rect 20800 10523 20858 10529
rect 20800 10489 20812 10523
rect 20846 10520 20858 10523
rect 22272 10520 22284 10529
rect 20846 10492 22094 10520
rect 22239 10492 22284 10520
rect 20846 10489 20858 10492
rect 20800 10483 20858 10489
rect 13004 10424 14872 10452
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 16209 10455 16267 10461
rect 16209 10452 16221 10455
rect 15252 10424 16221 10452
rect 15252 10412 15258 10424
rect 16209 10421 16221 10424
rect 16255 10421 16267 10455
rect 16209 10415 16267 10421
rect 16850 10412 16856 10464
rect 16908 10452 16914 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 16908 10424 18061 10452
rect 16908 10412 16914 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 21910 10412 21916 10464
rect 21968 10412 21974 10464
rect 22066 10452 22094 10492
rect 22272 10483 22284 10492
rect 22278 10480 22284 10483
rect 22336 10480 22342 10532
rect 23937 10523 23995 10529
rect 23937 10520 23949 10523
rect 22388 10492 23949 10520
rect 22388 10452 22416 10492
rect 23937 10489 23949 10492
rect 23983 10489 23995 10523
rect 23937 10483 23995 10489
rect 22066 10424 22416 10452
rect 24489 10455 24547 10461
rect 24489 10421 24501 10455
rect 24535 10452 24547 10455
rect 25406 10452 25412 10464
rect 24535 10424 25412 10452
rect 24535 10421 24547 10424
rect 24489 10415 24547 10421
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 9214 10208 9220 10260
rect 9272 10208 9278 10260
rect 9306 10208 9312 10260
rect 9364 10208 9370 10260
rect 9585 10251 9643 10257
rect 9585 10217 9597 10251
rect 9631 10248 9643 10251
rect 10042 10248 10048 10260
rect 9631 10220 10048 10248
rect 9631 10217 9643 10220
rect 9585 10211 9643 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10502 10248 10508 10260
rect 10183 10220 10508 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 10594 10208 10600 10260
rect 10652 10208 10658 10260
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 10778 10248 10784 10260
rect 10735 10220 10784 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 11146 10208 11152 10260
rect 11204 10208 11210 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 13354 10248 13360 10260
rect 11287 10220 13360 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 15378 10248 15384 10260
rect 14516 10220 15384 10248
rect 14516 10208 14522 10220
rect 15378 10208 15384 10220
rect 15436 10248 15442 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 15436 10220 15485 10248
rect 15436 10208 15442 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16758 10248 16764 10260
rect 16531 10220 16764 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 18782 10248 18788 10260
rect 17175 10220 18788 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 18969 10251 19027 10257
rect 18969 10217 18981 10251
rect 19015 10248 19027 10251
rect 24302 10248 24308 10260
rect 19015 10220 24308 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 24302 10208 24308 10220
rect 24360 10208 24366 10260
rect 24394 10208 24400 10260
rect 24452 10208 24458 10260
rect 9232 10180 9260 10208
rect 8956 10152 9260 10180
rect 9324 10152 9812 10180
rect 8956 10121 8984 10152
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10112 9183 10115
rect 9217 10115 9275 10121
rect 9217 10112 9229 10115
rect 9171 10084 9229 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9217 10081 9229 10084
rect 9263 10112 9275 10115
rect 9324 10112 9352 10152
rect 9508 10121 9536 10152
rect 9784 10124 9812 10152
rect 9858 10140 9864 10192
rect 9916 10140 9922 10192
rect 10612 10180 10640 10208
rect 11164 10180 11192 10208
rect 9968 10152 10640 10180
rect 10796 10152 11192 10180
rect 11517 10183 11575 10189
rect 9263 10084 9352 10112
rect 9401 10115 9459 10121
rect 9263 10081 9275 10084
rect 9217 10075 9275 10081
rect 9401 10081 9413 10115
rect 9447 10081 9459 10115
rect 9401 10075 9459 10081
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9416 10044 9444 10075
rect 9674 10072 9680 10124
rect 9732 10072 9738 10124
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 9968 10121 9996 10152
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10081 10011 10115
rect 9953 10075 10011 10081
rect 10042 10072 10048 10124
rect 10100 10072 10106 10124
rect 10134 10072 10140 10124
rect 10192 10072 10198 10124
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10152 10044 10180 10072
rect 9416 10016 10180 10044
rect 10244 10044 10272 10075
rect 10318 10072 10324 10124
rect 10376 10072 10382 10124
rect 10410 10072 10416 10124
rect 10468 10072 10474 10124
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10112 10655 10115
rect 10686 10112 10692 10124
rect 10643 10084 10692 10112
rect 10643 10081 10655 10084
rect 10597 10075 10655 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 10796 10121 10824 10152
rect 11517 10149 11529 10183
rect 11563 10180 11575 10183
rect 12618 10180 12624 10192
rect 11563 10152 12624 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 14093 10183 14151 10189
rect 14093 10149 14105 10183
rect 14139 10180 14151 10183
rect 16298 10180 16304 10192
rect 14139 10152 16304 10180
rect 14139 10149 14151 10152
rect 14093 10143 14151 10149
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 18417 10183 18475 10189
rect 18417 10149 18429 10183
rect 18463 10180 18475 10183
rect 20070 10180 20076 10192
rect 18463 10152 20076 10180
rect 18463 10149 18475 10152
rect 18417 10143 18475 10149
rect 20070 10140 20076 10152
rect 20128 10140 20134 10192
rect 20257 10183 20315 10189
rect 20257 10149 20269 10183
rect 20303 10180 20315 10183
rect 20303 10152 21404 10180
rect 20303 10149 20315 10152
rect 20257 10143 20315 10149
rect 21376 10124 21404 10152
rect 21910 10140 21916 10192
rect 21968 10180 21974 10192
rect 22186 10180 22192 10192
rect 21968 10152 22192 10180
rect 21968 10140 21974 10152
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 10870 10072 10876 10124
rect 10928 10072 10934 10124
rect 11146 10072 11152 10124
rect 11204 10072 11210 10124
rect 11330 10072 11336 10124
rect 11388 10072 11394 10124
rect 11422 10072 11428 10124
rect 11480 10072 11486 10124
rect 11877 10118 11935 10119
rect 11808 10113 11935 10118
rect 11808 10112 11889 10113
rect 11716 10090 11889 10112
rect 11716 10084 11836 10090
rect 10888 10044 10916 10072
rect 10244 10016 10916 10044
rect 11716 9988 11744 10084
rect 11877 10079 11889 10090
rect 11923 10079 11935 10113
rect 11877 10073 11935 10079
rect 12250 10072 12256 10124
rect 12308 10072 12314 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 13872 10084 14197 10112
rect 13872 10072 13878 10084
rect 14185 10081 14197 10084
rect 14231 10081 14243 10115
rect 14185 10075 14243 10081
rect 16206 10072 16212 10124
rect 16264 10072 16270 10124
rect 19518 10072 19524 10124
rect 19576 10072 19582 10124
rect 20162 10072 20168 10124
rect 20220 10112 20226 10124
rect 20441 10115 20499 10121
rect 20441 10112 20453 10115
rect 20220 10084 20453 10112
rect 20220 10072 20226 10084
rect 20441 10081 20453 10084
rect 20487 10081 20499 10115
rect 20441 10075 20499 10081
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 21085 10115 21143 10121
rect 21085 10112 21097 10115
rect 20772 10084 21097 10112
rect 20772 10072 20778 10084
rect 21085 10081 21097 10084
rect 21131 10081 21143 10115
rect 21085 10075 21143 10081
rect 21266 10072 21272 10124
rect 21324 10072 21330 10124
rect 21358 10072 21364 10124
rect 21416 10112 21422 10124
rect 23109 10115 23167 10121
rect 23109 10112 23121 10115
rect 21416 10084 23121 10112
rect 21416 10072 21422 10084
rect 23109 10081 23121 10084
rect 23155 10081 23167 10115
rect 24412 10112 24440 10208
rect 24949 10115 25007 10121
rect 24949 10112 24961 10115
rect 24412 10084 24961 10112
rect 23109 10075 23167 10081
rect 24949 10081 24961 10084
rect 24995 10081 25007 10115
rect 24949 10075 25007 10081
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 19536 10044 19564 10072
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 19536 10016 21005 10044
rect 12345 10007 12403 10013
rect 20993 10013 21005 10016
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 24857 10047 24915 10053
rect 24857 10013 24869 10047
rect 24903 10044 24915 10047
rect 25682 10044 25688 10056
rect 24903 10016 25688 10044
rect 24903 10013 24915 10016
rect 24857 10007 24915 10013
rect 9125 9979 9183 9985
rect 9125 9945 9137 9979
rect 9171 9976 9183 9979
rect 10226 9976 10232 9988
rect 9171 9948 10232 9976
rect 9171 9945 9183 9948
rect 9125 9939 9183 9945
rect 10226 9936 10232 9948
rect 10284 9936 10290 9988
rect 10686 9936 10692 9988
rect 10744 9936 10750 9988
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 12360 9976 12388 10007
rect 25682 10004 25688 10016
rect 25740 10004 25746 10056
rect 11756 9948 12388 9976
rect 20717 9979 20775 9985
rect 11756 9936 11762 9948
rect 20717 9945 20729 9979
rect 20763 9976 20775 9979
rect 20806 9976 20812 9988
rect 20763 9948 20812 9976
rect 20763 9945 20775 9948
rect 20717 9939 20775 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 24302 9936 24308 9988
rect 24360 9976 24366 9988
rect 25590 9976 25596 9988
rect 24360 9948 25596 9976
rect 24360 9936 24366 9948
rect 25590 9936 25596 9948
rect 25648 9936 25654 9988
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 10704 9908 10732 9936
rect 10100 9880 10732 9908
rect 10100 9868 10106 9880
rect 11790 9868 11796 9920
rect 11848 9868 11854 9920
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 14918 9908 14924 9920
rect 12952 9880 14924 9908
rect 12952 9868 12958 9880
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 22738 9868 22744 9920
rect 22796 9868 22802 9920
rect 23934 9868 23940 9920
rect 23992 9908 23998 9920
rect 25041 9911 25099 9917
rect 25041 9908 25053 9911
rect 23992 9880 25053 9908
rect 23992 9868 23998 9880
rect 25041 9877 25053 9880
rect 25087 9877 25099 9911
rect 25041 9871 25099 9877
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 9692 9676 9904 9704
rect 9692 9636 9720 9676
rect 9876 9648 9904 9676
rect 10226 9664 10232 9716
rect 10284 9664 10290 9716
rect 11146 9664 11152 9716
rect 11204 9664 11210 9716
rect 13814 9704 13820 9716
rect 13648 9676 13820 9704
rect 9600 9608 9720 9636
rect 9600 9509 9628 9608
rect 9858 9596 9864 9648
rect 9916 9596 9922 9648
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 11164 9636 11192 9664
rect 10827 9608 11192 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 13648 9636 13676 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 21358 9664 21364 9716
rect 21416 9664 21422 9716
rect 23198 9664 23204 9716
rect 23256 9664 23262 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23584 9676 23857 9704
rect 11296 9608 13676 9636
rect 15565 9639 15623 9645
rect 11296 9596 11302 9608
rect 15565 9605 15577 9639
rect 15611 9636 15623 9639
rect 16390 9636 16396 9648
rect 15611 9608 16396 9636
rect 15611 9605 15623 9608
rect 15565 9599 15623 9605
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 19153 9639 19211 9645
rect 19153 9605 19165 9639
rect 19199 9636 19211 9639
rect 19426 9636 19432 9648
rect 19199 9608 19432 9636
rect 19199 9605 19211 9608
rect 19153 9599 19211 9605
rect 11698 9568 11704 9580
rect 9876 9540 10364 9568
rect 9876 9509 9904 9540
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 10137 9503 10195 9509
rect 10137 9500 10149 9503
rect 10100 9472 10149 9500
rect 10100 9460 10106 9472
rect 10137 9469 10149 9472
rect 10183 9469 10195 9503
rect 10336 9502 10364 9540
rect 11440 9540 11704 9568
rect 10410 9502 10416 9512
rect 10336 9474 10416 9502
rect 10137 9463 10195 9469
rect 10410 9460 10416 9474
rect 10468 9460 10474 9512
rect 10594 9460 10600 9512
rect 10652 9460 10658 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10962 9500 10968 9512
rect 10744 9472 10968 9500
rect 10744 9460 10750 9472
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 11054 9460 11060 9512
rect 11112 9460 11118 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11440 9500 11468 9540
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 16868 9540 17264 9568
rect 11195 9472 11468 9500
rect 11517 9503 11575 9509
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11517 9469 11529 9503
rect 11563 9500 11575 9503
rect 11790 9500 11796 9512
rect 11563 9472 11796 9500
rect 11563 9469 11575 9472
rect 11517 9463 11575 9469
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 13630 9500 13636 9512
rect 12584 9472 13636 9500
rect 12584 9460 12590 9472
rect 13630 9460 13636 9472
rect 13688 9500 13694 9512
rect 15102 9500 15108 9512
rect 13688 9472 15108 9500
rect 13688 9460 13694 9472
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 16868 9509 16896 9540
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9469 17187 9503
rect 17236 9500 17264 9540
rect 19168 9500 19196 9599
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 20993 9639 21051 9645
rect 20993 9605 21005 9639
rect 21039 9636 21051 9639
rect 21376 9636 21404 9664
rect 21039 9608 21404 9636
rect 21039 9605 21051 9608
rect 20993 9599 21051 9605
rect 23474 9596 23480 9648
rect 23532 9636 23538 9648
rect 23584 9636 23612 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 24320 9676 25544 9704
rect 24320 9636 24348 9676
rect 23532 9608 23612 9636
rect 23676 9608 24348 9636
rect 23532 9596 23538 9608
rect 23676 9568 23704 9608
rect 22066 9540 23704 9568
rect 22066 9512 22094 9540
rect 20346 9500 20352 9512
rect 17236 9472 19196 9500
rect 19306 9472 20352 9500
rect 17129 9463 17187 9469
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 13357 9435 13415 9441
rect 13357 9432 13369 9435
rect 13320 9404 13369 9432
rect 13320 9392 13326 9404
rect 13357 9401 13369 9404
rect 13403 9401 13415 9435
rect 13357 9395 13415 9401
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 13878 9435 13936 9441
rect 13878 9432 13890 9435
rect 13780 9404 13890 9432
rect 13780 9392 13786 9404
rect 13878 9401 13890 9404
rect 13924 9401 13936 9435
rect 13878 9395 13936 9401
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 10045 9367 10103 9373
rect 10045 9333 10057 9367
rect 10091 9364 10103 9367
rect 10134 9364 10140 9376
rect 10091 9336 10140 9364
rect 10091 9333 10103 9336
rect 10045 9327 10103 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10410 9324 10416 9376
rect 10468 9324 10474 9376
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 10560 9336 11345 9364
rect 10560 9324 10566 9336
rect 11333 9333 11345 9336
rect 11379 9333 11391 9367
rect 11333 9327 11391 9333
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11848 9336 11897 9364
rect 11848 9324 11854 9336
rect 11885 9333 11897 9336
rect 11931 9333 11943 9367
rect 11885 9327 11943 9333
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 16206 9364 16212 9376
rect 15059 9336 16212 9364
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 17144 9364 17172 9463
rect 17218 9392 17224 9444
rect 17276 9432 17282 9444
rect 17374 9435 17432 9441
rect 17374 9432 17386 9435
rect 17276 9404 17386 9432
rect 17276 9392 17282 9404
rect 17374 9401 17386 9404
rect 17420 9401 17432 9435
rect 18598 9432 18604 9444
rect 17374 9395 17432 9401
rect 17512 9404 18604 9432
rect 17512 9364 17540 9404
rect 18598 9392 18604 9404
rect 18656 9432 18662 9444
rect 19306 9432 19334 9472
rect 20346 9460 20352 9472
rect 20404 9460 20410 9512
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 22002 9500 22008 9512
rect 20772 9472 22008 9500
rect 20772 9460 20778 9472
rect 22002 9460 22008 9472
rect 22060 9472 22094 9512
rect 22060 9460 22066 9472
rect 22186 9460 22192 9512
rect 22244 9460 22250 9512
rect 23676 9509 23704 9540
rect 25516 9512 25544 9676
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9500 22339 9503
rect 23661 9503 23719 9509
rect 22327 9472 23612 9500
rect 22327 9469 22339 9472
rect 22281 9463 22339 9469
rect 18656 9404 19334 9432
rect 18656 9392 18662 9404
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 20036 9404 20453 9432
rect 20036 9392 20042 9404
rect 20441 9401 20453 9404
rect 20487 9401 20499 9435
rect 22204 9432 22232 9460
rect 22465 9435 22523 9441
rect 22465 9432 22477 9435
rect 22204 9404 22477 9432
rect 20441 9395 20499 9401
rect 22465 9401 22477 9404
rect 22511 9401 22523 9435
rect 22465 9395 22523 9401
rect 23293 9435 23351 9441
rect 23293 9401 23305 9435
rect 23339 9432 23351 9435
rect 23474 9432 23480 9444
rect 23339 9404 23480 9432
rect 23339 9401 23351 9404
rect 23293 9395 23351 9401
rect 23474 9392 23480 9404
rect 23532 9392 23538 9444
rect 23584 9432 23612 9472
rect 23661 9469 23673 9503
rect 23707 9469 23719 9503
rect 23661 9463 23719 9469
rect 24026 9460 24032 9512
rect 24084 9500 24090 9512
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 24084 9472 25237 9500
rect 24084 9460 24090 9472
rect 25225 9469 25237 9472
rect 25271 9469 25283 9503
rect 25225 9463 25283 9469
rect 25498 9460 25504 9512
rect 25556 9460 25562 9512
rect 25590 9460 25596 9512
rect 25648 9460 25654 9512
rect 25682 9460 25688 9512
rect 25740 9500 25746 9512
rect 25869 9503 25927 9509
rect 25869 9500 25881 9503
rect 25740 9472 25881 9500
rect 25740 9460 25746 9472
rect 25869 9469 25881 9472
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 24854 9432 24860 9444
rect 23584 9404 24860 9432
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 24980 9435 25038 9441
rect 24980 9401 24992 9435
rect 25026 9432 25038 9435
rect 25961 9435 26019 9441
rect 25961 9432 25973 9435
rect 25026 9404 25973 9432
rect 25026 9401 25038 9404
rect 24980 9395 25038 9401
rect 25961 9401 25973 9404
rect 26007 9401 26019 9435
rect 25961 9395 26019 9401
rect 17144 9336 17540 9364
rect 18509 9367 18567 9373
rect 18509 9333 18521 9367
rect 18555 9364 18567 9367
rect 20162 9364 20168 9376
rect 18555 9336 20168 9364
rect 18555 9333 18567 9336
rect 18509 9327 18567 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 22741 9367 22799 9373
rect 22741 9333 22753 9367
rect 22787 9364 22799 9367
rect 22830 9364 22836 9376
rect 22787 9336 22836 9364
rect 22787 9333 22799 9336
rect 22741 9327 22799 9333
rect 22830 9324 22836 9336
rect 22888 9324 22894 9376
rect 23569 9367 23627 9373
rect 23569 9333 23581 9367
rect 23615 9364 23627 9367
rect 23750 9364 23756 9376
rect 23615 9336 23756 9364
rect 23615 9333 23627 9336
rect 23569 9327 23627 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 25130 9324 25136 9376
rect 25188 9364 25194 9376
rect 25409 9367 25467 9373
rect 25409 9364 25421 9367
rect 25188 9336 25421 9364
rect 25188 9324 25194 9336
rect 25409 9333 25421 9336
rect 25455 9333 25467 9367
rect 25409 9327 25467 9333
rect 25682 9324 25688 9376
rect 25740 9324 25746 9376
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10594 9160 10600 9172
rect 9824 9132 10600 9160
rect 9824 9120 9830 9132
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 11054 9120 11060 9172
rect 11112 9120 11118 9172
rect 15194 9160 15200 9172
rect 11808 9132 15200 9160
rect 10137 9095 10195 9101
rect 10137 9061 10149 9095
rect 10183 9092 10195 9095
rect 11072 9092 11100 9120
rect 10183 9064 11008 9092
rect 11072 9064 11284 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 9024 10287 9027
rect 10413 9027 10471 9033
rect 10413 9024 10425 9027
rect 10275 8996 10425 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 10413 8993 10425 8996
rect 10459 8993 10471 9027
rect 10413 8987 10471 8993
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 8993 10839 9027
rect 10980 9024 11008 9064
rect 11054 9024 11060 9036
rect 10980 8996 11060 9024
rect 10781 8987 10839 8993
rect 10520 8888 10548 8987
rect 10796 8956 10824 8987
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11256 9033 11284 9064
rect 11348 9064 11744 9092
rect 11348 9036 11376 9064
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 11241 9027 11299 9033
rect 11241 8993 11253 9027
rect 11287 8993 11299 9027
rect 11241 8987 11299 8993
rect 10962 8956 10968 8968
rect 10796 8928 10968 8956
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11164 8956 11192 8987
rect 11330 8984 11336 9036
rect 11388 8984 11394 9036
rect 11716 9033 11744 9064
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11471 8996 11621 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 11808 8956 11836 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 16264 9132 16528 9160
rect 16264 9120 16270 9132
rect 12161 9095 12219 9101
rect 12161 9061 12173 9095
rect 12207 9092 12219 9095
rect 12250 9092 12256 9104
rect 12207 9064 12256 9092
rect 12207 9061 12219 9064
rect 12161 9055 12219 9061
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 14185 9095 14243 9101
rect 14185 9092 14197 9095
rect 12406 9064 14197 9092
rect 11164 8928 11836 8956
rect 11238 8888 11244 8900
rect 10520 8860 11244 8888
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 11333 8891 11391 8897
rect 11333 8857 11345 8891
rect 11379 8888 11391 8891
rect 12406 8888 12434 9064
rect 14185 9061 14197 9064
rect 14231 9061 14243 9095
rect 16390 9092 16396 9104
rect 14185 9055 14243 9061
rect 16132 9064 16396 9092
rect 12526 8984 12532 9036
rect 12584 8984 12590 9036
rect 16132 9033 16160 9064
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 16500 9101 16528 9132
rect 17218 9120 17224 9172
rect 17276 9120 17282 9172
rect 18874 9160 18880 9172
rect 18708 9132 18880 9160
rect 16485 9095 16543 9101
rect 16485 9061 16497 9095
rect 16531 9061 16543 9095
rect 16485 9055 16543 9061
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 11379 8860 12434 8888
rect 14108 8888 14136 8987
rect 16209 8959 16267 8965
rect 16209 8925 16221 8959
rect 16255 8956 16267 8959
rect 17236 8956 17264 9120
rect 18708 9033 18736 9132
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 22557 9163 22615 9169
rect 22557 9160 22569 9163
rect 20404 9132 22569 9160
rect 20404 9120 20410 9132
rect 22557 9129 22569 9132
rect 22603 9160 22615 9163
rect 23658 9160 23664 9172
rect 22603 9132 23664 9160
rect 22603 9129 22615 9132
rect 22557 9123 22615 9129
rect 23658 9120 23664 9132
rect 23716 9160 23722 9172
rect 24026 9160 24032 9172
rect 23716 9132 24032 9160
rect 23716 9120 23722 9132
rect 24026 9120 24032 9132
rect 24084 9120 24090 9172
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 25317 9163 25375 9169
rect 25317 9160 25329 9163
rect 24912 9132 25329 9160
rect 24912 9120 24918 9132
rect 25317 9129 25329 9132
rect 25363 9129 25375 9163
rect 25317 9123 25375 9129
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 19306 9064 21281 9092
rect 18693 9027 18751 9033
rect 18693 8993 18705 9027
rect 18739 8993 18751 9027
rect 18693 8987 18751 8993
rect 18785 9027 18843 9033
rect 18785 8993 18797 9027
rect 18831 9024 18843 9027
rect 18966 9024 18972 9036
rect 18831 8996 18972 9024
rect 18831 8993 18843 8996
rect 18785 8987 18843 8993
rect 18966 8984 18972 8996
rect 19024 8984 19030 9036
rect 19306 8956 19334 9064
rect 21269 9061 21281 9064
rect 21315 9061 21327 9095
rect 21269 9055 21327 9061
rect 22922 9052 22928 9104
rect 22980 9092 22986 9104
rect 28166 9092 28172 9104
rect 22980 9064 28172 9092
rect 22980 9052 22986 9064
rect 28166 9052 28172 9064
rect 28224 9052 28230 9104
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 20717 9027 20775 9033
rect 20717 9024 20729 9027
rect 19576 8996 20729 9024
rect 19576 8984 19582 8996
rect 20717 8993 20729 8996
rect 20763 8993 20775 9027
rect 20717 8987 20775 8993
rect 23106 8984 23112 9036
rect 23164 8984 23170 9036
rect 23198 8984 23204 9036
rect 23256 9024 23262 9036
rect 23477 9027 23535 9033
rect 23477 9024 23489 9027
rect 23256 8996 23489 9024
rect 23256 8984 23262 8996
rect 23477 8993 23489 8996
rect 23523 8993 23535 9027
rect 23477 8987 23535 8993
rect 25314 8984 25320 9036
rect 25372 8984 25378 9036
rect 25406 8984 25412 9036
rect 25464 9024 25470 9036
rect 25501 9027 25559 9033
rect 25501 9024 25513 9027
rect 25464 8996 25513 9024
rect 25464 8984 25470 8996
rect 25501 8993 25513 8996
rect 25547 8993 25559 9027
rect 25501 8987 25559 8993
rect 16255 8928 17264 8956
rect 18616 8928 19334 8956
rect 16255 8925 16267 8928
rect 16209 8919 16267 8925
rect 17221 8891 17279 8897
rect 17221 8888 17233 8891
rect 14108 8860 17233 8888
rect 11379 8857 11391 8860
rect 11333 8851 11391 8857
rect 17221 8857 17233 8860
rect 17267 8888 17279 8891
rect 18616 8888 18644 8928
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 28258 8956 28264 8968
rect 23072 8928 28264 8956
rect 23072 8916 23078 8928
rect 28258 8916 28264 8928
rect 28316 8916 28322 8968
rect 17267 8860 18644 8888
rect 17267 8857 17279 8860
rect 17221 8851 17279 8857
rect 18874 8848 18880 8900
rect 18932 8888 18938 8900
rect 21910 8888 21916 8900
rect 18932 8860 21916 8888
rect 18932 8848 18938 8860
rect 21910 8848 21916 8860
rect 21968 8848 21974 8900
rect 10686 8780 10692 8832
rect 10744 8780 10750 8832
rect 11054 8780 11060 8832
rect 11112 8780 11118 8832
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 12802 8820 12808 8832
rect 12115 8792 12808 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 15657 8823 15715 8829
rect 15657 8789 15669 8823
rect 15703 8820 15715 8823
rect 16206 8820 16212 8832
rect 15703 8792 16212 8820
rect 15703 8789 15715 8792
rect 15657 8783 15715 8789
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16761 8823 16819 8829
rect 16761 8789 16773 8823
rect 16807 8820 16819 8823
rect 17586 8820 17592 8832
rect 16807 8792 17592 8820
rect 16807 8789 16819 8792
rect 16761 8783 16819 8789
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 17770 8780 17776 8832
rect 17828 8820 17834 8832
rect 20073 8823 20131 8829
rect 20073 8820 20085 8823
rect 17828 8792 20085 8820
rect 17828 8780 17834 8792
rect 20073 8789 20085 8792
rect 20119 8789 20131 8823
rect 20073 8783 20131 8789
rect 20990 8780 20996 8832
rect 21048 8780 21054 8832
rect 23382 8780 23388 8832
rect 23440 8820 23446 8832
rect 24765 8823 24823 8829
rect 24765 8820 24777 8823
rect 23440 8792 24777 8820
rect 23440 8780 23446 8792
rect 24765 8789 24777 8792
rect 24811 8789 24823 8823
rect 24765 8783 24823 8789
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 10229 8619 10287 8625
rect 10229 8585 10241 8619
rect 10275 8616 10287 8619
rect 10318 8616 10324 8628
rect 10275 8588 10324 8616
rect 10275 8585 10287 8588
rect 10229 8579 10287 8585
rect 10244 8548 10272 8579
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11480 8588 11897 8616
rect 11480 8576 11486 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 13354 8576 13360 8628
rect 13412 8576 13418 8628
rect 13633 8619 13691 8625
rect 13633 8585 13645 8619
rect 13679 8616 13691 8619
rect 13722 8616 13728 8628
rect 13679 8588 13728 8616
rect 13679 8585 13691 8588
rect 13633 8579 13691 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 13906 8616 13912 8628
rect 13863 8588 13912 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 15286 8616 15292 8628
rect 14292 8588 15292 8616
rect 9416 8520 10272 8548
rect 9416 8421 9444 8520
rect 10594 8480 10600 8492
rect 9508 8452 10600 8480
rect 9508 8421 9536 8452
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10704 8412 10732 8576
rect 13372 8548 13400 8576
rect 14292 8548 14320 8588
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16577 8619 16635 8625
rect 16577 8616 16589 8619
rect 16356 8588 16589 8616
rect 16356 8576 16362 8588
rect 16577 8585 16589 8588
rect 16623 8585 16635 8619
rect 16577 8579 16635 8585
rect 18509 8619 18567 8625
rect 18509 8585 18521 8619
rect 18555 8616 18567 8619
rect 19518 8616 19524 8628
rect 18555 8588 19524 8616
rect 18555 8585 18567 8588
rect 18509 8579 18567 8585
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 20772 8588 21833 8616
rect 20772 8576 20778 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 22649 8619 22707 8625
rect 22649 8585 22661 8619
rect 22695 8616 22707 8619
rect 22922 8616 22928 8628
rect 22695 8588 22928 8616
rect 22695 8585 22707 8588
rect 22649 8579 22707 8585
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 23014 8576 23020 8628
rect 23072 8576 23078 8628
rect 31662 8616 31668 8628
rect 23400 8588 31668 8616
rect 16850 8548 16856 8560
rect 13372 8520 14320 8548
rect 15396 8520 16856 8548
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 12342 8480 12348 8492
rect 11204 8452 12348 8480
rect 11204 8440 11210 8452
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 15396 8480 15424 8520
rect 16850 8508 16856 8520
rect 16908 8508 16914 8560
rect 23400 8557 23428 8588
rect 31662 8576 31668 8588
rect 31720 8576 31726 8628
rect 19153 8551 19211 8557
rect 19153 8517 19165 8551
rect 19199 8548 19211 8551
rect 23385 8551 23443 8557
rect 19199 8520 21680 8548
rect 19199 8517 19211 8520
rect 19153 8511 19211 8517
rect 21652 8492 21680 8520
rect 23385 8517 23397 8551
rect 23431 8517 23443 8551
rect 23385 8511 23443 8517
rect 15120 8452 15424 8480
rect 9723 8384 10732 8412
rect 11517 8415 11575 8421
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 13630 8412 13636 8424
rect 11563 8384 13636 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 15120 8412 15148 8452
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 15528 8452 17264 8480
rect 15528 8440 15534 8452
rect 13771 8384 15148 8412
rect 15197 8415 15255 8421
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 15197 8381 15209 8415
rect 15243 8412 15255 8415
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 15243 8384 17141 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17236 8412 17264 8452
rect 21634 8440 21640 8492
rect 21692 8480 21698 8492
rect 21692 8452 23980 8480
rect 21692 8440 21698 8452
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 17236 8384 20545 8412
rect 17129 8375 17187 8381
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 20533 8375 20591 8381
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8412 23259 8415
rect 23290 8412 23296 8424
rect 23247 8384 23296 8412
rect 23247 8381 23259 8384
rect 23201 8375 23259 8381
rect 9309 8347 9367 8353
rect 9309 8313 9321 8347
rect 9355 8344 9367 8347
rect 9355 8316 9812 8344
rect 9355 8313 9367 8316
rect 9309 8307 9367 8313
rect 9674 8236 9680 8288
rect 9732 8236 9738 8288
rect 9784 8276 9812 8316
rect 11238 8304 11244 8356
rect 11296 8344 11302 8356
rect 13357 8347 13415 8353
rect 11296 8316 12434 8344
rect 11296 8304 11302 8316
rect 11974 8276 11980 8288
rect 9784 8248 11980 8276
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 12406 8276 12434 8316
rect 13357 8313 13369 8347
rect 13403 8344 13415 8347
rect 13403 8316 14872 8344
rect 13403 8313 13415 8316
rect 13357 8307 13415 8313
rect 13722 8276 13728 8288
rect 12406 8248 13728 8276
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 14844 8276 14872 8316
rect 14918 8304 14924 8356
rect 14976 8353 14982 8356
rect 14976 8344 14988 8353
rect 14976 8316 15021 8344
rect 14976 8307 14988 8316
rect 14976 8304 14982 8307
rect 15102 8304 15108 8356
rect 15160 8344 15166 8356
rect 15212 8344 15240 8375
rect 23290 8372 23296 8384
rect 23348 8372 23354 8424
rect 23569 8415 23627 8421
rect 23569 8381 23581 8415
rect 23615 8381 23627 8415
rect 23569 8375 23627 8381
rect 15160 8316 15240 8344
rect 15160 8304 15166 8316
rect 15286 8304 15292 8356
rect 15344 8304 15350 8356
rect 16206 8344 16212 8356
rect 15396 8316 16212 8344
rect 15396 8276 15424 8316
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 17396 8347 17454 8353
rect 17396 8313 17408 8347
rect 17442 8344 17454 8347
rect 20441 8347 20499 8353
rect 17442 8316 18736 8344
rect 17442 8313 17454 8316
rect 17396 8307 17454 8313
rect 14844 8248 15424 8276
rect 18708 8276 18736 8316
rect 20441 8313 20453 8347
rect 20487 8344 20499 8347
rect 22646 8344 22652 8356
rect 20487 8316 22652 8344
rect 20487 8313 20499 8316
rect 20441 8307 20499 8313
rect 22646 8304 22652 8316
rect 22704 8304 22710 8356
rect 22741 8347 22799 8353
rect 22741 8313 22753 8347
rect 22787 8344 22799 8347
rect 23584 8344 23612 8375
rect 23658 8372 23664 8424
rect 23716 8412 23722 8424
rect 23845 8415 23903 8421
rect 23845 8412 23857 8415
rect 23716 8384 23857 8412
rect 23716 8372 23722 8384
rect 23845 8381 23857 8384
rect 23891 8381 23903 8415
rect 23952 8412 23980 8452
rect 25317 8415 25375 8421
rect 25317 8412 25329 8415
rect 23952 8384 25329 8412
rect 23845 8375 23903 8381
rect 25317 8381 25329 8384
rect 25363 8381 25375 8415
rect 25317 8375 25375 8381
rect 25498 8372 25504 8424
rect 25556 8412 25562 8424
rect 25593 8415 25651 8421
rect 25593 8412 25605 8415
rect 25556 8384 25605 8412
rect 25556 8372 25562 8384
rect 25593 8381 25605 8384
rect 25639 8381 25651 8415
rect 25593 8375 25651 8381
rect 23934 8344 23940 8356
rect 22787 8316 23520 8344
rect 23584 8316 23940 8344
rect 22787 8313 22799 8316
rect 22741 8307 22799 8313
rect 18874 8276 18880 8288
rect 18708 8248 18880 8276
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 20162 8236 20168 8288
rect 20220 8276 20226 8288
rect 23106 8276 23112 8288
rect 20220 8248 23112 8276
rect 20220 8236 20226 8248
rect 23106 8236 23112 8248
rect 23164 8236 23170 8288
rect 23492 8276 23520 8316
rect 23934 8304 23940 8316
rect 23992 8304 23998 8356
rect 24118 8353 24124 8356
rect 24090 8347 24124 8353
rect 24090 8313 24102 8347
rect 24090 8307 24124 8313
rect 24118 8304 24124 8307
rect 24176 8304 24182 8356
rect 24228 8316 24854 8344
rect 24228 8276 24256 8316
rect 23492 8248 24256 8276
rect 24826 8276 24854 8316
rect 25225 8279 25283 8285
rect 25225 8276 25237 8279
rect 24826 8248 25237 8276
rect 25225 8245 25237 8248
rect 25271 8245 25283 8279
rect 25225 8239 25283 8245
rect 25406 8236 25412 8288
rect 25464 8236 25470 8288
rect 25682 8236 25688 8288
rect 25740 8236 25746 8288
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10100 8044 10149 8072
rect 10100 8032 10106 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 11054 8032 11060 8084
rect 11112 8032 11118 8084
rect 11238 8032 11244 8084
rect 11296 8032 11302 8084
rect 11532 8044 12296 8072
rect 11072 8004 11100 8032
rect 11256 8004 11284 8032
rect 10336 7976 11100 8004
rect 11164 7976 11284 8004
rect 10336 7945 10364 7976
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7905 10287 7939
rect 10229 7899 10287 7905
rect 10321 7939 10379 7945
rect 10321 7905 10333 7939
rect 10367 7905 10379 7939
rect 10321 7899 10379 7905
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10244 7868 10272 7899
rect 10410 7868 10416 7880
rect 10244 7840 10416 7868
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 10520 7868 10548 7899
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 10689 7939 10747 7945
rect 10689 7936 10701 7939
rect 10652 7908 10701 7936
rect 10652 7896 10658 7908
rect 10689 7905 10701 7908
rect 10735 7905 10747 7939
rect 10689 7899 10747 7905
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7936 10839 7939
rect 11164 7936 11192 7976
rect 10827 7908 11192 7936
rect 10827 7905 10839 7908
rect 10781 7899 10839 7905
rect 11238 7896 11244 7948
rect 11296 7896 11302 7948
rect 11532 7945 11560 8044
rect 12268 8004 12296 8044
rect 13630 8032 13636 8084
rect 13688 8032 13694 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 13872 8044 15669 8072
rect 13872 8032 13878 8044
rect 15657 8041 15669 8044
rect 15703 8072 15715 8075
rect 16850 8072 16856 8084
rect 15703 8044 16856 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17034 8072 17040 8084
rect 16991 8044 17040 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 18509 8075 18567 8081
rect 18509 8072 18521 8075
rect 17552 8044 18521 8072
rect 17552 8032 17558 8044
rect 18509 8041 18521 8044
rect 18555 8041 18567 8075
rect 18509 8035 18567 8041
rect 20349 8075 20407 8081
rect 20349 8041 20361 8075
rect 20395 8072 20407 8075
rect 20438 8072 20444 8084
rect 20395 8044 20444 8072
rect 20395 8041 20407 8044
rect 20349 8035 20407 8041
rect 20438 8032 20444 8044
rect 20496 8032 20502 8084
rect 22646 8032 22652 8084
rect 22704 8072 22710 8084
rect 22741 8075 22799 8081
rect 22741 8072 22753 8075
rect 22704 8044 22753 8072
rect 22704 8032 22710 8044
rect 22741 8041 22753 8044
rect 22787 8072 22799 8075
rect 23198 8072 23204 8084
rect 22787 8044 23204 8072
rect 22787 8041 22799 8044
rect 22741 8035 22799 8041
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 12268 7976 17448 8004
rect 17420 7948 17448 7976
rect 21174 7964 21180 8016
rect 21232 8004 21238 8016
rect 23109 8007 23167 8013
rect 23109 8004 23121 8007
rect 21232 7976 23121 8004
rect 21232 7964 21238 7976
rect 23109 7973 23121 7976
rect 23155 7973 23167 8007
rect 23109 7967 23167 7973
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7905 11575 7939
rect 11885 7939 11943 7945
rect 11517 7899 11575 7905
rect 11624 7908 11836 7936
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 10520 7840 11161 7868
rect 11149 7837 11161 7840
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11624 7868 11652 7908
rect 11471 7840 11652 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11698 7760 11704 7812
rect 11756 7760 11762 7812
rect 11808 7800 11836 7908
rect 11885 7905 11897 7939
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 11900 7868 11928 7899
rect 11974 7896 11980 7948
rect 12032 7896 12038 7948
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 12124 7908 12357 7936
rect 12124 7896 12130 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 14056 7908 14197 7936
rect 14056 7896 14062 7908
rect 14185 7905 14197 7908
rect 14231 7936 14243 7939
rect 15378 7936 15384 7948
rect 14231 7908 15384 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 16209 7939 16267 7945
rect 16209 7905 16221 7939
rect 16255 7936 16267 7939
rect 16298 7936 16304 7948
rect 16255 7908 16304 7936
rect 16255 7905 16267 7908
rect 16209 7899 16267 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 17126 7896 17132 7948
rect 17184 7896 17190 7948
rect 17218 7896 17224 7948
rect 17276 7896 17282 7948
rect 17402 7896 17408 7948
rect 17460 7896 17466 7948
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 19061 7939 19119 7945
rect 19061 7936 19073 7939
rect 18196 7908 19073 7936
rect 18196 7896 18202 7908
rect 19061 7905 19073 7908
rect 19107 7905 19119 7939
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 19061 7899 19119 7905
rect 20640 7908 20913 7936
rect 11900 7840 12434 7868
rect 12406 7800 12434 7840
rect 17034 7828 17040 7880
rect 17092 7868 17098 7880
rect 17494 7868 17500 7880
rect 17092 7840 17500 7868
rect 17092 7828 17098 7840
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 20640 7812 20668 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7936 21327 7939
rect 22094 7936 22100 7948
rect 21315 7908 22100 7936
rect 21315 7905 21327 7908
rect 21269 7899 21327 7905
rect 22094 7896 22100 7908
rect 22152 7896 22158 7948
rect 12894 7800 12900 7812
rect 11808 7772 12296 7800
rect 12406 7772 12900 7800
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 12161 7735 12219 7741
rect 12161 7732 12173 7735
rect 11664 7704 12173 7732
rect 11664 7692 11670 7704
rect 12161 7701 12173 7704
rect 12207 7701 12219 7735
rect 12268 7732 12296 7772
rect 12894 7760 12900 7772
rect 12952 7760 12958 7812
rect 20622 7760 20628 7812
rect 20680 7760 20686 7812
rect 14642 7732 14648 7744
rect 12268 7704 14648 7732
rect 12161 7695 12219 7701
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 16485 7735 16543 7741
rect 16485 7701 16497 7735
rect 16531 7732 16543 7735
rect 16574 7732 16580 7744
rect 16531 7704 16580 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 16666 7692 16672 7744
rect 16724 7732 16730 7744
rect 20993 7735 21051 7741
rect 20993 7732 21005 7735
rect 16724 7704 21005 7732
rect 16724 7692 16730 7704
rect 20993 7701 21005 7704
rect 21039 7701 21051 7735
rect 20993 7695 21051 7701
rect 23198 7692 23204 7744
rect 23256 7732 23262 7744
rect 24397 7735 24455 7741
rect 24397 7732 24409 7735
rect 23256 7704 24409 7732
rect 23256 7692 23262 7704
rect 24397 7701 24409 7704
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 10410 7488 10416 7540
rect 10468 7488 10474 7540
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 10560 7500 15853 7528
rect 10560 7488 10566 7500
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 15841 7491 15899 7497
rect 19889 7531 19947 7537
rect 19889 7497 19901 7531
rect 19935 7528 19947 7531
rect 28442 7528 28448 7540
rect 19935 7500 28448 7528
rect 19935 7497 19947 7500
rect 19889 7491 19947 7497
rect 28442 7488 28448 7500
rect 28500 7488 28506 7540
rect 10428 7392 10456 7488
rect 16850 7420 16856 7472
rect 16908 7460 16914 7472
rect 19242 7460 19248 7472
rect 16908 7432 19248 7460
rect 16908 7420 16914 7432
rect 19242 7420 19248 7432
rect 19300 7420 19306 7472
rect 20717 7463 20775 7469
rect 20717 7429 20729 7463
rect 20763 7460 20775 7463
rect 21174 7460 21180 7472
rect 20763 7432 21180 7460
rect 20763 7429 20775 7432
rect 20717 7423 20775 7429
rect 21174 7420 21180 7432
rect 21232 7420 21238 7472
rect 23477 7395 23535 7401
rect 10428 7364 16436 7392
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11020 7296 11836 7324
rect 11020 7284 11026 7296
rect 11808 7265 11836 7296
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 12676 7296 13645 7324
rect 12676 7284 12682 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14553 7327 14611 7333
rect 14553 7324 14565 7327
rect 13780 7296 14565 7324
rect 13780 7284 13786 7296
rect 14553 7293 14565 7296
rect 14599 7293 14611 7327
rect 14553 7287 14611 7293
rect 14918 7284 14924 7336
rect 14976 7284 14982 7336
rect 16408 7333 16436 7364
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 24026 7392 24032 7404
rect 23523 7364 24032 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 24026 7352 24032 7364
rect 24084 7352 24090 7404
rect 16393 7327 16451 7333
rect 16393 7293 16405 7327
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 18506 7284 18512 7336
rect 18564 7284 18570 7336
rect 20073 7327 20131 7333
rect 20073 7293 20085 7327
rect 20119 7324 20131 7327
rect 20530 7324 20536 7336
rect 20119 7296 20536 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 20530 7284 20536 7296
rect 20588 7284 20594 7336
rect 11517 7259 11575 7265
rect 11517 7225 11529 7259
rect 11563 7225 11575 7259
rect 11517 7219 11575 7225
rect 11793 7259 11851 7265
rect 11793 7225 11805 7259
rect 11839 7256 11851 7259
rect 11882 7256 11888 7268
rect 11839 7228 11888 7256
rect 11839 7225 11851 7228
rect 11793 7219 11851 7225
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 11422 7188 11428 7200
rect 10275 7160 11428 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 11532 7188 11560 7219
rect 11882 7216 11888 7228
rect 11940 7216 11946 7268
rect 13357 7259 13415 7265
rect 13357 7225 13369 7259
rect 13403 7256 13415 7259
rect 13998 7256 14004 7268
rect 13403 7228 14004 7256
rect 13403 7225 13415 7228
rect 13357 7219 13415 7225
rect 13998 7216 14004 7228
rect 14056 7216 14062 7268
rect 14093 7259 14151 7265
rect 14093 7225 14105 7259
rect 14139 7256 14151 7259
rect 14936 7256 14964 7284
rect 14139 7228 14964 7256
rect 14139 7225 14151 7228
rect 14093 7219 14151 7225
rect 18230 7216 18236 7268
rect 18288 7256 18294 7268
rect 18785 7259 18843 7265
rect 18785 7256 18797 7259
rect 18288 7228 18797 7256
rect 18288 7216 18294 7228
rect 18785 7225 18797 7228
rect 18831 7225 18843 7259
rect 18785 7219 18843 7225
rect 19153 7259 19211 7265
rect 19153 7225 19165 7259
rect 19199 7225 19211 7259
rect 19153 7219 19211 7225
rect 19337 7259 19395 7265
rect 19337 7225 19349 7259
rect 19383 7256 19395 7259
rect 19610 7256 19616 7268
rect 19383 7228 19616 7256
rect 19383 7225 19395 7228
rect 19337 7219 19395 7225
rect 13262 7188 13268 7200
rect 11532 7160 13268 7188
rect 13262 7148 13268 7160
rect 13320 7188 13326 7200
rect 13630 7188 13636 7200
rect 13320 7160 13636 7188
rect 13320 7148 13326 7160
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13814 7148 13820 7200
rect 13872 7148 13878 7200
rect 14182 7148 14188 7200
rect 14240 7148 14246 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 17681 7191 17739 7197
rect 17681 7188 17693 7191
rect 15436 7160 17693 7188
rect 15436 7148 15442 7160
rect 17681 7157 17693 7160
rect 17727 7188 17739 7191
rect 18966 7188 18972 7200
rect 17727 7160 18972 7188
rect 17727 7157 17739 7160
rect 17681 7151 17739 7157
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 19168 7188 19196 7219
rect 19610 7216 19616 7228
rect 19668 7216 19674 7268
rect 19705 7259 19763 7265
rect 19705 7225 19717 7259
rect 19751 7256 19763 7259
rect 20254 7256 20260 7268
rect 19751 7228 20260 7256
rect 19751 7225 19763 7228
rect 19705 7219 19763 7225
rect 20254 7216 20260 7228
rect 20312 7216 20318 7268
rect 22005 7259 22063 7265
rect 22005 7225 22017 7259
rect 22051 7256 22063 7259
rect 22370 7256 22376 7268
rect 22051 7228 22376 7256
rect 22051 7225 22063 7228
rect 22005 7219 22063 7225
rect 22370 7216 22376 7228
rect 22428 7216 22434 7268
rect 23014 7216 23020 7268
rect 23072 7256 23078 7268
rect 23210 7259 23268 7265
rect 23210 7256 23222 7259
rect 23072 7228 23222 7256
rect 23072 7216 23078 7228
rect 23210 7225 23222 7228
rect 23256 7225 23268 7259
rect 23210 7219 23268 7225
rect 20346 7188 20352 7200
rect 19168 7160 20352 7188
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 22097 7191 22155 7197
rect 22097 7157 22109 7191
rect 22143 7188 22155 7191
rect 22186 7188 22192 7200
rect 22143 7160 22192 7188
rect 22143 7157 22155 7160
rect 22097 7151 22155 7157
rect 22186 7148 22192 7160
rect 22244 7148 22250 7200
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 13630 6944 13636 6996
rect 13688 6944 13694 6996
rect 17402 6944 17408 6996
rect 17460 6944 17466 6996
rect 22370 6944 22376 6996
rect 22428 6944 22434 6996
rect 23014 6944 23020 6996
rect 23072 6944 23078 6996
rect 17972 6888 18552 6916
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 11256 6780 11284 6811
rect 11422 6808 11428 6860
rect 11480 6808 11486 6860
rect 11701 6851 11759 6857
rect 11701 6817 11713 6851
rect 11747 6848 11759 6851
rect 11790 6848 11796 6860
rect 11747 6820 11796 6848
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11256 6752 11621 6780
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 12176 6780 12204 6811
rect 12342 6808 12348 6860
rect 12400 6808 12406 6860
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 12434 6780 12440 6792
rect 12176 6752 12440 6780
rect 11609 6743 11667 6749
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 11333 6715 11391 6721
rect 11333 6681 11345 6715
rect 11379 6712 11391 6715
rect 14200 6712 14228 6811
rect 16114 6808 16120 6860
rect 16172 6808 16178 6860
rect 17972 6857 18000 6888
rect 18524 6860 18552 6888
rect 19242 6876 19248 6928
rect 19300 6916 19306 6928
rect 20622 6916 20628 6928
rect 19300 6888 20628 6916
rect 19300 6876 19306 6888
rect 20622 6876 20628 6888
rect 20680 6876 20686 6928
rect 22186 6876 22192 6928
rect 22244 6876 22250 6928
rect 22296 6888 22876 6916
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17935 6820 17969 6848
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18213 6851 18271 6857
rect 18213 6848 18225 6851
rect 18104 6820 18225 6848
rect 18104 6808 18110 6820
rect 18213 6817 18225 6820
rect 18259 6817 18271 6851
rect 18213 6811 18271 6817
rect 18506 6808 18512 6860
rect 18564 6848 18570 6860
rect 18564 6820 19012 6848
rect 18564 6808 18570 6820
rect 18984 6780 19012 6820
rect 19150 6808 19156 6860
rect 19208 6848 19214 6860
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 19208 6820 19441 6848
rect 19208 6808 19214 6820
rect 19429 6817 19441 6820
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 19972 6851 20030 6857
rect 19972 6817 19984 6851
rect 20018 6848 20030 6851
rect 21361 6851 21419 6857
rect 20018 6820 20852 6848
rect 20018 6817 20030 6820
rect 19972 6811 20030 6817
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 18984 6752 19717 6780
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 11379 6684 14228 6712
rect 19337 6715 19395 6721
rect 11379 6681 11391 6684
rect 11333 6675 11391 6681
rect 19337 6681 19349 6715
rect 19383 6712 19395 6715
rect 19610 6712 19616 6724
rect 19383 6684 19616 6712
rect 19383 6681 19395 6684
rect 19337 6675 19395 6681
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 20824 6656 20852 6820
rect 21361 6817 21373 6851
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6848 21787 6851
rect 22296 6848 22324 6888
rect 21775 6820 22324 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 21085 6715 21143 6721
rect 21085 6681 21097 6715
rect 21131 6712 21143 6715
rect 21376 6712 21404 6811
rect 22370 6808 22376 6860
rect 22428 6808 22434 6860
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6817 22615 6851
rect 22557 6811 22615 6817
rect 22649 6851 22707 6857
rect 22649 6817 22661 6851
rect 22695 6848 22707 6851
rect 22738 6848 22744 6860
rect 22695 6820 22744 6848
rect 22695 6817 22707 6820
rect 22649 6811 22707 6817
rect 21818 6740 21824 6792
rect 21876 6780 21882 6792
rect 22572 6780 22600 6811
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 21876 6752 22600 6780
rect 22848 6780 22876 6888
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6848 23167 6851
rect 23382 6848 23388 6860
rect 23155 6820 23388 6848
rect 23155 6817 23167 6820
rect 23109 6811 23167 6817
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 28258 6780 28264 6792
rect 22848 6752 28264 6780
rect 21876 6740 21882 6752
rect 28258 6740 28264 6752
rect 28316 6740 28322 6792
rect 21131 6684 21404 6712
rect 21131 6681 21143 6684
rect 21085 6675 21143 6681
rect 21542 6672 21548 6724
rect 21600 6712 21606 6724
rect 23842 6712 23848 6724
rect 21600 6684 23848 6712
rect 21600 6672 21606 6684
rect 23842 6672 23848 6684
rect 23900 6672 23906 6724
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6644 12127 6647
rect 13538 6644 13544 6656
rect 12115 6616 13544 6644
rect 12115 6613 12127 6616
rect 12069 6607 12127 6613
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 15654 6604 15660 6656
rect 15712 6604 15718 6656
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 19242 6644 19248 6656
rect 17920 6616 19248 6644
rect 17920 6604 17926 6616
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19518 6604 19524 6656
rect 19576 6604 19582 6656
rect 20806 6604 20812 6656
rect 20864 6604 20870 6656
rect 21913 6647 21971 6653
rect 21913 6613 21925 6647
rect 21959 6644 21971 6647
rect 22002 6644 22008 6656
rect 21959 6616 22008 6644
rect 21959 6613 21971 6616
rect 21913 6607 21971 6613
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 22741 6647 22799 6653
rect 22741 6644 22753 6647
rect 22244 6616 22753 6644
rect 22244 6604 22250 6616
rect 22741 6613 22753 6616
rect 22787 6613 22799 6647
rect 22741 6607 22799 6613
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12434 6440 12440 6452
rect 12023 6412 12440 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 17129 6443 17187 6449
rect 17129 6409 17141 6443
rect 17175 6440 17187 6443
rect 18230 6440 18236 6452
rect 17175 6412 18236 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 18782 6400 18788 6452
rect 18840 6400 18846 6452
rect 19518 6400 19524 6452
rect 19576 6400 19582 6452
rect 21818 6400 21824 6452
rect 21876 6400 21882 6452
rect 22094 6400 22100 6452
rect 22152 6400 22158 6452
rect 14093 6375 14151 6381
rect 14093 6341 14105 6375
rect 14139 6341 14151 6375
rect 14093 6335 14151 6341
rect 17313 6375 17371 6381
rect 17313 6341 17325 6375
rect 17359 6372 17371 6375
rect 17954 6372 17960 6384
rect 17359 6344 17960 6372
rect 17359 6341 17371 6344
rect 17313 6335 17371 6341
rect 14108 6304 14136 6335
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 19536 6304 19564 6400
rect 22373 6375 22431 6381
rect 22373 6372 22385 6375
rect 14108 6276 15516 6304
rect 15488 6248 15516 6276
rect 17512 6276 19564 6304
rect 19720 6344 22385 6372
rect 12526 6196 12532 6248
rect 12584 6236 12590 6248
rect 13357 6239 13415 6245
rect 13357 6236 13369 6239
rect 12584 6208 13369 6236
rect 12584 6196 12590 6208
rect 13357 6205 13369 6208
rect 13403 6205 13415 6239
rect 13357 6199 13415 6205
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 13090 6171 13148 6177
rect 13090 6168 13102 6171
rect 12400 6140 13102 6168
rect 12400 6128 12406 6140
rect 13090 6137 13102 6140
rect 13136 6137 13148 6171
rect 13372 6168 13400 6199
rect 15378 6196 15384 6248
rect 15436 6196 15442 6248
rect 15470 6196 15476 6248
rect 15528 6196 15534 6248
rect 17512 6245 17540 6276
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 17497 6239 17555 6245
rect 17497 6205 17509 6239
rect 17543 6205 17555 6239
rect 17497 6199 17555 6205
rect 14550 6168 14556 6180
rect 13372 6140 14556 6168
rect 13090 6131 13148 6137
rect 14550 6128 14556 6140
rect 14608 6168 14614 6180
rect 15764 6168 15792 6199
rect 17770 6196 17776 6248
rect 17828 6196 17834 6248
rect 18322 6196 18328 6248
rect 18380 6196 18386 6248
rect 18690 6196 18696 6248
rect 18748 6196 18754 6248
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6236 19487 6239
rect 19720 6236 19748 6344
rect 22373 6341 22385 6344
rect 22419 6341 22431 6375
rect 22373 6335 22431 6341
rect 19886 6264 19892 6316
rect 19944 6304 19950 6316
rect 21542 6304 21548 6316
rect 19944 6276 21548 6304
rect 19944 6264 19950 6276
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 25682 6304 25688 6316
rect 22020 6276 25688 6304
rect 19475 6208 19748 6236
rect 19475 6205 19487 6208
rect 19429 6199 19487 6205
rect 19794 6196 19800 6248
rect 19852 6196 19858 6248
rect 21726 6196 21732 6248
rect 21784 6196 21790 6248
rect 22020 6247 22048 6276
rect 25682 6264 25688 6276
rect 25740 6264 25746 6316
rect 22005 6241 22063 6247
rect 22005 6207 22017 6241
rect 22051 6207 22063 6241
rect 22005 6201 22063 6207
rect 22186 6196 22192 6248
rect 22244 6196 22250 6248
rect 22281 6239 22339 6245
rect 22281 6205 22293 6239
rect 22327 6238 22339 6239
rect 22327 6210 22416 6238
rect 22327 6205 22339 6210
rect 22281 6199 22339 6205
rect 14608 6140 15792 6168
rect 16016 6171 16074 6177
rect 14608 6128 14614 6140
rect 16016 6137 16028 6171
rect 16062 6168 16074 6171
rect 16206 6168 16212 6180
rect 16062 6140 16212 6168
rect 16062 6137 16074 6140
rect 16016 6131 16074 6137
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 19334 6128 19340 6180
rect 19392 6168 19398 6180
rect 19889 6171 19947 6177
rect 19889 6168 19901 6171
rect 19392 6140 19901 6168
rect 19392 6128 19398 6140
rect 19889 6137 19901 6140
rect 19935 6137 19947 6171
rect 19889 6131 19947 6137
rect 15562 6060 15568 6112
rect 15620 6060 15626 6112
rect 17678 6060 17684 6112
rect 17736 6060 17742 6112
rect 18141 6103 18199 6109
rect 18141 6069 18153 6103
rect 18187 6100 18199 6103
rect 18690 6100 18696 6112
rect 18187 6072 18696 6100
rect 18187 6069 18199 6072
rect 18141 6063 18199 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 19242 6060 19248 6112
rect 19300 6060 19306 6112
rect 19613 6103 19671 6109
rect 19613 6069 19625 6103
rect 19659 6100 19671 6103
rect 21082 6100 21088 6112
rect 19659 6072 21088 6100
rect 19659 6069 19671 6072
rect 19613 6063 19671 6069
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 21174 6060 21180 6112
rect 21232 6060 21238 6112
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 22388 6100 22416 6210
rect 22060 6072 22416 6100
rect 22060 6060 22066 6072
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 11422 5856 11428 5908
rect 11480 5856 11486 5908
rect 12342 5856 12348 5908
rect 12400 5856 12406 5908
rect 12894 5856 12900 5908
rect 12952 5856 12958 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15620 5868 16574 5896
rect 15620 5856 15626 5868
rect 11440 5692 11468 5856
rect 11790 5788 11796 5840
rect 11848 5828 11854 5840
rect 11848 5800 13308 5828
rect 11848 5788 11854 5800
rect 11514 5720 11520 5772
rect 11572 5760 11578 5772
rect 13280 5769 13308 5800
rect 15654 5788 15660 5840
rect 15712 5828 15718 5840
rect 15749 5831 15807 5837
rect 15749 5828 15761 5831
rect 15712 5800 15761 5828
rect 15712 5788 15718 5800
rect 15749 5797 15761 5800
rect 15795 5797 15807 5831
rect 15749 5791 15807 5797
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 11572 5732 12449 5760
rect 11572 5720 11578 5732
rect 12437 5729 12449 5732
rect 12483 5760 12495 5763
rect 12805 5763 12863 5769
rect 12805 5760 12817 5763
rect 12483 5732 12817 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 12805 5729 12817 5732
rect 12851 5729 12863 5763
rect 12805 5723 12863 5729
rect 13265 5763 13323 5769
rect 13265 5729 13277 5763
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 13906 5720 13912 5772
rect 13964 5720 13970 5772
rect 15562 5720 15568 5772
rect 15620 5760 15626 5772
rect 16209 5763 16267 5769
rect 16209 5760 16221 5763
rect 15620 5732 16221 5760
rect 15620 5720 15626 5732
rect 16209 5729 16221 5732
rect 16255 5729 16267 5763
rect 16546 5760 16574 5868
rect 19150 5856 19156 5908
rect 19208 5856 19214 5908
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19484 5868 19625 5896
rect 19484 5856 19490 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 19613 5859 19671 5865
rect 19981 5899 20039 5905
rect 19981 5865 19993 5899
rect 20027 5896 20039 5899
rect 20162 5896 20168 5908
rect 20027 5868 20168 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 20714 5856 20720 5908
rect 20772 5856 20778 5908
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 21637 5899 21695 5905
rect 21637 5896 21649 5899
rect 20864 5868 21649 5896
rect 20864 5856 20870 5868
rect 21637 5865 21649 5868
rect 21683 5865 21695 5899
rect 22370 5896 22376 5908
rect 21637 5859 21695 5865
rect 21744 5868 22376 5896
rect 17034 5788 17040 5840
rect 17092 5828 17098 5840
rect 17221 5831 17279 5837
rect 17221 5828 17233 5831
rect 17092 5800 17233 5828
rect 17092 5788 17098 5800
rect 17221 5797 17233 5800
rect 17267 5797 17279 5831
rect 17221 5791 17279 5797
rect 18969 5831 19027 5837
rect 18969 5797 18981 5831
rect 19015 5828 19027 5831
rect 19168 5828 19196 5856
rect 19886 5828 19892 5840
rect 19015 5800 19196 5828
rect 19536 5800 19892 5828
rect 19015 5797 19027 5800
rect 18969 5791 19027 5797
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 16546 5732 16681 5760
rect 16209 5723 16267 5729
rect 16669 5729 16681 5732
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 19058 5720 19064 5772
rect 19116 5720 19122 5772
rect 19536 5769 19564 5800
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 20732 5828 20760 5856
rect 21744 5828 21772 5868
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 20088 5800 20760 5828
rect 19153 5763 19211 5769
rect 19153 5729 19165 5763
rect 19199 5760 19211 5763
rect 19337 5763 19395 5769
rect 19337 5760 19349 5763
rect 19199 5732 19349 5760
rect 19199 5729 19211 5732
rect 19153 5723 19211 5729
rect 19337 5729 19349 5732
rect 19383 5729 19395 5763
rect 19337 5723 19395 5729
rect 19521 5763 19579 5769
rect 19521 5729 19533 5763
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 19610 5720 19616 5772
rect 19668 5720 19674 5772
rect 19794 5720 19800 5772
rect 19852 5720 19858 5772
rect 19978 5720 19984 5772
rect 20036 5720 20042 5772
rect 20088 5769 20116 5800
rect 20073 5763 20131 5769
rect 20073 5729 20085 5763
rect 20119 5729 20131 5763
rect 20073 5723 20131 5729
rect 20165 5763 20223 5769
rect 20165 5729 20177 5763
rect 20211 5760 20223 5763
rect 20530 5760 20536 5772
rect 20211 5732 20536 5760
rect 20211 5729 20223 5732
rect 20165 5723 20223 5729
rect 20530 5720 20536 5732
rect 20588 5720 20594 5772
rect 20622 5720 20628 5772
rect 20680 5720 20686 5772
rect 20732 5769 20760 5800
rect 20824 5800 21772 5828
rect 20824 5769 20852 5800
rect 22002 5788 22008 5840
rect 22060 5788 22066 5840
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5729 20775 5763
rect 20717 5723 20775 5729
rect 20809 5763 20867 5769
rect 20809 5729 20821 5763
rect 20855 5729 20867 5763
rect 20809 5723 20867 5729
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5729 21511 5763
rect 21453 5723 21511 5729
rect 21729 5763 21787 5769
rect 21729 5729 21741 5763
rect 21775 5760 21787 5763
rect 22020 5760 22048 5788
rect 21775 5732 22048 5760
rect 21775 5729 21787 5732
rect 21729 5723 21787 5729
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 11440 5664 13369 5692
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 19429 5695 19487 5701
rect 19429 5661 19441 5695
rect 19475 5692 19487 5695
rect 19996 5692 20024 5720
rect 19475 5664 20024 5692
rect 21468 5692 21496 5723
rect 23198 5692 23204 5704
rect 21468 5664 23204 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 23198 5652 23204 5664
rect 23256 5652 23262 5704
rect 19242 5584 19248 5636
rect 19300 5624 19306 5636
rect 21361 5627 21419 5633
rect 19300 5596 21312 5624
rect 19300 5584 19306 5596
rect 13725 5559 13783 5565
rect 13725 5525 13737 5559
rect 13771 5556 13783 5559
rect 14182 5556 14188 5568
rect 13771 5528 14188 5556
rect 13771 5525 13783 5528
rect 13725 5519 13783 5525
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 14458 5516 14464 5568
rect 14516 5516 14522 5568
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 15712 5528 16313 5556
rect 15712 5516 15718 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 16301 5519 16359 5525
rect 16390 5516 16396 5568
rect 16448 5556 16454 5568
rect 16853 5559 16911 5565
rect 16853 5556 16865 5559
rect 16448 5528 16865 5556
rect 16448 5516 16454 5528
rect 16853 5525 16865 5528
rect 16899 5525 16911 5559
rect 16853 5519 16911 5525
rect 20254 5516 20260 5568
rect 20312 5516 20318 5568
rect 20530 5516 20536 5568
rect 20588 5516 20594 5568
rect 21284 5556 21312 5596
rect 21361 5593 21373 5627
rect 21407 5624 21419 5627
rect 24118 5624 24124 5636
rect 21407 5596 24124 5624
rect 21407 5593 21419 5596
rect 21361 5587 21419 5593
rect 24118 5584 24124 5596
rect 24176 5584 24182 5636
rect 22554 5556 22560 5568
rect 21284 5528 22560 5556
rect 22554 5516 22560 5528
rect 22612 5516 22618 5568
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14093 5355 14151 5361
rect 14093 5352 14105 5355
rect 13964 5324 14105 5352
rect 13964 5312 13970 5324
rect 14093 5321 14105 5324
rect 14139 5321 14151 5355
rect 14093 5315 14151 5321
rect 16117 5355 16175 5361
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 16206 5352 16212 5364
rect 16163 5324 16212 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 16298 5312 16304 5364
rect 16356 5312 16362 5364
rect 16577 5355 16635 5361
rect 16577 5321 16589 5355
rect 16623 5352 16635 5355
rect 17126 5352 17132 5364
rect 16623 5324 17132 5352
rect 16623 5321 16635 5324
rect 16577 5315 16635 5321
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 18138 5352 18144 5364
rect 18095 5324 18144 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 18322 5312 18328 5364
rect 18380 5312 18386 5364
rect 18598 5312 18604 5364
rect 18656 5352 18662 5364
rect 18969 5355 19027 5361
rect 18969 5352 18981 5355
rect 18656 5324 18981 5352
rect 18656 5312 18662 5324
rect 18969 5321 18981 5324
rect 19015 5352 19027 5355
rect 20622 5352 20628 5364
rect 19015 5324 20628 5352
rect 19015 5321 19027 5324
rect 18969 5315 19027 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 22002 5312 22008 5364
rect 22060 5312 22066 5364
rect 15933 5287 15991 5293
rect 15933 5253 15945 5287
rect 15979 5284 15991 5287
rect 16316 5284 16344 5312
rect 19150 5284 19156 5296
rect 15979 5256 16344 5284
rect 17604 5256 19156 5284
rect 15979 5253 15991 5256
rect 15933 5247 15991 5253
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 14550 5216 14556 5228
rect 14332 5188 14556 5216
rect 14332 5176 14338 5188
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 17494 5216 17500 5228
rect 16500 5188 17500 5216
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5148 14243 5151
rect 14458 5148 14464 5160
rect 14231 5120 14464 5148
rect 14231 5117 14243 5120
rect 14185 5111 14243 5117
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 14809 5151 14867 5157
rect 14809 5148 14821 5151
rect 14700 5120 14821 5148
rect 14700 5108 14706 5120
rect 14809 5117 14821 5120
rect 14855 5117 14867 5151
rect 14809 5111 14867 5117
rect 15562 5108 15568 5160
rect 15620 5148 15626 5160
rect 16500 5157 16528 5188
rect 17494 5176 17500 5188
rect 17552 5176 17558 5228
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15620 5120 16037 5148
rect 15620 5108 15626 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 16485 5151 16543 5157
rect 16485 5117 16497 5151
rect 16531 5117 16543 5151
rect 16485 5111 16543 5117
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 17604 5157 17632 5256
rect 19150 5244 19156 5256
rect 19208 5244 19214 5296
rect 17773 5219 17831 5225
rect 17773 5185 17785 5219
rect 17819 5216 17831 5219
rect 17819 5188 18184 5216
rect 17819 5185 17831 5188
rect 17773 5179 17831 5185
rect 17589 5151 17647 5157
rect 17589 5117 17601 5151
rect 17635 5117 17647 5151
rect 17589 5111 17647 5117
rect 17678 5108 17684 5160
rect 17736 5108 17742 5160
rect 18156 5157 18184 5188
rect 17957 5151 18015 5157
rect 17957 5117 17969 5151
rect 18003 5117 18015 5151
rect 17957 5111 18015 5117
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 17497 5083 17555 5089
rect 17497 5049 17509 5083
rect 17543 5080 17555 5083
rect 17972 5080 18000 5111
rect 18414 5108 18420 5160
rect 18472 5108 18478 5160
rect 20438 5108 20444 5160
rect 20496 5108 20502 5160
rect 20533 5151 20591 5157
rect 20533 5117 20545 5151
rect 20579 5148 20591 5151
rect 21174 5148 21180 5160
rect 20579 5120 21180 5148
rect 20579 5117 20591 5120
rect 20533 5111 20591 5117
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 17543 5052 18000 5080
rect 17543 5049 17555 5052
rect 17497 5043 17555 5049
rect 14366 4972 14372 5024
rect 14424 4972 14430 5024
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 15746 5012 15752 5024
rect 15528 4984 15752 5012
rect 15528 4972 15534 4984
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 14274 4768 14280 4820
rect 14332 4768 14338 4820
rect 14366 4768 14372 4820
rect 14424 4768 14430 4820
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 15654 4808 15660 4820
rect 15519 4780 15660 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 18046 4768 18052 4820
rect 18104 4768 18110 4820
rect 18598 4808 18604 4820
rect 18156 4780 18604 4808
rect 14093 4675 14151 4681
rect 14093 4641 14105 4675
rect 14139 4672 14151 4675
rect 14292 4672 14320 4768
rect 14384 4681 14412 4768
rect 18156 4681 18184 4780
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 18693 4811 18751 4817
rect 18693 4777 18705 4811
rect 18739 4808 18751 4811
rect 19334 4808 19340 4820
rect 18739 4780 19340 4808
rect 18739 4777 18751 4780
rect 18693 4771 18751 4777
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 20254 4740 20260 4752
rect 18524 4712 20260 4740
rect 18524 4681 18552 4712
rect 20254 4700 20260 4712
rect 20312 4700 20318 4752
rect 14139 4644 14320 4672
rect 14360 4675 14418 4681
rect 14139 4641 14151 4644
rect 14093 4635 14151 4641
rect 14360 4641 14372 4675
rect 14406 4641 14418 4675
rect 14360 4635 14418 4641
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 18509 4675 18567 4681
rect 18509 4641 18521 4675
rect 18555 4641 18567 4675
rect 18509 4635 18567 4641
rect 18693 4675 18751 4681
rect 18693 4641 18705 4675
rect 18739 4672 18751 4675
rect 20530 4672 20536 4684
rect 18739 4644 20536 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 20530 4632 20536 4644
rect 20588 4632 20594 4684
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 14090 3584 14096 3596
rect 9732 3556 14096 3584
rect 9732 3544 9738 3556
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 13814 3516 13820 3528
rect 11020 3488 13820 3516
rect 11020 3476 11026 3488
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 10226 3408 10232 3460
rect 10284 3448 10290 3460
rect 23198 3448 23204 3460
rect 10284 3420 23204 3448
rect 10284 3408 10290 3420
rect 23198 3408 23204 3420
rect 23256 3408 23262 3460
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 20990 2836 20996 2848
rect 19392 2808 20996 2836
rect 19392 2796 19398 2808
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
rect 16022 416 16028 468
rect 16080 456 16086 468
rect 16390 456 16396 468
rect 16080 428 16396 456
rect 16080 416 16086 428
rect 16390 416 16396 428
rect 16448 416 16454 468
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 13544 18912 13596 18964
rect 13452 18572 13504 18624
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 18696 15988 18748 16040
rect 20812 15988 20864 16040
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 19984 15376 20036 15428
rect 22192 15376 22244 15428
rect 20628 15308 20680 15360
rect 24216 15308 24268 15360
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 18144 14220 18196 14272
rect 23848 14288 23900 14340
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 18420 13948 18472 14000
rect 19524 13880 19576 13932
rect 18144 13855 18196 13864
rect 18144 13821 18153 13855
rect 18153 13821 18187 13855
rect 18187 13821 18196 13855
rect 18144 13812 18196 13821
rect 19340 13812 19392 13864
rect 20720 13948 20772 14000
rect 18328 13787 18380 13796
rect 18328 13753 18337 13787
rect 18337 13753 18371 13787
rect 18371 13753 18380 13787
rect 18328 13744 18380 13753
rect 18604 13744 18656 13796
rect 19432 13744 19484 13796
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 18052 13719 18104 13728
rect 18052 13685 18061 13719
rect 18061 13685 18095 13719
rect 18095 13685 18104 13719
rect 18052 13676 18104 13685
rect 18144 13676 18196 13728
rect 21456 13880 21508 13932
rect 21640 13812 21692 13864
rect 19892 13719 19944 13728
rect 19892 13685 19901 13719
rect 19901 13685 19935 13719
rect 19935 13685 19944 13719
rect 19892 13676 19944 13685
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 14648 13268 14700 13320
rect 18144 13404 18196 13456
rect 18696 13404 18748 13456
rect 19892 13404 19944 13456
rect 15292 13243 15344 13252
rect 15292 13209 15301 13243
rect 15301 13209 15335 13243
rect 15335 13209 15344 13243
rect 15292 13200 15344 13209
rect 18328 13379 18380 13388
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 18328 13345 18337 13379
rect 18337 13345 18371 13379
rect 18371 13345 18380 13379
rect 18328 13336 18380 13345
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 17960 13200 18012 13252
rect 20628 13336 20680 13388
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 18512 13132 18564 13184
rect 19248 13132 19300 13184
rect 21824 13132 21876 13184
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 19432 12928 19484 12980
rect 21824 12971 21876 12980
rect 21824 12937 21833 12971
rect 21833 12937 21867 12971
rect 21867 12937 21876 12971
rect 21824 12928 21876 12937
rect 13452 12724 13504 12776
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 14464 12792 14516 12844
rect 14188 12724 14240 12776
rect 15200 12792 15252 12844
rect 16212 12792 16264 12844
rect 18880 12792 18932 12844
rect 12348 12656 12400 12708
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 17684 12656 17736 12708
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 13820 12588 13872 12640
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 17960 12588 18012 12640
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 13636 12384 13688 12436
rect 11520 12316 11572 12368
rect 9588 12248 9640 12300
rect 11060 12248 11112 12300
rect 11244 12180 11296 12232
rect 12440 12248 12492 12300
rect 12716 12291 12768 12300
rect 12716 12257 12725 12291
rect 12725 12257 12759 12291
rect 12759 12257 12768 12291
rect 12716 12248 12768 12257
rect 13268 12248 13320 12300
rect 13820 12316 13872 12368
rect 18880 12427 18932 12436
rect 18880 12393 18889 12427
rect 18889 12393 18923 12427
rect 18923 12393 18932 12427
rect 18880 12384 18932 12393
rect 18788 12316 18840 12368
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 16212 12248 16264 12300
rect 19064 12248 19116 12300
rect 20720 12316 20772 12368
rect 21456 12359 21508 12368
rect 21456 12325 21465 12359
rect 21465 12325 21499 12359
rect 21499 12325 21508 12359
rect 21456 12316 21508 12325
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 22192 12427 22244 12436
rect 22192 12393 22201 12427
rect 22201 12393 22235 12427
rect 22235 12393 22244 12427
rect 22192 12384 22244 12393
rect 11612 12112 11664 12164
rect 9956 12044 10008 12096
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 12900 12044 12952 12053
rect 13820 12044 13872 12096
rect 14004 12087 14056 12096
rect 14004 12053 14013 12087
rect 14013 12053 14047 12087
rect 14047 12053 14056 12087
rect 14004 12044 14056 12053
rect 14648 12044 14700 12096
rect 20536 12112 20588 12164
rect 20352 12044 20404 12096
rect 20628 12044 20680 12096
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 11060 11883 11112 11892
rect 11060 11849 11069 11883
rect 11069 11849 11103 11883
rect 11103 11849 11112 11883
rect 11060 11840 11112 11849
rect 11244 11840 11296 11892
rect 11796 11840 11848 11892
rect 12440 11840 12492 11892
rect 12716 11840 12768 11892
rect 13544 11840 13596 11892
rect 14096 11840 14148 11892
rect 14464 11883 14516 11892
rect 14464 11849 14473 11883
rect 14473 11849 14507 11883
rect 14507 11849 14516 11883
rect 14464 11840 14516 11849
rect 15752 11840 15804 11892
rect 17684 11840 17736 11892
rect 18696 11840 18748 11892
rect 9680 11772 9732 11824
rect 9772 11704 9824 11756
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 9864 11568 9916 11620
rect 11428 11679 11480 11688
rect 11428 11645 11437 11679
rect 11437 11645 11471 11679
rect 11471 11645 11480 11679
rect 11428 11636 11480 11645
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 13176 11772 13228 11824
rect 13820 11815 13872 11824
rect 13820 11781 13829 11815
rect 13829 11781 13863 11815
rect 13863 11781 13872 11815
rect 13820 11772 13872 11781
rect 14648 11772 14700 11824
rect 12532 11636 12584 11688
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 13636 11636 13688 11688
rect 13912 11636 13964 11688
rect 14188 11636 14240 11688
rect 15752 11679 15804 11688
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 16948 11772 17000 11824
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 13268 11568 13320 11620
rect 15016 11568 15068 11620
rect 17960 11636 18012 11688
rect 18052 11636 18104 11688
rect 18328 11679 18380 11688
rect 18328 11645 18337 11679
rect 18337 11645 18371 11679
rect 18371 11645 18380 11679
rect 18328 11636 18380 11645
rect 18420 11636 18472 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 19248 11636 19300 11688
rect 22284 11636 22336 11688
rect 19432 11568 19484 11620
rect 21088 11611 21140 11620
rect 21088 11577 21097 11611
rect 21097 11577 21131 11611
rect 21131 11577 21140 11611
rect 21088 11568 21140 11577
rect 21180 11611 21232 11620
rect 21180 11577 21189 11611
rect 21189 11577 21223 11611
rect 21223 11577 21232 11611
rect 21180 11568 21232 11577
rect 24032 11568 24084 11620
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 12256 11500 12308 11552
rect 12532 11500 12584 11552
rect 14096 11500 14148 11552
rect 14556 11500 14608 11552
rect 16672 11500 16724 11552
rect 17132 11500 17184 11552
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 9588 11339 9640 11348
rect 9588 11305 9597 11339
rect 9597 11305 9631 11339
rect 9631 11305 9640 11339
rect 9588 11296 9640 11305
rect 9864 11339 9916 11348
rect 9864 11305 9873 11339
rect 9873 11305 9907 11339
rect 9907 11305 9916 11339
rect 9864 11296 9916 11305
rect 10140 11296 10192 11348
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 12256 11296 12308 11348
rect 13544 11296 13596 11348
rect 13636 11296 13688 11348
rect 9404 11160 9456 11212
rect 14464 11228 14516 11280
rect 15016 11296 15068 11348
rect 16396 11296 16448 11348
rect 18328 11296 18380 11348
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10416 11160 10468 11212
rect 9864 11092 9916 11144
rect 13912 11160 13964 11212
rect 14004 11160 14056 11212
rect 14280 11160 14332 11212
rect 18144 11228 18196 11280
rect 28264 11296 28316 11348
rect 18512 11228 18564 11280
rect 17500 11160 17552 11212
rect 19340 11203 19392 11212
rect 19340 11169 19349 11203
rect 19349 11169 19383 11203
rect 19383 11169 19392 11203
rect 19340 11160 19392 11169
rect 9680 11024 9732 11076
rect 14372 11092 14424 11144
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 22008 11160 22060 11212
rect 23204 11203 23256 11212
rect 23204 11169 23213 11203
rect 23213 11169 23247 11203
rect 23247 11169 23256 11203
rect 23204 11160 23256 11169
rect 23572 11092 23624 11144
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 10324 10956 10376 11008
rect 11336 10956 11388 11008
rect 12900 10956 12952 11008
rect 13636 10956 13688 11008
rect 16120 10956 16172 11008
rect 20076 10956 20128 11008
rect 25320 11024 25372 11076
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 9772 10752 9824 10804
rect 10232 10752 10284 10804
rect 11428 10752 11480 10804
rect 14280 10752 14332 10804
rect 14096 10684 14148 10736
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 9588 10591 9640 10600
rect 9588 10557 9607 10591
rect 9607 10557 9640 10591
rect 9588 10548 9640 10557
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 10324 10548 10376 10600
rect 10692 10616 10744 10668
rect 9772 10412 9824 10464
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 12256 10616 12308 10668
rect 13636 10616 13688 10668
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 12348 10548 12400 10600
rect 15384 10616 15436 10668
rect 14648 10591 14700 10600
rect 14648 10557 14657 10591
rect 14657 10557 14691 10591
rect 14691 10557 14700 10591
rect 14648 10548 14700 10557
rect 14832 10548 14884 10600
rect 20352 10548 20404 10600
rect 23204 10752 23256 10804
rect 23848 10752 23900 10804
rect 24032 10684 24084 10736
rect 23296 10616 23348 10668
rect 21088 10548 21140 10600
rect 23572 10548 23624 10600
rect 24308 10591 24360 10600
rect 24308 10557 24317 10591
rect 24317 10557 24351 10591
rect 24351 10557 24360 10591
rect 24308 10548 24360 10557
rect 24400 10591 24452 10600
rect 24400 10557 24409 10591
rect 24409 10557 24443 10591
rect 24443 10557 24452 10591
rect 24400 10548 24452 10557
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 10876 10455 10928 10464
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 12348 10412 12400 10464
rect 13084 10523 13136 10532
rect 13084 10489 13102 10523
rect 13102 10489 13136 10523
rect 13084 10480 13136 10489
rect 15660 10480 15712 10532
rect 16304 10480 16356 10532
rect 18420 10480 18472 10532
rect 20444 10523 20496 10532
rect 20444 10489 20453 10523
rect 20453 10489 20487 10523
rect 20487 10489 20496 10523
rect 20444 10480 20496 10489
rect 22284 10523 22336 10532
rect 15200 10412 15252 10464
rect 16856 10412 16908 10464
rect 21916 10455 21968 10464
rect 21916 10421 21925 10455
rect 21925 10421 21959 10455
rect 21959 10421 21968 10455
rect 21916 10412 21968 10421
rect 22284 10489 22318 10523
rect 22318 10489 22336 10523
rect 22284 10480 22336 10489
rect 25412 10412 25464 10464
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 9220 10208 9272 10260
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 10048 10208 10100 10260
rect 10508 10208 10560 10260
rect 10600 10208 10652 10260
rect 10784 10208 10836 10260
rect 11152 10208 11204 10260
rect 13360 10208 13412 10260
rect 14464 10208 14516 10260
rect 15384 10208 15436 10260
rect 16764 10208 16816 10260
rect 18788 10208 18840 10260
rect 24308 10208 24360 10260
rect 24400 10208 24452 10260
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 10140 10072 10192 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 10416 10115 10468 10124
rect 10416 10081 10425 10115
rect 10425 10081 10459 10115
rect 10459 10081 10468 10115
rect 10416 10072 10468 10081
rect 10692 10072 10744 10124
rect 12624 10140 12676 10192
rect 16304 10140 16356 10192
rect 20076 10140 20128 10192
rect 21916 10140 21968 10192
rect 22192 10140 22244 10192
rect 10876 10072 10928 10124
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 12256 10115 12308 10124
rect 12256 10081 12265 10115
rect 12265 10081 12299 10115
rect 12299 10081 12308 10115
rect 12256 10072 12308 10081
rect 13820 10072 13872 10124
rect 16212 10115 16264 10124
rect 16212 10081 16221 10115
rect 16221 10081 16255 10115
rect 16255 10081 16264 10115
rect 16212 10072 16264 10081
rect 19524 10072 19576 10124
rect 20168 10072 20220 10124
rect 20720 10072 20772 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 21364 10072 21416 10124
rect 10232 9936 10284 9988
rect 10692 9936 10744 9988
rect 11704 9936 11756 9988
rect 25688 10004 25740 10056
rect 20812 9936 20864 9988
rect 24308 9936 24360 9988
rect 25596 9936 25648 9988
rect 10048 9868 10100 9920
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 12900 9868 12952 9920
rect 14924 9868 14976 9920
rect 22744 9911 22796 9920
rect 22744 9877 22753 9911
rect 22753 9877 22787 9911
rect 22787 9877 22796 9911
rect 22744 9868 22796 9877
rect 23940 9868 23992 9920
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 11152 9664 11204 9716
rect 9864 9596 9916 9648
rect 11244 9596 11296 9648
rect 13820 9664 13872 9716
rect 21364 9664 21416 9716
rect 23204 9707 23256 9716
rect 23204 9673 23213 9707
rect 23213 9673 23247 9707
rect 23247 9673 23256 9707
rect 23204 9664 23256 9673
rect 16396 9596 16448 9648
rect 10048 9460 10100 9512
rect 10416 9460 10468 9512
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 10968 9460 11020 9512
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 11704 9528 11756 9580
rect 11796 9460 11848 9512
rect 12532 9460 12584 9512
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 15108 9460 15160 9512
rect 19432 9596 19484 9648
rect 23480 9596 23532 9648
rect 13268 9392 13320 9444
rect 13728 9392 13780 9444
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 10140 9324 10192 9376
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 10508 9324 10560 9376
rect 11796 9324 11848 9376
rect 16212 9324 16264 9376
rect 17224 9392 17276 9444
rect 18604 9392 18656 9444
rect 20352 9460 20404 9512
rect 20720 9460 20772 9512
rect 22008 9460 22060 9512
rect 22192 9460 22244 9512
rect 19984 9392 20036 9444
rect 23480 9392 23532 9444
rect 24032 9460 24084 9512
rect 25504 9503 25556 9512
rect 25504 9469 25513 9503
rect 25513 9469 25547 9503
rect 25547 9469 25556 9503
rect 25504 9460 25556 9469
rect 25596 9503 25648 9512
rect 25596 9469 25605 9503
rect 25605 9469 25639 9503
rect 25639 9469 25648 9503
rect 25596 9460 25648 9469
rect 25688 9460 25740 9512
rect 24860 9392 24912 9444
rect 20168 9324 20220 9376
rect 22836 9324 22888 9376
rect 23756 9324 23808 9376
rect 25136 9324 25188 9376
rect 25688 9367 25740 9376
rect 25688 9333 25697 9367
rect 25697 9333 25731 9367
rect 25731 9333 25740 9367
rect 25688 9324 25740 9333
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 9772 9120 9824 9172
rect 10600 9120 10652 9172
rect 11060 9120 11112 9172
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 11060 8984 11112 9036
rect 10968 8916 11020 8968
rect 11336 8984 11388 9036
rect 15200 9120 15252 9172
rect 16212 9120 16264 9172
rect 12256 9052 12308 9104
rect 11244 8848 11296 8900
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 16396 9052 16448 9104
rect 17224 9120 17276 9172
rect 18880 9120 18932 9172
rect 20352 9120 20404 9172
rect 23664 9120 23716 9172
rect 24032 9120 24084 9172
rect 24860 9120 24912 9172
rect 18972 8984 19024 9036
rect 22928 9052 22980 9104
rect 28172 9052 28224 9104
rect 19524 8984 19576 9036
rect 23112 9027 23164 9036
rect 23112 8993 23121 9027
rect 23121 8993 23155 9027
rect 23155 8993 23164 9027
rect 23112 8984 23164 8993
rect 23204 8984 23256 9036
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 25412 8984 25464 9036
rect 23020 8916 23072 8968
rect 28264 8916 28316 8968
rect 18880 8848 18932 8900
rect 21916 8848 21968 8900
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 12808 8780 12860 8832
rect 16212 8780 16264 8832
rect 17592 8780 17644 8832
rect 17776 8780 17828 8832
rect 20996 8823 21048 8832
rect 20996 8789 21005 8823
rect 21005 8789 21039 8823
rect 21039 8789 21048 8823
rect 20996 8780 21048 8789
rect 23388 8780 23440 8832
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 10324 8576 10376 8628
rect 10692 8576 10744 8628
rect 11428 8576 11480 8628
rect 13360 8576 13412 8628
rect 13728 8576 13780 8628
rect 13912 8576 13964 8628
rect 10600 8440 10652 8492
rect 15292 8576 15344 8628
rect 16304 8576 16356 8628
rect 19524 8576 19576 8628
rect 20720 8576 20772 8628
rect 22928 8576 22980 8628
rect 23020 8619 23072 8628
rect 23020 8585 23029 8619
rect 23029 8585 23063 8619
rect 23063 8585 23072 8619
rect 23020 8576 23072 8585
rect 11152 8440 11204 8492
rect 12348 8440 12400 8492
rect 16856 8508 16908 8560
rect 31668 8576 31720 8628
rect 13636 8372 13688 8424
rect 15476 8440 15528 8492
rect 21640 8440 21692 8492
rect 9680 8279 9732 8288
rect 9680 8245 9689 8279
rect 9689 8245 9723 8279
rect 9723 8245 9732 8279
rect 9680 8236 9732 8245
rect 11244 8304 11296 8356
rect 11980 8236 12032 8288
rect 13728 8236 13780 8288
rect 14924 8347 14976 8356
rect 14924 8313 14942 8347
rect 14942 8313 14976 8347
rect 14924 8304 14976 8313
rect 15108 8304 15160 8356
rect 23296 8372 23348 8424
rect 15292 8347 15344 8356
rect 15292 8313 15301 8347
rect 15301 8313 15335 8347
rect 15335 8313 15344 8347
rect 15292 8304 15344 8313
rect 16212 8304 16264 8356
rect 22652 8304 22704 8356
rect 23664 8372 23716 8424
rect 25504 8372 25556 8424
rect 18880 8236 18932 8288
rect 20168 8236 20220 8288
rect 23112 8236 23164 8288
rect 23940 8304 23992 8356
rect 24124 8347 24176 8356
rect 24124 8313 24136 8347
rect 24136 8313 24176 8347
rect 24124 8304 24176 8313
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 25688 8279 25740 8288
rect 25688 8245 25697 8279
rect 25697 8245 25731 8279
rect 25731 8245 25740 8279
rect 25688 8236 25740 8245
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 10048 8032 10100 8084
rect 11060 8032 11112 8084
rect 11244 8032 11296 8084
rect 10416 7828 10468 7880
rect 10600 7896 10652 7948
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 13636 8075 13688 8084
rect 13636 8041 13645 8075
rect 13645 8041 13679 8075
rect 13679 8041 13688 8075
rect 13636 8032 13688 8041
rect 13820 8032 13872 8084
rect 16856 8032 16908 8084
rect 17040 8032 17092 8084
rect 17500 8032 17552 8084
rect 20444 8032 20496 8084
rect 22652 8032 22704 8084
rect 23204 8032 23256 8084
rect 21180 7964 21232 8016
rect 11704 7803 11756 7812
rect 11704 7769 11713 7803
rect 11713 7769 11747 7803
rect 11747 7769 11756 7803
rect 11704 7760 11756 7769
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 12072 7896 12124 7948
rect 14004 7896 14056 7948
rect 15384 7896 15436 7948
rect 16304 7896 16356 7948
rect 17132 7939 17184 7948
rect 17132 7905 17141 7939
rect 17141 7905 17175 7939
rect 17175 7905 17184 7939
rect 17132 7896 17184 7905
rect 17224 7939 17276 7948
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 17408 7896 17460 7948
rect 18144 7896 18196 7948
rect 17040 7828 17092 7880
rect 17500 7828 17552 7880
rect 22100 7896 22152 7948
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 11612 7692 11664 7744
rect 12900 7760 12952 7812
rect 20628 7760 20680 7812
rect 14648 7692 14700 7744
rect 16580 7692 16632 7744
rect 16672 7692 16724 7744
rect 23204 7692 23256 7744
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 10416 7488 10468 7540
rect 10508 7488 10560 7540
rect 28448 7488 28500 7540
rect 16856 7420 16908 7472
rect 19248 7420 19300 7472
rect 21180 7420 21232 7472
rect 10968 7284 11020 7336
rect 12624 7284 12676 7336
rect 13728 7284 13780 7336
rect 14924 7284 14976 7336
rect 24032 7352 24084 7404
rect 18512 7327 18564 7336
rect 18512 7293 18521 7327
rect 18521 7293 18555 7327
rect 18555 7293 18564 7327
rect 18512 7284 18564 7293
rect 20536 7284 20588 7336
rect 11428 7148 11480 7200
rect 11888 7216 11940 7268
rect 14004 7216 14056 7268
rect 18236 7216 18288 7268
rect 13268 7148 13320 7200
rect 13636 7148 13688 7200
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 15384 7148 15436 7200
rect 18972 7148 19024 7200
rect 19616 7216 19668 7268
rect 20260 7216 20312 7268
rect 22376 7216 22428 7268
rect 23020 7216 23072 7268
rect 20352 7148 20404 7200
rect 22192 7148 22244 7200
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 22376 6987 22428 6996
rect 22376 6953 22385 6987
rect 22385 6953 22419 6987
rect 22419 6953 22428 6987
rect 22376 6944 22428 6953
rect 23020 6987 23072 6996
rect 23020 6953 23029 6987
rect 23029 6953 23063 6987
rect 23063 6953 23072 6987
rect 23020 6944 23072 6953
rect 11428 6851 11480 6860
rect 11428 6817 11437 6851
rect 11437 6817 11471 6851
rect 11471 6817 11480 6851
rect 11428 6808 11480 6817
rect 11796 6808 11848 6860
rect 12348 6851 12400 6860
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 12440 6740 12492 6792
rect 16120 6851 16172 6860
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 19248 6876 19300 6928
rect 20628 6876 20680 6928
rect 22192 6919 22244 6928
rect 22192 6885 22201 6919
rect 22201 6885 22235 6919
rect 22235 6885 22244 6919
rect 22192 6876 22244 6885
rect 18052 6808 18104 6860
rect 18512 6808 18564 6860
rect 19156 6808 19208 6860
rect 19616 6672 19668 6724
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 21824 6740 21876 6792
rect 22744 6808 22796 6860
rect 23388 6808 23440 6860
rect 28264 6740 28316 6792
rect 21548 6672 21600 6724
rect 23848 6672 23900 6724
rect 13544 6604 13596 6656
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 17868 6604 17920 6656
rect 19248 6604 19300 6656
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 20812 6604 20864 6656
rect 22008 6604 22060 6656
rect 22192 6604 22244 6656
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 12440 6400 12492 6452
rect 18236 6400 18288 6452
rect 18788 6443 18840 6452
rect 18788 6409 18797 6443
rect 18797 6409 18831 6443
rect 18831 6409 18840 6443
rect 18788 6400 18840 6409
rect 19524 6400 19576 6452
rect 21824 6443 21876 6452
rect 21824 6409 21833 6443
rect 21833 6409 21867 6443
rect 21867 6409 21876 6443
rect 21824 6400 21876 6409
rect 22100 6443 22152 6452
rect 22100 6409 22109 6443
rect 22109 6409 22143 6443
rect 22143 6409 22152 6443
rect 22100 6400 22152 6409
rect 17960 6332 18012 6384
rect 12532 6196 12584 6248
rect 12348 6128 12400 6180
rect 15384 6239 15436 6248
rect 15384 6205 15393 6239
rect 15393 6205 15427 6239
rect 15427 6205 15436 6239
rect 15384 6196 15436 6205
rect 15476 6239 15528 6248
rect 15476 6205 15485 6239
rect 15485 6205 15519 6239
rect 15519 6205 15528 6239
rect 15476 6196 15528 6205
rect 14556 6128 14608 6180
rect 17776 6239 17828 6248
rect 17776 6205 17785 6239
rect 17785 6205 17819 6239
rect 17819 6205 17828 6239
rect 17776 6196 17828 6205
rect 18328 6239 18380 6248
rect 18328 6205 18337 6239
rect 18337 6205 18371 6239
rect 18371 6205 18380 6239
rect 18328 6196 18380 6205
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 19892 6264 19944 6316
rect 21548 6264 21600 6316
rect 19800 6239 19852 6248
rect 19800 6205 19809 6239
rect 19809 6205 19843 6239
rect 19843 6205 19852 6239
rect 19800 6196 19852 6205
rect 21732 6239 21784 6248
rect 21732 6205 21741 6239
rect 21741 6205 21775 6239
rect 21775 6205 21784 6239
rect 21732 6196 21784 6205
rect 25688 6264 25740 6316
rect 22192 6239 22244 6248
rect 22192 6205 22201 6239
rect 22201 6205 22235 6239
rect 22235 6205 22244 6239
rect 22192 6196 22244 6205
rect 16212 6128 16264 6180
rect 19340 6128 19392 6180
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 18696 6060 18748 6112
rect 19248 6103 19300 6112
rect 19248 6069 19257 6103
rect 19257 6069 19291 6103
rect 19291 6069 19300 6103
rect 19248 6060 19300 6069
rect 21088 6060 21140 6112
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 22008 6060 22060 6112
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 11428 5856 11480 5908
rect 12348 5899 12400 5908
rect 12348 5865 12357 5899
rect 12357 5865 12391 5899
rect 12391 5865 12400 5899
rect 12348 5856 12400 5865
rect 12900 5899 12952 5908
rect 12900 5865 12909 5899
rect 12909 5865 12943 5899
rect 12943 5865 12952 5899
rect 12900 5856 12952 5865
rect 15568 5856 15620 5908
rect 11796 5788 11848 5840
rect 11520 5720 11572 5772
rect 15660 5788 15712 5840
rect 13912 5763 13964 5772
rect 13912 5729 13921 5763
rect 13921 5729 13955 5763
rect 13955 5729 13964 5763
rect 13912 5720 13964 5729
rect 15568 5720 15620 5772
rect 19156 5856 19208 5908
rect 19432 5856 19484 5908
rect 20168 5856 20220 5908
rect 20720 5856 20772 5908
rect 20812 5856 20864 5908
rect 17040 5788 17092 5840
rect 19064 5763 19116 5772
rect 19064 5729 19073 5763
rect 19073 5729 19107 5763
rect 19107 5729 19116 5763
rect 19064 5720 19116 5729
rect 19892 5788 19944 5840
rect 22376 5856 22428 5908
rect 19616 5763 19668 5772
rect 19616 5729 19625 5763
rect 19625 5729 19659 5763
rect 19659 5729 19668 5763
rect 19616 5720 19668 5729
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 19984 5720 20036 5772
rect 20536 5720 20588 5772
rect 20628 5763 20680 5772
rect 20628 5729 20637 5763
rect 20637 5729 20671 5763
rect 20671 5729 20680 5763
rect 20628 5720 20680 5729
rect 22008 5788 22060 5840
rect 23204 5652 23256 5704
rect 19248 5584 19300 5636
rect 14188 5516 14240 5568
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 15660 5516 15712 5568
rect 16396 5516 16448 5568
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 20536 5559 20588 5568
rect 20536 5525 20545 5559
rect 20545 5525 20579 5559
rect 20579 5525 20588 5559
rect 20536 5516 20588 5525
rect 24124 5584 24176 5636
rect 22560 5516 22612 5568
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 13912 5312 13964 5364
rect 16212 5312 16264 5364
rect 16304 5312 16356 5364
rect 17132 5312 17184 5364
rect 18144 5312 18196 5364
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 18604 5312 18656 5364
rect 20628 5312 20680 5364
rect 22008 5355 22060 5364
rect 22008 5321 22017 5355
rect 22017 5321 22051 5355
rect 22051 5321 22060 5355
rect 22008 5312 22060 5321
rect 14280 5176 14332 5228
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 14648 5108 14700 5160
rect 15568 5108 15620 5160
rect 17500 5176 17552 5228
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 19156 5244 19208 5296
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 18420 5151 18472 5160
rect 18420 5117 18429 5151
rect 18429 5117 18463 5151
rect 18463 5117 18472 5151
rect 18420 5108 18472 5117
rect 20444 5151 20496 5160
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 21180 5108 21232 5160
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 14372 4972 14424 4981
rect 15476 4972 15528 5024
rect 15752 4972 15804 5024
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 14280 4768 14332 4820
rect 14372 4768 14424 4820
rect 15660 4768 15712 4820
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 18604 4768 18656 4820
rect 19340 4768 19392 4820
rect 20260 4700 20312 4752
rect 20536 4632 20588 4684
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 9680 3544 9732 3596
rect 14096 3544 14148 3596
rect 10968 3476 11020 3528
rect 13820 3476 13872 3528
rect 10232 3408 10284 3460
rect 23204 3408 23256 3460
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 19340 2796 19392 2848
rect 20996 2796 21048 2848
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
rect 16028 416 16080 468
rect 16396 416 16448 468
<< metal2 >>
rect 13542 19600 13598 20000
rect 14186 19600 14242 20000
rect 14830 19600 14886 20000
rect 15474 19600 15530 20000
rect 16762 19600 16818 20000
rect 17052 19638 17356 19666
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 13556 18970 13584 19600
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 4250 18459 4558 18468
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 4250 15260 4558 15269
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 13464 12866 13492 18566
rect 13464 12838 13676 12866
rect 13464 12782 13492 12838
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 9600 11354 9628 12242
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9404 11212 9456 11218
rect 9692 11200 9720 11766
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9404 11154 9456 11160
rect 9600 11172 9720 11200
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 9416 10606 9444 11154
rect 9600 10606 9628 11172
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 8102 10299 8410 10308
rect 9232 10266 9260 10406
rect 9324 10266 9352 10542
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9692 10130 9720 11018
rect 9784 10810 9812 11698
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9876 11354 9904 11562
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9968 11218 9996 12038
rect 11072 11898 11100 12242
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 11898 11284 12174
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 11354 10180 11494
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10130 9812 10406
rect 9876 10198 9904 11086
rect 10060 10266 10088 11154
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 10152 10130 10180 10950
rect 10244 10810 10272 11630
rect 11440 11354 11468 11630
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10336 10606 10364 10950
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10428 10282 10456 11154
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10244 10254 10456 10282
rect 10520 10266 10548 10542
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10266 10640 10406
rect 10508 10260 10560 10266
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10060 9926 10088 10066
rect 10244 9994 10272 10254
rect 10508 10202 10560 10208
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10414 10160 10470 10169
rect 10324 10124 10376 10130
rect 10704 10130 10732 10610
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10796 10266 10824 10542
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10888 10130 10916 10406
rect 11164 10266 11192 10406
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11348 10130 11376 10950
rect 11440 10810 11468 11290
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10606 11560 12310
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11624 11694 11652 12106
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11898 11836 12038
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12268 11354 12296 11494
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11955 10843 12263 10852
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 12268 10130 12296 10610
rect 12360 10606 12388 12650
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12452 11898 12480 12242
rect 12728 11898 12756 12242
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12544 11558 12572 11630
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12912 11014 12940 12038
rect 13188 11830 13216 12582
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13280 11626 13308 12242
rect 13556 11898 13584 12718
rect 13648 12442 13676 12838
rect 14200 12782 14228 19600
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13832 12374 13860 12582
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13832 11830 13860 12038
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13924 11694 13952 12582
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13556 11354 13584 11630
rect 13648 11354 13676 11630
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 14016 11218 14044 12038
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14108 11558 14136 11834
rect 14200 11694 14228 12718
rect 14476 11898 14504 12786
rect 14660 12102 14688 13262
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14660 11830 14688 12038
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 10414 10095 10416 10104
rect 10324 10066 10376 10072
rect 10468 10095 10470 10104
rect 10692 10124 10744 10130
rect 10416 10066 10468 10072
rect 10692 10066 10744 10072
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 9784 9178 9812 9318
rect 9876 9217 9904 9590
rect 10060 9518 10088 9862
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10138 9616 10194 9625
rect 10138 9551 10194 9560
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10152 9382 10180 9551
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9862 9208 9918 9217
rect 9772 9172 9824 9178
rect 9862 9143 9918 9152
rect 9772 9114 9824 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 9692 8129 9720 8230
rect 9678 8120 9734 8129
rect 10060 8090 10088 8978
rect 9678 8055 9734 8064
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 9692 400 9720 3538
rect 10244 3466 10272 9658
rect 10336 8634 10364 10066
rect 10704 9994 10732 10066
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9518 10732 9930
rect 11164 9722 11192 10066
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11244 9648 11296 9654
rect 11242 9616 11244 9625
rect 11296 9616 11298 9625
rect 11242 9551 11298 9560
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10428 9382 10456 9454
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10520 7970 10548 9318
rect 10612 9178 10640 9454
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10980 8974 11008 9454
rect 11072 9178 11100 9454
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11060 9036 11112 9042
rect 11336 9036 11388 9042
rect 11112 8996 11192 9024
rect 11060 8978 11112 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8634 10732 8774
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10336 7942 10548 7970
rect 10612 7954 10640 8434
rect 10600 7948 10652 7954
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 10336 400 10364 7942
rect 10600 7890 10652 7896
rect 10416 7880 10468 7886
rect 10468 7828 10548 7834
rect 10416 7822 10548 7828
rect 10428 7806 10548 7822
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7546 10456 7686
rect 10520 7546 10548 7806
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10980 7342 11008 8910
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8090 11100 8774
rect 11164 8498 11192 8996
rect 11256 8996 11336 9024
rect 11256 8906 11284 8996
rect 11336 8978 11388 8984
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11256 8362 11284 8842
rect 11440 8634 11468 10066
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11716 9586 11744 9930
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11808 9518 11836 9862
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11256 8242 11284 8298
rect 11164 8214 11284 8242
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 7970 11192 8214
rect 11440 8106 11468 8570
rect 11256 8090 11468 8106
rect 11244 8084 11468 8090
rect 11296 8078 11468 8084
rect 11244 8026 11296 8032
rect 11808 7970 11836 9318
rect 12360 9194 12388 10406
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12268 9166 12388 9194
rect 12438 9208 12494 9217
rect 12268 9110 12296 9166
rect 12544 9194 12572 9454
rect 12494 9166 12572 9194
rect 12438 9143 12494 9152
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12544 9042 12572 9166
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11164 7954 11284 7970
rect 11164 7948 11296 7954
rect 11164 7942 11244 7948
rect 11808 7942 11928 7970
rect 11992 7954 12020 8230
rect 12070 8120 12126 8129
rect 12070 8055 12126 8064
rect 12084 7954 12112 8055
rect 11244 7890 11296 7896
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 7018 11468 7142
rect 11440 6990 11560 7018
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11440 5914 11468 6802
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11532 5778 11560 6990
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10980 400 11008 3470
rect 11624 400 11652 7686
rect 11716 2774 11744 7754
rect 11900 7698 11928 7942
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11808 7670 11928 7698
rect 11808 6866 11836 7670
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11900 6746 11928 7210
rect 12360 6866 12388 8434
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 11808 6718 11928 6746
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 11808 5846 11836 6718
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11955 6491 12263 6500
rect 12452 6458 12480 6734
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12544 6254 12572 8978
rect 12636 7342 12664 10134
rect 12912 9926 12940 10950
rect 13648 10674 13676 10950
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 10169 13124 10474
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13082 10160 13138 10169
rect 13082 10095 13138 10104
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12360 5914 12388 6122
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 12820 3482 12848 8774
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12912 5914 12940 7754
rect 13280 7206 13308 9386
rect 13372 8634 13400 10202
rect 13648 9518 13676 10610
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13832 9722 13860 10066
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 8634 13768 9386
rect 13924 8634 13952 11154
rect 14108 10742 14136 11494
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14292 10810 14320 11154
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14384 8922 14412 11086
rect 14476 10266 14504 11222
rect 14568 11150 14596 11494
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14660 10606 14688 11766
rect 14844 10606 14872 19600
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15212 12850 15240 13806
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13258 15332 13670
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15488 12434 15516 19600
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12866 15792 13126
rect 15396 12406 15516 12434
rect 15672 12838 15792 12866
rect 16212 12844 16264 12850
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15028 11354 15056 11562
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15396 10674 15424 12406
rect 15672 12306 15700 12838
rect 16212 12786 16264 12792
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 16224 12306 16252 12786
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15764 11694 15792 11834
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 16684 11558 16712 13262
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 15807 11452 16115 11461
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15807 11387 16115 11396
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 16132 10554 16160 10950
rect 15660 10532 15712 10538
rect 16132 10526 16252 10554
rect 15660 10474 15712 10480
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14384 8894 14872 8922
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13648 8090 13676 8366
rect 13728 8288 13780 8294
rect 13780 8236 13860 8242
rect 13728 8230 13860 8236
rect 13740 8214 13860 8230
rect 13832 8090 13860 8214
rect 13636 8084 13688 8090
rect 13820 8084 13872 8090
rect 13688 8044 13768 8072
rect 13636 8026 13688 8032
rect 13740 7342 13768 8044
rect 13820 8026 13872 8032
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 14016 7274 14044 7890
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 13648 7002 13676 7142
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12820 3454 12940 3482
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 11716 2746 11836 2774
rect 9678 0 9734 400
rect 10322 0 10378 400
rect 10966 0 11022 400
rect 11610 0 11666 400
rect 11808 354 11836 2746
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 12176 462 12296 490
rect 12176 354 12204 462
rect 12268 400 12296 462
rect 12912 400 12940 3454
rect 13556 400 13584 6598
rect 13832 3534 13860 7142
rect 14200 6914 14228 7142
rect 14108 6886 14228 6914
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13924 5370 13952 5714
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 14108 3602 14136 6886
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 14200 400 14228 5510
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14292 4826 14320 5170
rect 14476 5166 14504 5510
rect 14568 5234 14596 6122
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14660 5166 14688 7686
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14384 4826 14412 4966
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14844 400 14872 8894
rect 14936 8362 14964 9862
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 8362 15148 9454
rect 15212 9178 15240 10406
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15304 8362 15332 8570
rect 15396 8514 15424 10202
rect 15396 8498 15516 8514
rect 15396 8492 15528 8498
rect 15396 8486 15476 8492
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 14936 7342 14964 8298
rect 15396 7954 15424 8486
rect 15476 8434 15528 8440
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 6254 15424 7142
rect 15672 6662 15700 10474
rect 15807 10364 16115 10373
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 16224 10130 16252 10526
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 16316 10198 16344 10474
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 16224 9178 16252 9318
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8362 16252 8774
rect 16316 8634 16344 10134
rect 16408 9654 16436 11290
rect 16776 10266 16804 19600
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16960 11830 16988 12718
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16408 9110 16436 9590
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16868 8566 16896 10406
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15807 8123 16115 8132
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 16224 6882 16252 8298
rect 17052 8090 17080 19638
rect 17328 19530 17356 19638
rect 17406 19600 17462 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 19338 19600 19394 20000
rect 19982 19600 20038 20000
rect 20626 19600 20682 20000
rect 17420 19530 17448 19600
rect 17328 19502 17448 19530
rect 18064 14362 18092 19600
rect 18708 16046 18736 19600
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18064 14334 18276 14362
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 13870 18184 14214
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17696 11898 17724 12650
rect 17972 12646 18000 13194
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17972 11694 18000 12582
rect 18064 11694 18092 13670
rect 18156 13462 18184 13670
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 18248 12434 18276 14334
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18340 13394 18368 13738
rect 18328 13388 18380 13394
rect 18328 13330 18380 13336
rect 18156 12406 18276 12434
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16132 6866 16252 6882
rect 16120 6860 16252 6866
rect 16172 6854 16252 6860
rect 16120 6802 16172 6808
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5250 15516 6190
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5914 15608 6054
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15672 5846 15700 6598
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15580 5386 15608 5714
rect 15660 5568 15712 5574
rect 15712 5516 15792 5534
rect 15660 5510 15792 5516
rect 15672 5506 15792 5510
rect 15580 5358 15700 5386
rect 15488 5222 15608 5250
rect 15580 5166 15608 5222
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 400 15516 4966
rect 15672 4826 15700 5358
rect 15764 5030 15792 5506
rect 16224 5370 16252 6122
rect 16316 5370 16344 7890
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 16408 474 16436 5510
rect 16592 2802 16620 7686
rect 16684 5166 16712 7686
rect 16868 7478 16896 8026
rect 17144 7954 17172 11494
rect 18156 11286 18184 12406
rect 18432 11694 18460 13942
rect 19352 13870 19380 19600
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 19996 15434 20024 19600
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 20640 15366 20668 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 31217 19068 31525 19077
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 18616 13394 18644 13738
rect 18696 13456 18748 13462
rect 18696 13398 18748 13404
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18340 11354 18368 11630
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18524 11286 18552 13126
rect 18708 11898 18736 13398
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18892 12442 18920 12786
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18788 12368 18840 12374
rect 18788 12310 18840 12316
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17236 9178 17264 9386
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17512 8090 17540 11154
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 17052 5846 17080 7822
rect 17236 6914 17264 7890
rect 17420 7002 17448 7890
rect 17512 7886 17540 8026
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17604 6914 17632 8774
rect 17144 6886 17264 6914
rect 17512 6886 17632 6914
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 17144 5370 17172 6886
rect 17512 5534 17540 6886
rect 17788 6254 17816 8774
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5534 17724 6054
rect 17420 5506 17540 5534
rect 17604 5506 17724 5534
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16592 2774 16804 2802
rect 16028 468 16080 474
rect 16396 468 16448 474
rect 16080 428 16160 456
rect 16028 410 16080 416
rect 16132 400 16160 428
rect 16396 410 16448 416
rect 16776 400 16804 2774
rect 17420 400 17448 5506
rect 17604 5386 17632 5506
rect 17880 5386 17908 6598
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17512 5358 17632 5386
rect 17696 5358 17908 5386
rect 17512 5234 17540 5358
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17696 5166 17724 5358
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17972 2802 18000 6326
rect 18064 4826 18092 6802
rect 18156 5370 18184 7890
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18248 6458 18276 7210
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18340 5370 18368 6190
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18432 5166 18460 10474
rect 18604 9444 18656 9450
rect 18524 9404 18604 9432
rect 18524 7342 18552 9404
rect 18604 9386 18656 9392
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18524 6866 18552 7278
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18708 6254 18736 11086
rect 18800 10266 18828 12310
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19076 11694 19104 12242
rect 19260 11694 19288 13126
rect 19444 12986 19472 13738
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19432 11620 19484 11626
rect 19432 11562 19484 11568
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18800 9674 18828 10202
rect 18800 9646 19104 9674
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18892 8906 18920 9114
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18892 6914 18920 8230
rect 18984 7206 19012 8978
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18800 6886 18920 6914
rect 18800 6458 18828 6886
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18616 4826 18644 5306
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 17972 2774 18092 2802
rect 18064 400 18092 2774
rect 18708 400 18736 6054
rect 19076 5778 19104 9646
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19260 6934 19288 7414
rect 19248 6928 19300 6934
rect 19352 6914 19380 11154
rect 19444 9654 19472 11562
rect 19536 10130 19564 13874
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 13462 19932 13670
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 20088 10198 20116 10950
rect 20364 10606 20392 12038
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20076 10192 20128 10198
rect 20076 10134 20128 10140
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19536 8634 19564 8978
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 19616 7268 19668 7274
rect 19616 7210 19668 7216
rect 19352 6886 19472 6914
rect 19248 6870 19300 6876
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19168 5914 19196 6802
rect 19260 6662 19288 6870
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19168 5302 19196 5850
rect 19260 5642 19288 6054
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19156 5296 19208 5302
rect 19156 5238 19208 5244
rect 19352 4826 19380 6122
rect 19444 5914 19472 6886
rect 19628 6730 19656 7210
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19536 6458 19564 6598
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19798 6352 19854 6361
rect 19798 6287 19854 6296
rect 19892 6316 19944 6322
rect 19812 6254 19840 6287
rect 19892 6258 19944 6264
rect 19800 6248 19852 6254
rect 19614 6216 19670 6225
rect 19800 6190 19852 6196
rect 19614 6151 19670 6160
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19628 5778 19656 6151
rect 19904 5846 19932 6258
rect 19892 5840 19944 5846
rect 19798 5808 19854 5817
rect 19616 5772 19668 5778
rect 19892 5782 19944 5788
rect 19996 5778 20024 9386
rect 20180 9382 20208 10066
rect 20364 9518 20392 10542
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20364 9178 20392 9454
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20180 5914 20208 8230
rect 20456 8090 20484 10474
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 19798 5743 19800 5752
rect 19616 5714 19668 5720
rect 19852 5743 19854 5752
rect 19984 5772 20036 5778
rect 19800 5714 19852 5720
rect 19984 5714 20036 5720
rect 20272 5658 20300 7210
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 19996 5630 20300 5658
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19352 400 19380 2790
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 19996 400 20024 5630
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 4758 20300 5510
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 11808 326 12204 354
rect 12254 0 12310 400
rect 12898 0 12954 400
rect 13542 0 13598 400
rect 14186 0 14242 400
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16118 0 16174 400
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 18050 0 18106 400
rect 18694 0 18750 400
rect 19338 0 19394 400
rect 19982 0 20038 400
rect 20364 354 20392 7142
rect 20456 5166 20484 8026
rect 20548 7342 20576 12106
rect 20640 12102 20668 13330
rect 20732 12374 20760 13942
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20732 9518 20760 10066
rect 20824 9994 20852 15982
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21468 12374 21496 13874
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21652 12442 21680 13806
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21836 12986 21864 13126
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 22204 12442 22232 15370
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 21180 11620 21232 11626
rect 21180 11562 21232 11568
rect 21100 10606 21128 11562
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20732 8634 20760 9454
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20640 6934 20668 7754
rect 20628 6928 20680 6934
rect 20628 6870 20680 6876
rect 20640 5778 20668 6870
rect 20732 5914 20760 8570
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 5914 20852 6598
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20548 5658 20576 5714
rect 20548 5630 20668 5658
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20548 4690 20576 5510
rect 20640 5370 20668 5630
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 21008 2854 21036 8774
rect 21192 8022 21220 11562
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 10198 21956 10406
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21192 7478 21220 7958
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21284 6914 21312 10066
rect 21376 9722 21404 10066
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 22020 9518 22048 11154
rect 22296 10538 22324 11630
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23216 10810 23244 11154
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22204 9518 22232 10134
rect 23202 10024 23258 10033
rect 23202 9959 23258 9968
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21192 6886 21312 6914
rect 21192 6118 21220 6886
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21560 6322 21588 6666
rect 21652 6610 21680 8434
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21652 6582 21772 6610
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21744 6254 21772 6582
rect 21836 6458 21864 6734
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21100 2802 21128 6054
rect 21192 5166 21220 6054
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21100 2774 21312 2802
rect 20548 462 20668 490
rect 20548 354 20576 462
rect 20640 400 20668 462
rect 21284 400 21312 2774
rect 21928 400 21956 8842
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22664 8090 22692 8298
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22006 6760 22062 6769
rect 22006 6695 22062 6704
rect 22020 6662 22048 6695
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 22112 6458 22140 7890
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22204 6934 22232 7142
rect 22388 7002 22416 7210
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22756 6866 22784 9862
rect 23216 9722 23244 9959
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22848 9081 22876 9318
rect 22928 9104 22980 9110
rect 22834 9072 22890 9081
rect 22928 9046 22980 9052
rect 22834 9007 22890 9016
rect 22940 8634 22968 9046
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23204 9036 23256 9042
rect 23204 8978 23256 8984
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23032 8634 23060 8910
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 23124 8294 23152 8978
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 23216 8090 23244 8978
rect 23308 8430 23336 10610
rect 23584 10606 23612 11086
rect 23860 10810 23888 14282
rect 24228 11762 24256 15302
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 31217 13628 31525 13637
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 28446 12336 28502 12345
rect 28446 12271 28502 12280
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 28262 11656 28318 11665
rect 24032 11620 24084 11626
rect 28262 11591 28318 11600
rect 24032 11562 24084 11568
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 24044 10742 24072 11562
rect 28276 11354 28304 11591
rect 28264 11348 28316 11354
rect 28264 11290 28316 11296
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 24032 10736 24084 10742
rect 24032 10678 24084 10684
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 24320 10266 24348 10542
rect 24412 10266 24440 10542
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24400 10260 24452 10266
rect 24400 10202 24452 10208
rect 24320 9994 24348 10202
rect 24308 9988 24360 9994
rect 24308 9930 24360 9936
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23492 9450 23520 9590
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 23768 9438 23888 9466
rect 23768 9382 23796 9438
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23020 7268 23072 7274
rect 23020 7210 23072 7216
rect 23032 7002 23060 7210
rect 23020 6996 23072 7002
rect 23020 6938 23072 6944
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22204 6254 22232 6598
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 5846 22048 6054
rect 22388 5914 22416 6802
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 22020 5370 22048 5782
rect 23216 5710 23244 7686
rect 23400 6866 23428 8774
rect 23676 8430 23704 9114
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23860 6730 23888 9438
rect 23952 8362 23980 9862
rect 24032 9512 24084 9518
rect 24032 9454 24084 9460
rect 24044 9178 24072 9454
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24872 9178 24900 9386
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 24044 7410 24072 9114
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23848 6724 23900 6730
rect 23848 6666 23900 6672
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 24136 5642 24164 8298
rect 25148 6225 25176 9318
rect 25332 9042 25360 11018
rect 28354 10976 28410 10985
rect 27365 10908 27673 10917
rect 28354 10911 28410 10920
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25424 9042 25452 10406
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25608 9518 25636 9930
rect 25700 9518 25728 9998
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 28262 9616 28318 9625
rect 28262 9551 28318 9560
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25596 9512 25648 9518
rect 25596 9454 25648 9460
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25516 8430 25544 9454
rect 25688 9376 25740 9382
rect 25688 9318 25740 9324
rect 25504 8424 25556 8430
rect 25700 8378 25728 9318
rect 28172 9104 28224 9110
rect 28172 9046 28224 9052
rect 28184 8945 28212 9046
rect 28276 8974 28304 9551
rect 28368 9081 28396 10911
rect 28354 9072 28410 9081
rect 28354 9007 28410 9016
rect 28264 8968 28316 8974
rect 28170 8936 28226 8945
rect 28264 8910 28316 8916
rect 28170 8871 28226 8880
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 25504 8366 25556 8372
rect 25608 8350 25728 8378
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25424 6361 25452 8230
rect 25410 6352 25466 6361
rect 25410 6287 25466 6296
rect 25134 6216 25190 6225
rect 25134 6151 25190 6160
rect 25608 5817 25636 8350
rect 25688 8288 25740 8294
rect 25688 8230 25740 8236
rect 25700 6322 25728 8230
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 27365 7579 27673 7588
rect 28460 7546 28488 12271
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31666 10296 31722 10305
rect 31666 10231 31722 10240
rect 31680 10033 31708 10231
rect 31666 10024 31722 10033
rect 31666 9959 31722 9968
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 31217 9211 31525 9220
rect 31668 8628 31720 8634
rect 31668 8570 31720 8576
rect 31680 8265 31708 8570
rect 31666 8256 31722 8265
rect 31217 8188 31525 8197
rect 31666 8191 31722 8200
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 31217 8123 31525 8132
rect 28448 7540 28500 7546
rect 28448 7482 28500 7488
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 28262 6896 28318 6905
rect 28262 6831 28318 6840
rect 28276 6798 28304 6831
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 25594 5808 25650 5817
rect 25594 5743 25650 5752
rect 24124 5636 24176 5642
rect 24124 5578 24176 5584
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 22572 400 22600 5510
rect 27365 5468 27673 5477
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 23204 3460 23256 3466
rect 23204 3402 23256 3408
rect 23216 400 23244 3402
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 31217 2748 31525 2757
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 20364 326 20576 354
rect 20626 0 20682 400
rect 21270 0 21326 400
rect 21914 0 21970 400
rect 22558 0 22614 400
rect 23202 0 23258 400
<< via2 >>
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 10414 10124 10470 10160
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 10414 10104 10416 10124
rect 10416 10104 10468 10124
rect 10468 10104 10470 10124
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 10138 9560 10194 9616
rect 9862 9152 9918 9208
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 9678 8064 9734 8120
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 11242 9596 11244 9616
rect 11244 9596 11296 9616
rect 11296 9596 11298 9616
rect 11242 9560 11298 9596
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 12438 9152 12494 9208
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 12070 8064 12126 8120
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 13082 10104 13138 10160
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 19798 6296 19854 6352
rect 19614 6160 19670 6216
rect 19798 5772 19854 5808
rect 19798 5752 19800 5772
rect 19800 5752 19852 5772
rect 19852 5752 19854 5772
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 23202 9968 23258 10024
rect 22006 6704 22062 6760
rect 22834 9016 22890 9072
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 28446 12280 28502 12336
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 28262 11600 28318 11656
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 28354 10920 28410 10976
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 28262 9560 28318 9616
rect 28354 9016 28410 9072
rect 28170 8880 28226 8936
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 25410 6296 25466 6352
rect 25134 6160 25190 6216
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10240 31722 10296
rect 31666 9968 31722 10024
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 31666 8200 31722 8256
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 28262 6840 28318 6896
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 25594 5752 25650 5808
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
<< metal3 >>
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31213 19007 31529 19008
rect 4246 18528 4562 18529
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31213 13567 31529 13568
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 28441 12338 28507 12341
rect 31600 12338 32000 12368
rect 28441 12336 32000 12338
rect 28441 12280 28446 12336
rect 28502 12280 32000 12336
rect 28441 12278 32000 12280
rect 28441 12275 28507 12278
rect 31600 12248 32000 12278
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 28257 11658 28323 11661
rect 31600 11658 32000 11688
rect 28257 11656 32000 11658
rect 28257 11600 28262 11656
rect 28318 11600 32000 11656
rect 28257 11598 32000 11600
rect 28257 11595 28323 11598
rect 31600 11568 32000 11598
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 28349 10978 28415 10981
rect 31600 10978 32000 11008
rect 28349 10976 32000 10978
rect 28349 10920 28354 10976
rect 28410 10920 32000 10976
rect 28349 10918 32000 10920
rect 28349 10915 28415 10918
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 31600 10888 32000 10918
rect 27361 10847 27677 10848
rect 8098 10368 8414 10369
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 10409 10162 10475 10165
rect 13077 10162 13143 10165
rect 10409 10160 13143 10162
rect 10409 10104 10414 10160
rect 10470 10104 13082 10160
rect 13138 10104 13143 10160
rect 10409 10102 13143 10104
rect 10409 10099 10475 10102
rect 13077 10099 13143 10102
rect 23197 10026 23263 10029
rect 31661 10026 31727 10029
rect 23197 10024 31727 10026
rect 23197 9968 23202 10024
rect 23258 9968 31666 10024
rect 31722 9968 31727 10024
rect 23197 9966 31727 9968
rect 23197 9963 23263 9966
rect 31661 9963 31727 9966
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 10133 9618 10199 9621
rect 11237 9618 11303 9621
rect 10133 9616 11303 9618
rect 10133 9560 10138 9616
rect 10194 9560 11242 9616
rect 11298 9560 11303 9616
rect 10133 9558 11303 9560
rect 10133 9555 10199 9558
rect 11237 9555 11303 9558
rect 28257 9618 28323 9621
rect 31600 9618 32000 9648
rect 28257 9616 32000 9618
rect 28257 9560 28262 9616
rect 28318 9560 32000 9616
rect 28257 9558 32000 9560
rect 28257 9555 28323 9558
rect 31600 9528 32000 9558
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 9857 9210 9923 9213
rect 12433 9210 12499 9213
rect 9857 9208 12499 9210
rect 9857 9152 9862 9208
rect 9918 9152 12438 9208
rect 12494 9152 12499 9208
rect 9857 9150 12499 9152
rect 9857 9147 9923 9150
rect 12433 9147 12499 9150
rect 22829 9074 22895 9077
rect 28349 9074 28415 9077
rect 22829 9072 28415 9074
rect 22829 9016 22834 9072
rect 22890 9016 28354 9072
rect 28410 9016 28415 9072
rect 22829 9014 28415 9016
rect 22829 9011 22895 9014
rect 28349 9011 28415 9014
rect 28165 8938 28231 8941
rect 31600 8938 32000 8968
rect 28165 8936 32000 8938
rect 28165 8880 28170 8936
rect 28226 8880 32000 8936
rect 28165 8878 32000 8880
rect 28165 8875 28231 8878
rect 31600 8848 32000 8878
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 31600 8256 32000 8288
rect 31600 8200 31666 8256
rect 31722 8200 32000 8256
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31600 8168 32000 8200
rect 31213 8127 31529 8128
rect 9673 8122 9739 8125
rect 12065 8122 12131 8125
rect 9673 8120 12131 8122
rect 9673 8064 9678 8120
rect 9734 8064 12070 8120
rect 12126 8064 12131 8120
rect 9673 8062 12131 8064
rect 9673 8059 9739 8062
rect 12065 8059 12131 8062
rect 4246 7648 4562 7649
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 31600 7578 32000 7608
rect 28214 7518 32000 7578
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 28214 7034 28274 7518
rect 31600 7488 32000 7518
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 24810 6974 28274 7034
rect 22001 6762 22067 6765
rect 24810 6762 24870 6974
rect 28257 6898 28323 6901
rect 31600 6898 32000 6928
rect 28257 6896 32000 6898
rect 28257 6840 28262 6896
rect 28318 6840 32000 6896
rect 28257 6838 32000 6840
rect 28257 6835 28323 6838
rect 31600 6808 32000 6838
rect 22001 6760 24870 6762
rect 22001 6704 22006 6760
rect 22062 6704 24870 6760
rect 22001 6702 24870 6704
rect 22001 6699 22067 6702
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 19793 6354 19859 6357
rect 25405 6354 25471 6357
rect 19793 6352 25471 6354
rect 19793 6296 19798 6352
rect 19854 6296 25410 6352
rect 25466 6296 25471 6352
rect 19793 6294 25471 6296
rect 19793 6291 19859 6294
rect 25405 6291 25471 6294
rect 19609 6218 19675 6221
rect 25129 6218 25195 6221
rect 19609 6216 25195 6218
rect 19609 6160 19614 6216
rect 19670 6160 25134 6216
rect 25190 6160 25195 6216
rect 19609 6158 25195 6160
rect 19609 6155 19675 6158
rect 25129 6155 25195 6158
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 19793 5810 19859 5813
rect 25589 5810 25655 5813
rect 19793 5808 25655 5810
rect 19793 5752 19798 5808
rect 19854 5752 25594 5808
rect 25650 5752 25655 5808
rect 19793 5750 25655 5752
rect 19793 5747 19859 5750
rect 25589 5747 25655 5750
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 27361 5407 27677 5408
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11949 12000 12269 13024
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 11949 8736 12269 9760
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 11949 6560 12269 7584
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 15801 15808 16121 16832
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 15801 10368 16121 11392
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15801 4928 16121 5952
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15801 3840 16121 4864
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19654 12000 19974 13024
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19654 7648 19974 8672
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 19654 4384 19974 5408
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 23506 15808 23826 16832
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
use sky130_fd_sc_hd__or2b_1  _10_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13524 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _11_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _12_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 16100 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _13__1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 20700 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__2
timestamp 1701704242
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__3
timestamp 1701704242
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__4
timestamp 1701704242
transform -1 0 11316 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__5
timestamp 1701704242
transform 1 0 13248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__6
timestamp 1701704242
transform -1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__7
timestamp 1701704242
transform -1 0 10856 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__8
timestamp 1701704242
transform -1 0 11776 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__9
timestamp 1701704242
transform 1 0 10672 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__10
timestamp 1701704242
transform -1 0 23736 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__11
timestamp 1701704242
transform -1 0 25576 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__12
timestamp 1701704242
transform 1 0 23644 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__15
timestamp 1701704242
transform -1 0 21160 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13_
timestamp 1701704242
transform 1 0 10120 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__13
timestamp 1701704242
transform 1 0 20700 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__14
timestamp 1701704242
transform 1 0 25576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _13__16
timestamp 1701704242
transform -1 0 20148 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _14_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13432 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _15_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _16_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14904 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _17_
timestamp 1701704242
transform 1 0 15548 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _18_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 19320 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _19_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15824 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _20_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18860 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _21_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18584 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _22_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 21252 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _23_
timestamp 1701704242
transform -1 0 20148 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _24_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16008 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _25_
timestamp 1701704242
transform 1 0 16652 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _26_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 20516 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _27_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14536 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _28_
timestamp 1701704242
transform -1 0 15272 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _29_
timestamp 1701704242
transform 1 0 13616 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _30_
timestamp 1701704242
transform 1 0 14536 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _31_
timestamp 1701704242
transform -1 0 13432 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _32_
timestamp 1701704242
transform -1 0 13432 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _33_
timestamp 1701704242
transform 1 0 14076 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _34_
timestamp 1701704242
transform 1 0 15732 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _35_
timestamp 1701704242
transform 1 0 17112 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _36_
timestamp 1701704242
transform 1 0 17940 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _37_
timestamp 1701704242
transform 1 0 19688 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _38_
timestamp 1701704242
transform -1 0 23552 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _39_
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _40_
timestamp 1701704242
transform -1 0 25300 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _41_
timestamp 1701704242
transform 1 0 20516 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _42_
timestamp 1701704242
transform 1 0 17112 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _43_
timestamp 1701704242
transform 1 0 16652 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _44_
timestamp 1701704242
transform 1 0 19412 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _45_
timestamp 1701704242
transform 1 0 21988 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _46_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 13432 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1701704242
transform -1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _48_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13984 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1701704242
transform -1 0 11592 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1701704242
transform 1 0 13616 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1701704242
transform 1 0 11960 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1701704242
transform -1 0 11960 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1701704242
transform -1 0 13984 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1701704242
transform 1 0 16652 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1701704242
transform -1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1701704242
transform -1 0 18400 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1701704242
transform -1 0 19504 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1701704242
transform -1 0 19872 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1701704242
transform -1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1701704242
transform -1 0 23276 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1701704242
transform -1 0 20148 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1701704242
transform -1 0 17204 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _63_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _64_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18768 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _65_
timestamp 1701704242
transform 1 0 23828 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _66_
timestamp 1701704242
transform 1 0 18768 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _67_
timestamp 1701704242
transform 1 0 21804 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _68_
timestamp 1701704242
transform 1 0 23092 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _69_
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _70_
timestamp 1701704242
transform -1 0 13524 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _71_
timestamp 1701704242
transform 1 0 16376 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _72_
timestamp 1701704242
transform 1 0 16100 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _73_
timestamp 1701704242
transform -1 0 12328 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _74_
timestamp 1701704242
transform -1 0 12328 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _75_
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _76_
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _77_
timestamp 1701704242
transform 1 0 20608 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _78_
timestamp 1701704242
transform 1 0 19228 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _79_
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _80_
timestamp 1701704242
transform -1 0 22356 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _81_
timestamp 1701704242
transform -1 0 22908 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _82_
timestamp 1701704242
transform -1 0 23460 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _83_
timestamp 1701704242
transform 1 0 22356 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _84_
timestamp 1701704242
transform 1 0 20332 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1701704242
transform -1 0 18584 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1701704242
transform -1 0 12328 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1701704242
transform 1 0 23092 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1701704242
transform -1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_stop pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18768 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[1\]
timestamp 1701704242
transform 1 0 15272 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[2\]
timestamp 1701704242
transform 1 0 14168 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[3\]
timestamp 1701704242
transform 1 0 12328 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[4\]
timestamp 1701704242
transform 1 0 12328 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[5\]
timestamp 1701704242
transform 1 0 14168 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[6\]
timestamp 1701704242
transform 1 0 16376 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[7\]
timestamp 1701704242
transform 1 0 17204 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[8\]
timestamp 1701704242
transform 1 0 19044 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[9\]
timestamp 1701704242
transform 1 0 19872 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[10\]
timestamp 1701704242
transform 1 0 21252 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[11\]
timestamp 1701704242
transform -1 0 22080 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[12\]
timestamp 1701704242
transform -1 0 22356 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[13\]
timestamp 1701704242
transform 1 0 19320 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[14\]
timestamp 1701704242
transform -1 0 20516 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_sig1_n_ana_\[15\]
timestamp 1701704242
transform -1 0 18308 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_dly_stop
timestamp 1701704242
transform 1 0 14168 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w_ring_ctr_clk
timestamp 1701704242
transform 1 0 17572 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_i_stop
timestamp 1701704242
transform -1 0 14168 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[1\]
timestamp 1701704242
transform -1 0 14168 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[2\]
timestamp 1701704242
transform -1 0 13432 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[3\]
timestamp 1701704242
transform -1 0 11592 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[4\]
timestamp 1701704242
transform -1 0 11592 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[5\]
timestamp 1701704242
transform -1 0 15824 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[6\]
timestamp 1701704242
transform -1 0 15456 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[7\]
timestamp 1701704242
transform 1 0 17204 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[8\]
timestamp 1701704242
transform -1 0 20516 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[9\]
timestamp 1701704242
transform 1 0 20516 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[10\]
timestamp 1701704242
transform -1 0 20516 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[11\]
timestamp 1701704242
transform 1 0 21160 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[12\]
timestamp 1701704242
transform -1 0 20332 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[13\]
timestamp 1701704242
transform -1 0 18492 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[14\]
timestamp 1701704242
transform -1 0 16928 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_dly_sig1_n_ana_\[15\]
timestamp 1701704242
transform -1 0 15824 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_w_ring_ctr_clk
timestamp 1701704242
transform -1 0 16652 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_i_stop
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[1\]
timestamp 1701704242
transform 1 0 16744 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[2\]
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[3\]
timestamp 1701704242
transform 1 0 14536 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[4\]
timestamp 1701704242
transform -1 0 13432 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[5\]
timestamp 1701704242
transform 1 0 14904 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[6\]
timestamp 1701704242
transform 1 0 18768 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[7\]
timestamp 1701704242
transform 1 0 16928 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[8\]
timestamp 1701704242
transform -1 0 20516 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[9\]
timestamp 1701704242
transform 1 0 21252 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[10\]
timestamp 1701704242
transform 1 0 23460 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[11\]
timestamp 1701704242
transform 1 0 23092 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[12\]
timestamp 1701704242
transform 1 0 23092 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[13\]
timestamp 1701704242
transform 1 0 21252 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[14\]
timestamp 1701704242
transform 1 0 19320 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_dly_sig1_n_ana_\[15\]
timestamp 1701704242
transform 1 0 18676 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_w_ring_ctr_clk
timestamp 1701704242
transform 1 0 20516 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_w_dly_stop
timestamp 1701704242
transform -1 0 13432 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_w_dly_stop
timestamp 1701704242
transform -1 0 12788 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_w_dly_stop
timestamp 1701704242
transform 1 0 14168 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_w_dly_stop
timestamp 1701704242
transform 1 0 20516 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__nor2_2  dly_stg01 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  dly_stg02
timestamp 1701704242
transform -1 0 13064 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  dly_stg03 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12512 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  dly_stg04
timestamp 1701704242
transform -1 0 12788 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  dly_stg09 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 18216 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_74
timestamp 1701704242
transform -1 0 12512 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_75
timestamp 1701704242
transform -1 0 14720 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_76
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_77
timestamp 1701704242
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_78
timestamp 1701704242
transform -1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_79
timestamp 1701704242
transform 1 0 15180 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_80
timestamp 1701704242
transform -1 0 14076 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  dly_stg11 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_73
timestamp 1701704242
transform 1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1701704242
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1701704242
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1701704242
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1701704242
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1701704242
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1701704242
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1701704242
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1701704242
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1701704242
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_329
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1701704242
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1701704242
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1701704242
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1701704242
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1701704242
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1701704242
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1701704242
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1701704242
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1701704242
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1701704242
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1701704242
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1701704242
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1701704242
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1701704242
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1701704242
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1701704242
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1701704242
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1701704242
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1701704242
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1701704242
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1701704242
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1701704242
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1701704242
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1701704242
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1701704242
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1701704242
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1701704242
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1701704242
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1701704242
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1701704242
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1701704242
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1701704242
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1701704242
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1701704242
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1701704242
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1701704242
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1701704242
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1701704242
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1701704242
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1701704242
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1701704242
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_329
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1701704242
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1701704242
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1701704242
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1701704242
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1701704242
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1701704242
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1701704242
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1701704242
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1701704242
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1701704242
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1701704242
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1701704242
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1701704242
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1701704242
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1701704242
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1701704242
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1701704242
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1701704242
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1701704242
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1701704242
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1701704242
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1701704242
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1701704242
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1701704242
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1701704242
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1701704242
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1701704242
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1701704242
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1701704242
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1701704242
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1701704242
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1701704242
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1701704242
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1701704242
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1701704242
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1701704242
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1701704242
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1701704242
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1701704242
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1701704242
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1701704242
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1701704242
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1701704242
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_329
timestamp 1701704242
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1701704242
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1701704242
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1701704242
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1701704242
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1701704242
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_137
timestamp 1701704242
transform 1 0 13156 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_145 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_163
timestamp 1701704242
transform 1 0 15548 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1701704242
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 1701704242
transform 1 0 17204 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_192
timestamp 1701704242
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_198
timestamp 1701704242
transform 1 0 18768 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_210
timestamp 1701704242
transform 1 0 19872 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1701704242
transform 1 0 20976 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1701704242
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1701704242
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1701704242
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1701704242
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1701704242
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1701704242
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1701704242
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_329
timestamp 1701704242
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1701704242
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1701704242
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1701704242
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1701704242
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1701704242
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1701704242
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1701704242
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1701704242
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_171
timestamp 1701704242
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_176
timestamp 1701704242
transform 1 0 16744 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_182
timestamp 1701704242
transform 1 0 17296 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1701704242
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_237
timestamp 1701704242
transform 1 0 22356 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 1701704242
transform 1 0 23460 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1701704242
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1701704242
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1701704242
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1701704242
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1701704242
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1701704242
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 1701704242
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_329
timestamp 1701704242
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1701704242
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1701704242
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1701704242
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1701704242
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1701704242
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1701704242
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_125
timestamp 1701704242
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_130
timestamp 1701704242
transform 1 0 12512 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_136
timestamp 1701704242
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_141
timestamp 1701704242
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1701704242
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_179
timestamp 1701704242
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1701704242
transform 1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_231
timestamp 1701704242
transform 1 0 21804 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_243
timestamp 1701704242
transform 1 0 22908 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_255
timestamp 1701704242
transform 1 0 24012 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_267
timestamp 1701704242
transform 1 0 25116 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1701704242
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1701704242
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1701704242
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1701704242
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1701704242
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_329
timestamp 1701704242
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1701704242
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1701704242
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1701704242
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1701704242
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1701704242
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1701704242
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1701704242
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_121
timestamp 1701704242
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_188
timestamp 1701704242
transform 1 0 17848 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1701704242
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_200
timestamp 1701704242
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_239
timestamp 1701704242
transform 1 0 22540 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1701704242
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1701704242
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1701704242
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1701704242
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1701704242
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1701704242
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1701704242
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_321
timestamp 1701704242
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 1701704242
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1701704242
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1701704242
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1701704242
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1701704242
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1701704242
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1701704242
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_246
timestamp 1701704242
transform 1 0 23184 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_258
timestamp 1701704242
transform 1 0 24288 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_270
timestamp 1701704242
transform 1 0 25392 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1701704242
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1701704242
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1701704242
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1701704242
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_329
timestamp 1701704242
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1701704242
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1701704242
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1701704242
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1701704242
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1701704242
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1701704242
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1701704242
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_97
timestamp 1701704242
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_213
timestamp 1701704242
transform 1 0 20148 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1701704242
transform 1 0 23552 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1701704242
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1701704242
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1701704242
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1701704242
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1701704242
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1701704242
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_321
timestamp 1701704242
transform 1 0 30084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_329
timestamp 1701704242
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1701704242
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1701704242
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1701704242
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1701704242
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1701704242
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1701704242
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_93
timestamp 1701704242
transform 1 0 9108 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_101
timestamp 1701704242
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_175
timestamp 1701704242
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_265
timestamp 1701704242
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1701704242
transform 1 0 26036 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1701704242
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1701704242
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1701704242
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_329
timestamp 1701704242
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1701704242
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1701704242
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1701704242
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1701704242
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1701704242
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_275
timestamp 1701704242
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_287
timestamp 1701704242
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_299
timestamp 1701704242
transform 1 0 28060 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1701704242
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1701704242
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_321
timestamp 1701704242
transform 1 0 30084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_329
timestamp 1701704242
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1701704242
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1701704242
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1701704242
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1701704242
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_93
timestamp 1701704242
transform 1 0 9108 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_101
timestamp 1701704242
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_272
timestamp 1701704242
transform 1 0 25576 0 -1 9248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1701704242
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1701704242
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1701704242
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1701704242
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_329
timestamp 1701704242
transform 1 0 30820 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1701704242
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1701704242
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1701704242
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1701704242
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1701704242
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_97
timestamp 1701704242
transform 1 0 9476 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_178
timestamp 1701704242
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_278
timestamp 1701704242
transform 1 0 26128 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_290
timestamp 1701704242
transform 1 0 27232 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_302
timestamp 1701704242
transform 1 0 28336 0 1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1701704242
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1701704242
transform 1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_329
timestamp 1701704242
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1701704242
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1701704242
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1701704242
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_81
timestamp 1701704242
transform 1 0 8004 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_89
timestamp 1701704242
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_268
timestamp 1701704242
transform 1 0 25208 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1701704242
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1701704242
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1701704242
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_329
timestamp 1701704242
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1701704242
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1701704242
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1701704242
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1701704242
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1701704242
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1701704242
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_262
timestamp 1701704242
transform 1 0 24656 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_274
timestamp 1701704242
transform 1 0 25760 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_286
timestamp 1701704242
transform 1 0 26864 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_298
timestamp 1701704242
transform 1 0 27968 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_306
timestamp 1701704242
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_321
timestamp 1701704242
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_329
timestamp 1701704242
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1701704242
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1701704242
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1701704242
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1701704242
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1701704242
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1701704242
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_93
timestamp 1701704242
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_133
timestamp 1701704242
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_141
timestamp 1701704242
transform 1 0 13524 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_151
timestamp 1701704242
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_176
timestamp 1701704242
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_254
timestamp 1701704242
transform 1 0 23920 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_266
timestamp 1701704242
transform 1 0 25024 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_278
timestamp 1701704242
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1701704242
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1701704242
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1701704242
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1701704242
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_329
timestamp 1701704242
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1701704242
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1701704242
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1701704242
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1701704242
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1701704242
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1701704242
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_97
timestamp 1701704242
transform 1 0 9476 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_244
timestamp 1701704242
transform 1 0 23000 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_262
timestamp 1701704242
transform 1 0 24656 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_274
timestamp 1701704242
transform 1 0 25760 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_286
timestamp 1701704242
transform 1 0 26864 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_298
timestamp 1701704242
transform 1 0 27968 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 1701704242
transform 1 0 28704 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1701704242
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_329
timestamp 1701704242
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1701704242
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1701704242
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1701704242
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1701704242
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1701704242
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1701704242
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_116
timestamp 1701704242
transform 1 0 11224 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_120
timestamp 1701704242
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_140
timestamp 1701704242
transform 1 0 13432 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_147
timestamp 1701704242
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_181
timestamp 1701704242
transform 1 0 17204 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1701704242
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1701704242
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1701704242
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1701704242
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1701704242
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1701704242
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1701704242
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1701704242
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_329
timestamp 1701704242
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1701704242
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1701704242
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1701704242
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1701704242
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1701704242
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1701704242
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1701704242
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1701704242
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_133
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_154
timestamp 1701704242
transform 1 0 14720 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1701704242
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_237
timestamp 1701704242
transform 1 0 22356 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1701704242
transform 1 0 23460 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1701704242
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1701704242
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1701704242
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1701704242
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1701704242
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 1701704242
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1701704242
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1701704242
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1701704242
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1701704242
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1701704242
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1701704242
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1701704242
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1701704242
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1701704242
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1701704242
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1701704242
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1701704242
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1701704242
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_149
timestamp 1701704242
transform 1 0 14260 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_155
timestamp 1701704242
transform 1 0 14812 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1701704242
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_169
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_191
timestamp 1701704242
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_199
timestamp 1701704242
transform 1 0 18860 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1701704242
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1701704242
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1701704242
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1701704242
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1701704242
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1701704242
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1701704242
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1701704242
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1701704242
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1701704242
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_329
timestamp 1701704242
transform 1 0 30820 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1701704242
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1701704242
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1701704242
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1701704242
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1701704242
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1701704242
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1701704242
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1701704242
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1701704242
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1701704242
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1701704242
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_153
timestamp 1701704242
transform 1 0 14628 0 1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_162
timestamp 1701704242
transform 1 0 15456 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_174
timestamp 1701704242
transform 1 0 16560 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_182
timestamp 1701704242
transform 1 0 17296 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_186
timestamp 1701704242
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_213
timestamp 1701704242
transform 1 0 20148 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_225
timestamp 1701704242
transform 1 0 21252 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_237
timestamp 1701704242
transform 1 0 22356 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_249
timestamp 1701704242
transform 1 0 23460 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1701704242
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1701704242
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1701704242
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1701704242
transform 1 0 27140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1701704242
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1701704242
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 1701704242
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_329
timestamp 1701704242
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1701704242
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1701704242
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1701704242
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1701704242
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1701704242
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1701704242
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1701704242
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1701704242
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1701704242
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1701704242
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1701704242
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1701704242
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1701704242
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1701704242
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1701704242
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1701704242
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1701704242
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1701704242
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1701704242
transform 1 0 20516 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1701704242
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1701704242
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1701704242
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1701704242
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1701704242
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1701704242
transform 1 0 25668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1701704242
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1701704242
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1701704242
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1701704242
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_329
timestamp 1701704242
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1701704242
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1701704242
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1701704242
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1701704242
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1701704242
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1701704242
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1701704242
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1701704242
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1701704242
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1701704242
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1701704242
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1701704242
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1701704242
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1701704242
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1701704242
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1701704242
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1701704242
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1701704242
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1701704242
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1701704242
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1701704242
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1701704242
transform 1 0 23092 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1701704242
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1701704242
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1701704242
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1701704242
transform 1 0 27140 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1701704242
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1701704242
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1701704242
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1701704242
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1701704242
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1701704242
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1701704242
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1701704242
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1701704242
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1701704242
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1701704242
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1701704242
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1701704242
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1701704242
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1701704242
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1701704242
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1701704242
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1701704242
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1701704242
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1701704242
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1701704242
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1701704242
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1701704242
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1701704242
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1701704242
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1701704242
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1701704242
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_329
timestamp 1701704242
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1701704242
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1701704242
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1701704242
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1701704242
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1701704242
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1701704242
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1701704242
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1701704242
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1701704242
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1701704242
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1701704242
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1701704242
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1701704242
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1701704242
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1701704242
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1701704242
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1701704242
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1701704242
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1701704242
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1701704242
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1701704242
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1701704242
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1701704242
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1701704242
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1701704242
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1701704242
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1701704242
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1701704242
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1701704242
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1701704242
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1701704242
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1701704242
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1701704242
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1701704242
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1701704242
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1701704242
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1701704242
transform 1 0 20516 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1701704242
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1701704242
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1701704242
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1701704242
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1701704242
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1701704242
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1701704242
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1701704242
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1701704242
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1701704242
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1701704242
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1701704242
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1701704242
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1701704242
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1701704242
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1701704242
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1701704242
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1701704242
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1701704242
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1701704242
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1701704242
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1701704242
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1701704242
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1701704242
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1701704242
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1701704242
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1701704242
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1701704242
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1701704242
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1701704242
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1701704242
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1701704242
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1701704242
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1701704242
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1701704242
transform 1 0 20516 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1701704242
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1701704242
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1701704242
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1701704242
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1701704242
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1701704242
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1701704242
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1701704242
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1701704242
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1701704242
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1701704242
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1701704242
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1701704242
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1701704242
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1701704242
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1701704242
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1701704242
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1701704242
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1701704242
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_137
timestamp 1701704242
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_145
timestamp 1701704242
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_157
timestamp 1701704242
transform 1 0 14996 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1701704242
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 1701704242
transform 1 0 19780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1701704242
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22356 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_249
timestamp 1701704242
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1701704242
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1701704242
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_305
timestamp 1701704242
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_329
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[1\].dly_stg05
timestamp 1701704242
transform -1 0 11408 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg06_18
timestamp 1701704242
transform -1 0 11224 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg06_19
timestamp 1701704242
transform -1 0 11960 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg06_20
timestamp 1701704242
transform -1 0 13800 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[1\].dly_stg07
timestamp 1701704242
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg08_17
timestamp 1701704242
transform -1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[2\].dly_stg05
timestamp 1701704242
transform 1 0 11224 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg06_22
timestamp 1701704242
transform -1 0 10856 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg06_23
timestamp 1701704242
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg06_24
timestamp 1701704242
transform -1 0 11592 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[2\].dly_stg07
timestamp 1701704242
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg08_21
timestamp 1701704242
transform 1 0 10764 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[3\].dly_stg05
timestamp 1701704242
transform 1 0 9476 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg06_26
timestamp 1701704242
transform -1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg06_27
timestamp 1701704242
transform -1 0 9476 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg06_28
timestamp 1701704242
transform 1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[3\].dly_stg07
timestamp 1701704242
transform 1 0 10028 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg08_25
timestamp 1701704242
transform 1 0 10488 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[4\].dly_stg05
timestamp 1701704242
transform 1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg06_30
timestamp 1701704242
transform -1 0 11776 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg06_31
timestamp 1701704242
transform 1 0 12788 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg06_32
timestamp 1701704242
transform -1 0 12512 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[4\].dly_stg07
timestamp 1701704242
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg08_29
timestamp 1701704242
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[5\].dly_stg05
timestamp 1701704242
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg06_34
timestamp 1701704242
transform -1 0 11224 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg06_35
timestamp 1701704242
transform -1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg06_36
timestamp 1701704242
transform -1 0 14536 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[5\].dly_stg07
timestamp 1701704242
transform 1 0 9476 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg08_33
timestamp 1701704242
transform 1 0 10028 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[6\].dly_stg05
timestamp 1701704242
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg06_38
timestamp 1701704242
transform -1 0 17848 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg06_39
timestamp 1701704242
transform 1 0 15456 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg06_40
timestamp 1701704242
transform 1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[6\].dly_stg07
timestamp 1701704242
transform 1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg08_37
timestamp 1701704242
transform -1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[7\].dly_stg05
timestamp 1701704242
transform 1 0 16468 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg06_42
timestamp 1701704242
transform -1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg06_43
timestamp 1701704242
transform 1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg06_44
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[7\].dly_stg07
timestamp 1701704242
transform -1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg08_41
timestamp 1701704242
transform 1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[8\].dly_stg05
timestamp 1701704242
transform 1 0 17940 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg06_46
timestamp 1701704242
transform 1 0 20148 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg06_47
timestamp 1701704242
transform -1 0 18492 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg06_48
timestamp 1701704242
transform -1 0 18216 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[8\].dly_stg07
timestamp 1701704242
transform 1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg08_45
timestamp 1701704242
transform 1 0 10304 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[9\].dly_stg05
timestamp 1701704242
transform 1 0 18492 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg06_50
timestamp 1701704242
transform 1 0 22632 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg06_51
timestamp 1701704242
transform 1 0 22264 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg06_52
timestamp 1701704242
transform -1 0 21804 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[9\].dly_stg07
timestamp 1701704242
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg08_49
timestamp 1701704242
transform 1 0 9936 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[10\].dly_stg05
timestamp 1701704242
transform -1 0 22264 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg06_54
timestamp 1701704242
transform 1 0 21712 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg06_55
timestamp 1701704242
transform 1 0 25300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg06_56
timestamp 1701704242
transform -1 0 23184 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[10\].dly_stg07
timestamp 1701704242
transform -1 0 10488 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg08_53
timestamp 1701704242
transform -1 0 10304 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[11\].dly_stg05
timestamp 1701704242
transform -1 0 22632 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg06_58
timestamp 1701704242
transform 1 0 24380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg06_59
timestamp 1701704242
transform 1 0 24932 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg06_60
timestamp 1701704242
transform -1 0 21528 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[11\].dly_stg07
timestamp 1701704242
transform 1 0 9476 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg08_57
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[12\].dly_stg05
timestamp 1701704242
transform -1 0 25576 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg06_62
timestamp 1701704242
transform 1 0 25576 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg06_63
timestamp 1701704242
transform -1 0 24380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg06_64
timestamp 1701704242
transform 1 0 25852 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[12\].dly_stg07
timestamp 1701704242
transform 1 0 9752 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg08_61
timestamp 1701704242
transform 1 0 10580 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[13\].dly_stg05
timestamp 1701704242
transform -1 0 19872 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg06_66
timestamp 1701704242
transform 1 0 19044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg06_67
timestamp 1701704242
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg06_68
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[13\].dly_stg07
timestamp 1701704242
transform -1 0 11132 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg08_65
timestamp 1701704242
transform 1 0 11684 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[14\].dly_stg05
timestamp 1701704242
transform 1 0 19320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg06_70
timestamp 1701704242
transform 1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg06_71
timestamp 1701704242
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg06_72
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  g_dly_chain\[14\].dly_stg07
timestamp 1701704242
transform 1 0 11132 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg08_69
timestamp 1701704242
transform 1 0 11960 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  g_dly_stp\[0\].dly_stp
timestamp 1701704242
transform 1 0 9568 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  g_dly_stp\[1\].dly_stp
timestamp 1701704242
transform -1 0 10672 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  g_dly_stp\[2\].dly_stp
timestamp 1701704242
transform 1 0 9844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  g_dly_strt\[0\].buf_chain
timestamp 1701704242
transform -1 0 13432 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  g_dly_strt\[1\].buf_chain
timestamp 1701704242
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  g_dly_strt\[2\].buf_chain
timestamp 1701704242
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1701704242
transform -1 0 13892 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 23202 0 23258 400 0 FreeSans 224 90 0 0 dbg_delay_stop
port 2 nsew signal tristate
flabel metal2 s 14830 19600 14886 20000 0 FreeSans 224 90 0 0 dbg_dly_sig[0]
port 3 nsew signal tristate
flabel metal2 s 22558 0 22614 400 0 FreeSans 224 90 0 0 dbg_dly_sig[10]
port 4 nsew signal tristate
flabel metal2 s 21270 0 21326 400 0 FreeSans 224 90 0 0 dbg_dly_sig[11]
port 5 nsew signal tristate
flabel metal3 s 31600 8168 32000 8288 0 FreeSans 480 0 0 0 dbg_dly_sig[12]
port 6 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 dbg_dly_sig[13]
port 7 nsew signal tristate
flabel metal3 s 31600 12248 32000 12368 0 FreeSans 480 0 0 0 dbg_dly_sig[14]
port 8 nsew signal tristate
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 dbg_dly_sig[15]
port 9 nsew signal tristate
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 dbg_dly_sig[1]
port 10 nsew signal tristate
flabel metal2 s 10322 0 10378 400 0 FreeSans 224 90 0 0 dbg_dly_sig[2]
port 11 nsew signal tristate
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 dbg_dly_sig[3]
port 12 nsew signal tristate
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 dbg_dly_sig[4]
port 13 nsew signal tristate
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 dbg_dly_sig[5]
port 14 nsew signal tristate
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 dbg_dly_sig[6]
port 15 nsew signal tristate
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 dbg_dly_sig[7]
port 16 nsew signal tristate
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 dbg_dly_sig[8]
port 17 nsew signal tristate
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 dbg_dly_sig[9]
port 18 nsew signal tristate
flabel metal2 s 15474 19600 15530 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[0]
port 19 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[1]
port 20 nsew signal tristate
flabel metal2 s 20626 19600 20682 20000 0 FreeSans 224 90 0 0 dbg_ring_ctr[2]
port 21 nsew signal tristate
flabel metal2 s 14186 19600 14242 20000 0 FreeSans 224 90 0 0 dbg_start_pulse
port 22 nsew signal tristate
flabel metal2 s 13542 19600 13598 20000 0 FreeSans 224 90 0 0 i_start
port 23 nsew signal input
flabel metal2 s 21914 0 21970 400 0 FreeSans 224 90 0 0 i_stop
port 24 nsew signal input
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 o_result_ctr[0]
port 25 nsew signal tristate
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 o_result_ctr[1]
port 26 nsew signal tristate
flabel metal3 s 31600 11568 32000 11688 0 FreeSans 480 0 0 0 o_result_ctr[2]
port 27 nsew signal tristate
flabel metal2 s 16762 19600 16818 20000 0 FreeSans 224 90 0 0 o_result_ring[0]
port 28 nsew signal tristate
flabel metal3 s 31600 6808 32000 6928 0 FreeSans 480 0 0 0 o_result_ring[10]
port 29 nsew signal tristate
flabel metal3 s 31600 7488 32000 7608 0 FreeSans 480 0 0 0 o_result_ring[11]
port 30 nsew signal tristate
flabel metal3 s 31600 8848 32000 8968 0 FreeSans 480 0 0 0 o_result_ring[12]
port 31 nsew signal tristate
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 o_result_ring[13]
port 32 nsew signal tristate
flabel metal3 s 31600 10888 32000 11008 0 FreeSans 480 0 0 0 o_result_ring[14]
port 33 nsew signal tristate
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 o_result_ring[15]
port 34 nsew signal tristate
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 o_result_ring[1]
port 35 nsew signal tristate
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 o_result_ring[2]
port 36 nsew signal tristate
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 o_result_ring[3]
port 37 nsew signal tristate
flabel metal2 s 12898 0 12954 400 0 FreeSans 224 90 0 0 o_result_ring[4]
port 38 nsew signal tristate
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 o_result_ring[5]
port 39 nsew signal tristate
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 o_result_ring[6]
port 40 nsew signal tristate
flabel metal2 s 20626 0 20682 400 0 FreeSans 224 90 0 0 o_result_ring[7]
port 41 nsew signal tristate
flabel metal2 s 19338 0 19394 400 0 FreeSans 224 90 0 0 o_result_ring[8]
port 42 nsew signal tristate
flabel metal2 s 19982 0 20038 400 0 FreeSans 224 90 0 0 o_result_ring[9]
port 43 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal2 15732 12852 15732 12852 0 _00_
rlabel metal1 16652 11798 16652 11798 0 _01_
rlabel metal1 20060 13430 20060 13430 0 _02_
rlabel metal1 14122 11186 14122 11186 0 _03_
rlabel metal1 13340 11866 13340 11866 0 _04_
rlabel metal1 15502 13362 15502 13362 0 _05_
rlabel metal1 17618 11730 17618 11730 0 _06_
rlabel metal1 21068 12070 21068 12070 0 _07_
rlabel metal1 20598 13906 20598 13906 0 _08_
rlabel metal1 20884 13838 20884 13838 0 _09_
rlabel metal1 20309 9078 20309 9078 0 clknet_0_i_stop
rlabel metal1 23000 8058 23000 8058 0 clknet_0_w_dly_sig1_n_ana_\[10\]
rlabel metal1 20976 7446 20976 7446 0 clknet_0_w_dly_sig1_n_ana_\[11\]
rlabel metal1 21206 9622 21206 9622 0 clknet_0_w_dly_sig1_n_ana_\[12\]
rlabel metal1 20654 11016 20654 11016 0 clknet_0_w_dly_sig1_n_ana_\[13\]
rlabel metal1 19320 9622 19320 9622 0 clknet_0_w_dly_sig1_n_ana_\[14\]
rlabel metal1 17250 11866 17250 11866 0 clknet_0_w_dly_sig1_n_ana_\[15\]
rlabel metal2 16330 10336 16330 10336 0 clknet_0_w_dly_sig1_n_ana_\[1\]
rlabel metal2 16192 6868 16192 6868 0 clknet_0_w_dly_sig1_n_ana_\[2\]
rlabel metal2 13662 8228 13662 8228 0 clknet_0_w_dly_sig1_n_ana_\[3\]
rlabel metal2 13662 7072 13662 7072 0 clknet_0_w_dly_sig1_n_ana_\[4\]
rlabel metal1 15732 5814 15732 5814 0 clknet_0_w_dly_sig1_n_ana_\[5\]
rlabel metal1 16560 7174 16560 7174 0 clknet_0_w_dly_sig1_n_ana_\[6\]
rlabel metal1 17158 5814 17158 5814 0 clknet_0_w_dly_sig1_n_ana_\[7\]
rlabel metal1 20424 8058 20424 8058 0 clknet_0_w_dly_sig1_n_ana_\[8\]
rlabel metal2 21206 6493 21206 6493 0 clknet_0_w_dly_sig1_n_ana_\[9\]
rlabel metal1 17250 8432 17250 8432 0 clknet_0_w_dly_stop
rlabel metal1 17894 12818 17894 12818 0 clknet_0_w_ring_ctr_clk
rlabel metal2 14582 11322 14582 11322 0 clknet_1_0__leaf_i_stop
rlabel metal2 21712 6596 21712 6596 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[10\]
rlabel metal1 24426 10642 24426 10642 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[11\]
rlabel metal2 24334 10404 24334 10404 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[12\]
rlabel metal1 17986 10234 17986 10234 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[13\]
rlabel metal2 18354 11492 18354 11492 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[14\]
rlabel metal1 14674 12784 14674 12784 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[15\]
rlabel metal1 11592 9554 11592 9554 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[1\]
rlabel metal1 11684 8602 11684 8602 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[2\]
rlabel metal1 10304 8602 10304 8602 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[3\]
rlabel metal1 12650 5746 12650 5746 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[4\]
rlabel metal2 14490 5338 14490 5338 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[5\]
rlabel metal1 15502 6256 15502 6256 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[6\]
rlabel metal1 19090 5814 19090 5814 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[7\]
rlabel metal2 20608 5644 20608 5644 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[8\]
rlabel metal1 21896 5746 21896 5746 0 clknet_1_0__leaf_w_dly_sig1_n_ana_\[9\]
rlabel metal1 16100 12274 16100 12274 0 clknet_1_0__leaf_w_ring_ctr_clk
rlabel metal1 18768 6834 18768 6834 0 clknet_1_1__leaf_i_stop
rlabel metal1 23276 6834 23276 6834 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[10\]
rlabel metal1 21482 5712 21482 5712 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[11\]
rlabel metal1 25806 9486 25806 9486 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[12\]
rlabel metal1 23736 10574 23736 10574 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[13\]
rlabel metal1 21942 10575 21942 10575 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[14\]
rlabel metal1 19550 13838 19550 13838 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[15\]
rlabel metal2 16882 9486 16882 9486 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[1\]
rlabel metal1 11546 7990 11546 7990 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[2\]
rlabel metal2 10534 7667 10534 7667 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[3\]
rlabel metal1 11776 6834 11776 6834 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[4\]
rlabel metal2 15226 9792 15226 9792 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[5\]
rlabel metal1 18952 8806 18952 8806 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[6\]
rlabel metal2 18722 8670 18722 8670 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[7\]
rlabel metal1 18584 10506 18584 10506 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[8\]
rlabel metal1 22724 6834 22724 6834 0 clknet_1_1__leaf_w_dly_sig1_n_ana_\[9\]
rlabel metal1 21160 13294 21160 13294 0 clknet_1_1__leaf_w_ring_ctr_clk
rlabel metal1 13294 5780 13294 5780 0 clknet_2_0__leaf_w_dly_stop
rlabel metal2 11454 11492 11454 11492 0 clknet_2_1__leaf_w_dly_stop
rlabel metal1 18584 6630 18584 6630 0 clknet_2_2__leaf_w_dly_stop
rlabel metal1 20746 5814 20746 5814 0 clknet_2_3__leaf_w_dly_stop
rlabel metal2 10258 6562 10258 6562 0 dbg_delay_stop
rlabel metal1 13018 10472 13018 10472 0 dbg_dly_sig[0]
rlabel metal1 21298 5576 21298 5576 0 dbg_dly_sig[10]
rlabel metal1 20378 6086 20378 6086 0 dbg_dly_sig[11]
rlabel metal1 23414 8568 23414 8568 0 dbg_dly_sig[12]
rlabel metal2 23046 8772 23046 8772 0 dbg_dly_sig[13]
rlabel metal3 30092 12308 30092 12308 0 dbg_dly_sig[14]
rlabel metal1 17020 8058 17020 8058 0 dbg_dly_sig[15]
rlabel metal2 14122 5235 14122 5235 0 dbg_dly_sig[1]
rlabel metal2 10442 7956 10442 7956 0 dbg_dly_sig[2]
rlabel metal2 13846 5338 13846 5338 0 dbg_dly_sig[3]
rlabel metal1 11914 7718 11914 7718 0 dbg_dly_sig[4]
rlabel metal2 12282 415 12282 415 0 dbg_dly_sig[5]
rlabel metal1 13984 5542 13984 5542 0 dbg_dly_sig[6]
rlabel metal1 16652 5542 16652 5542 0 dbg_dly_sig[7]
rlabel metal1 17664 6358 17664 6358 0 dbg_dly_sig[8]
rlabel metal1 18446 6086 18446 6086 0 dbg_dly_sig[9]
rlabel metal1 14950 10642 14950 10642 0 dbg_ring_ctr[0]
rlabel metal1 19320 13838 19320 13838 0 dbg_ring_ctr[1]
rlabel metal2 20654 17486 20654 17486 0 dbg_ring_ctr[2]
rlabel metal1 13800 11662 13800 11662 0 dbg_start_pulse
rlabel metal1 13708 18802 13708 18802 0 i_start
rlabel metal2 18906 9010 18906 9010 0 i_stop
rlabel metal1 13616 12274 13616 12274 0 net1
rlabel metal1 10994 9622 10994 9622 0 net10
rlabel metal2 21574 6494 21574 6494 0 net11
rlabel metal2 19642 5967 19642 5967 0 net12
rlabel metal1 24564 11050 24564 11050 0 net13
rlabel metal1 20838 5780 20838 5780 0 net14
rlabel metal1 22034 6257 22034 6257 0 net15
rlabel metal1 20286 10030 20286 10030 0 net16
rlabel metal1 20102 5882 20102 5882 0 net17
rlabel metal1 10810 10132 10810 10132 0 net18
rlabel metal1 11270 9044 11270 9044 0 net19
rlabel metal1 19642 4658 19642 4658 0 net2
rlabel metal1 11684 9486 11684 9486 0 net20
rlabel metal1 13708 8602 13708 8602 0 net21
rlabel metal1 10258 10064 10258 10064 0 net22
rlabel metal1 10672 7922 10672 7922 0 net23
rlabel metal1 13156 7310 13156 7310 0 net24
rlabel metal1 14756 5134 14756 5134 0 net25
rlabel metal1 9982 10132 9982 10132 0 net26
rlabel metal1 10120 8058 10120 8058 0 net27
rlabel metal2 12006 8092 12006 8092 0 net28
rlabel via2 10442 10115 10442 10115 0 net29
rlabel metal1 18170 5168 18170 5168 0 net3
rlabel metal2 9706 10574 9706 10574 0 net30
rlabel metal1 11270 6800 11270 6800 0 net31
rlabel metal2 12926 6834 12926 6834 0 net32
rlabel metal2 12374 6018 12374 6018 0 net33
rlabel metal1 9430 10064 9430 10064 0 net34
rlabel metal1 10350 7956 10350 7956 0 net35
rlabel metal1 14030 5338 14030 5338 0 net36
rlabel viali 14393 4658 14393 4658 0 net37
rlabel metal1 8970 10132 8970 10132 0 net38
rlabel metal2 17710 5803 17710 5803 0 net39
rlabel metal1 18860 7718 18860 7718 0 net4
rlabel metal1 16629 5746 16629 5746 0 net40
rlabel metal1 16141 6154 16141 6154 0 net41
rlabel metal1 9890 10540 9890 10540 0 net42
rlabel metal1 17986 5100 17986 5100 0 net43
rlabel metal1 17526 6256 17526 6256 0 net44
rlabel metal2 18814 6663 18814 6663 0 net45
rlabel via1 9602 10574 9602 10574 0 net46
rlabel metal1 19412 4726 19412 4726 0 net47
rlabel metal2 18354 5780 18354 5780 0 net48
rlabel metal1 18160 6834 18160 6834 0 net49
rlabel metal1 10534 7888 10534 7888 0 net5
rlabel metal1 10166 10574 10166 10574 0 net50
rlabel metal2 22218 6426 22218 6426 0 net51
rlabel metal1 19596 6222 19596 6222 0 net52
rlabel metal1 20419 6834 20419 6834 0 net53
rlabel metal1 9706 11220 9706 11220 0 net54
rlabel metal2 21850 6596 21850 6596 0 net55
rlabel metal2 19826 6273 19826 6273 0 net56
rlabel metal2 23046 7106 23046 7106 0 net57
rlabel metal2 9982 11628 9982 11628 0 net58
rlabel metal2 25438 9724 25438 9724 0 net59
rlabel metal1 11454 5780 11454 5780 0 net6
rlabel metal1 23598 8364 23598 8364 0 net60
rlabel metal2 24150 6970 24150 6970 0 net61
rlabel metal1 10810 11662 10810 11662 0 net62
rlabel via2 19826 5763 19826 5763 0 net63
rlabel metal1 23276 8398 23276 8398 0 net64
rlabel metal1 25499 9418 25499 9418 0 net65
rlabel metal1 11362 11696 11362 11696 0 net66
rlabel metal1 19274 5746 19274 5746 0 net67
rlabel metal1 20332 7310 20332 7310 0 net68
rlabel metal1 21454 10506 21454 10506 0 net69
rlabel metal1 10350 9010 10350 9010 0 net7
rlabel metal2 11638 11900 11638 11900 0 net70
rlabel metal1 22977 14314 22977 14314 0 net71
rlabel metal2 17158 9724 17158 9724 0 net72
rlabel metal1 17250 9044 17250 9044 0 net73
rlabel metal1 12650 11696 12650 11696 0 net74
rlabel metal2 13570 11492 13570 11492 0 net75
rlabel metal1 13478 12682 13478 12682 0 net76
rlabel metal1 13984 10778 13984 10778 0 net77
rlabel metal1 21022 12342 21022 12342 0 net78
rlabel metal1 18584 11662 18584 11662 0 net79
rlabel metal1 10212 8398 10212 8398 0 net8
rlabel metal2 15318 13464 15318 13464 0 net80
rlabel metal1 13662 11594 13662 11594 0 net81
rlabel metal1 11546 9010 11546 9010 0 net9
rlabel metal1 18308 11254 18308 11254 0 o_result_ctr[0]
rlabel metal2 20010 17520 20010 17520 0 o_result_ctr[1]
rlabel metal2 28290 11475 28290 11475 0 o_result_ctr[2]
rlabel metal1 16652 10234 16652 10234 0 o_result_ring[0]
rlabel metal1 22310 6868 22310 6868 0 o_result_ring[10]
rlabel metal2 22034 6681 22034 6681 0 o_result_ring[11]
rlabel metal1 22816 8602 22816 8602 0 o_result_ring[12]
rlabel metal2 23230 9843 23230 9843 0 o_result_ring[13]
rlabel metal1 22816 9350 22816 9350 0 o_result_ring[14]
rlabel metal1 20792 9962 20792 9962 0 o_result_ring[15]
rlabel metal2 14628 8908 14628 8908 0 o_result_ring[1]
rlabel metal2 17572 6900 17572 6900 0 o_result_ring[2]
rlabel metal1 16560 7718 16560 7718 0 o_result_ring[3]
rlabel metal2 12880 3468 12880 3468 0 o_result_ring[4]
rlabel metal2 13570 3492 13570 3492 0 o_result_ring[5]
rlabel metal1 16008 5542 16008 5542 0 o_result_ring[6]
rlabel metal1 19780 7174 19780 7174 0 o_result_ring[7]
rlabel metal2 19366 1588 19366 1588 0 o_result_ring[8]
rlabel metal2 20148 5644 20148 5644 0 o_result_ring[9]
rlabel metal1 18722 11254 18722 11254 0 r_dly_store_ctr\[0\]
rlabel metal1 21758 12342 21758 12342 0 r_dly_store_ctr\[1\]
rlabel metal1 23322 10778 23322 10778 0 r_dly_store_ctr\[2\]
rlabel metal2 16238 10319 16238 10319 0 r_dly_store_ring\[0\]
rlabel metal1 21252 6698 21252 6698 0 r_dly_store_ring\[10\]
rlabel metal2 22218 7038 22218 7038 0 r_dly_store_ring\[11\]
rlabel metal1 23138 8330 23138 8330 0 r_dly_store_ring\[12\]
rlabel metal1 23414 9418 23414 9418 0 r_dly_store_ring\[13\]
rlabel metal2 21942 10302 21942 10302 0 r_dly_store_ring\[14\]
rlabel metal1 19366 9350 19366 9350 0 r_dly_store_ring\[15\]
rlabel metal1 13892 8602 13892 8602 0 r_dly_store_ring\[1\]
rlabel metal1 16514 9112 16514 9112 0 r_dly_store_ring\[2\]
rlabel metal1 16284 7922 16284 7922 0 r_dly_store_ring\[3\]
rlabel metal1 12236 9078 12236 9078 0 r_dly_store_ring\[4\]
rlabel metal2 12466 6596 12466 6596 0 r_dly_store_ring\[5\]
rlabel metal1 15916 5746 15916 5746 0 r_dly_store_ring\[6\]
rlabel metal1 17710 6426 17710 6426 0 r_dly_store_ring\[7\]
rlabel metal1 19044 8602 19044 8602 0 r_dly_store_ring\[8\]
rlabel metal1 19504 6698 19504 6698 0 r_dly_store_ring\[9\]
rlabel metal1 14628 12070 14628 12070 0 r_ring_ctr\[0\]
rlabel metal1 19090 11628 19090 11628 0 r_ring_ctr\[1\]
rlabel metal1 19182 13158 19182 13158 0 r_ring_ctr\[2\]
rlabel metal2 12926 11526 12926 11526 0 w_dly_sig1_ana_\[1\]
rlabel metal1 13018 12240 13018 12240 0 w_dly_sig1_n_ana_\[0\]
rlabel metal2 22126 7174 22126 7174 0 w_dly_sig1_n_ana_\[10\]
rlabel metal2 22402 7106 22402 7106 0 w_dly_sig1_n_ana_\[11\]
rlabel metal1 23598 9452 23598 9452 0 w_dly_sig1_n_ana_\[12\]
rlabel metal1 19550 5882 19550 5882 0 w_dly_sig1_n_ana_\[13\]
rlabel metal1 19734 5678 19734 5678 0 w_dly_sig1_n_ana_\[14\]
rlabel metal1 18170 11662 18170 11662 0 w_dly_sig1_n_ana_\[15\]
rlabel metal2 15318 8466 15318 8466 0 w_dly_sig1_n_ana_\[1\]
rlabel metal1 13317 9078 13317 9078 0 w_dly_sig1_n_ana_\[2\]
rlabel metal2 9706 8177 9706 8177 0 w_dly_sig1_n_ana_\[3\]
rlabel metal2 12374 7650 12374 7650 0 w_dly_sig1_n_ana_\[4\]
rlabel metal1 14214 6766 14214 6766 0 w_dly_sig1_n_ana_\[5\]
rlabel metal1 16422 7344 16422 7344 0 w_dly_sig1_n_ana_\[6\]
rlabel metal2 17204 6900 17204 6900 0 w_dly_sig1_n_ana_\[7\]
rlabel metal1 18630 7922 18630 7922 0 w_dly_sig1_n_ana_\[8\]
rlabel metal1 19642 6154 19642 6154 0 w_dly_sig1_n_ana_\[9\]
rlabel metal2 11546 11458 11546 11458 0 w_dly_sig2_ana_\[1\]
rlabel metal1 12696 11866 12696 11866 0 w_dly_sig2_n_ana_\[0\]
rlabel metal1 10350 10778 10350 10778 0 w_dly_sig2_n_ana_\[10\]
rlabel metal2 9614 11798 9614 11798 0 w_dly_sig2_n_ana_\[11\]
rlabel metal2 9890 11458 9890 11458 0 w_dly_sig2_n_ana_\[12\]
rlabel metal2 11086 12070 11086 12070 0 w_dly_sig2_n_ana_\[13\]
rlabel metal1 11224 11866 11224 11866 0 w_dly_sig2_n_ana_\[14\]
rlabel metal1 12006 11628 12006 11628 0 w_dly_sig2_n_ana_\[15\]
rlabel metal1 11270 10540 11270 10540 0 w_dly_sig2_n_ana_\[1\]
rlabel metal1 10764 10234 10764 10234 0 w_dly_sig2_n_ana_\[2\]
rlabel metal1 10350 10234 10350 10234 0 w_dly_sig2_n_ana_\[3\]
rlabel metal2 9890 10642 9890 10642 0 w_dly_sig2_n_ana_\[4\]
rlabel metal1 9844 10234 9844 10234 0 w_dly_sig2_n_ana_\[5\]
rlabel metal2 9338 10404 9338 10404 0 w_dly_sig2_n_ana_\[6\]
rlabel metal1 9706 9962 9706 9962 0 w_dly_sig2_n_ana_\[7\]
rlabel metal1 9752 10778 9752 10778 0 w_dly_sig2_n_ana_\[8\]
rlabel metal1 9982 10608 9982 10608 0 w_dly_sig2_n_ana_\[9\]
rlabel metal1 13754 9690 13754 9690 0 w_dly_stop
rlabel metal2 10626 9316 10626 9316 0 w_dly_stop_ana_\[1\]
rlabel metal1 9890 9520 9890 9520 0 w_dly_stop_ana_\[2\]
rlabel metal2 13202 12206 13202 12206 0 w_dly_strt_ana_\[1\]
rlabel metal2 12466 12070 12466 12070 0 w_dly_strt_ana_\[2\]
rlabel metal1 13662 12104 13662 12104 0 w_dly_strt_ana_\[3\]
rlabel metal1 17089 12342 17089 12342 0 w_ring_ctr_clk
rlabel metal1 14628 11322 14628 11322 0 w_strt_pulse_n
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
