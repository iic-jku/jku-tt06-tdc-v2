magic
tech sky130A
magscale 1 2
timestamp 1711752330
<< viali >>
rect 857 21641 891 21675
rect 1593 21641 1627 21675
rect 2329 21641 2363 21675
rect 3249 21641 3283 21675
rect 3801 21641 3835 21675
rect 4537 21641 4571 21675
rect 5273 21641 5307 21675
rect 6009 21641 6043 21675
rect 6745 21641 6779 21675
rect 7481 21641 7515 21675
rect 8217 21641 8251 21675
rect 8769 21641 8803 21675
rect 9689 21641 9723 21675
rect 10425 21641 10459 21675
rect 11161 21641 11195 21675
rect 27721 21641 27755 21675
rect 12909 21573 12943 21607
rect 16221 21573 16255 21607
rect 23305 21573 23339 21607
rect 29009 21573 29043 21607
rect 14381 21505 14415 21539
rect 14565 21505 14599 21539
rect 21741 21505 21775 21539
rect 29285 21505 29319 21539
rect 9137 21437 9171 21471
rect 9229 21437 9263 21471
rect 9413 21437 9447 21471
rect 11529 21437 11563 21471
rect 14657 21437 14691 21471
rect 15853 21437 15887 21471
rect 16405 21437 16439 21471
rect 20085 21437 20119 21471
rect 21465 21437 21499 21471
rect 23489 21437 23523 21471
rect 24041 21437 24075 21471
rect 24593 21437 24627 21471
rect 24685 21437 24719 21471
rect 25237 21437 25271 21471
rect 25789 21437 25823 21471
rect 25881 21437 25915 21471
rect 26801 21437 26835 21471
rect 28549 21437 28583 21471
rect 29193 21437 29227 21471
rect 29561 21437 29595 21471
rect 30021 21437 30055 21471
rect 11774 21369 11808 21403
rect 13829 21369 13863 21403
rect 19818 21369 19852 21403
rect 22008 21369 22042 21403
rect 23857 21369 23891 21403
rect 24869 21369 24903 21403
rect 27813 21369 27847 21403
rect 27997 21369 28031 21403
rect 28181 21369 28215 21403
rect 8953 21301 8987 21335
rect 14105 21301 14139 21335
rect 15025 21301 15059 21335
rect 15761 21301 15795 21335
rect 18705 21301 18739 21335
rect 23121 21301 23155 21335
rect 24593 21301 24627 21335
rect 26065 21301 26099 21335
rect 26709 21301 26743 21335
rect 28457 21301 28491 21335
rect 29745 21301 29779 21335
rect 29837 21301 29871 21335
rect 10149 21097 10183 21131
rect 11437 21097 11471 21131
rect 12541 21097 12575 21131
rect 13369 21097 13403 21131
rect 16129 21097 16163 21131
rect 16681 21097 16715 21131
rect 19073 21097 19107 21131
rect 21005 21097 21039 21131
rect 21833 21097 21867 21131
rect 22201 21097 22235 21131
rect 29469 21097 29503 21131
rect 13185 21029 13219 21063
rect 14832 21029 14866 21063
rect 23274 21029 23308 21063
rect 26709 21029 26743 21063
rect 27629 21029 27663 21063
rect 29561 21029 29595 21063
rect 9025 20961 9059 20995
rect 10425 20961 10459 20995
rect 10977 20961 11011 20995
rect 11161 20961 11195 20995
rect 11253 20961 11287 20995
rect 11897 20961 11931 20995
rect 12449 20961 12483 20995
rect 13921 20961 13955 20995
rect 14289 20961 14323 20995
rect 14381 20961 14415 20995
rect 16313 20961 16347 20995
rect 17794 20961 17828 20995
rect 18429 20961 18463 20995
rect 18613 20961 18647 20995
rect 18889 20961 18923 20995
rect 20545 20961 20579 20995
rect 20913 20961 20947 20995
rect 21097 20961 21131 20995
rect 21281 20961 21315 20995
rect 21649 20961 21683 20995
rect 21925 20961 21959 20995
rect 22109 20961 22143 20995
rect 22385 20961 22419 20995
rect 23029 20961 23063 20995
rect 24685 20961 24719 20995
rect 24777 20961 24811 20995
rect 25145 20961 25179 20995
rect 25329 20961 25363 20995
rect 25513 20961 25547 20995
rect 25697 20961 25731 20995
rect 25789 20961 25823 20995
rect 26249 20961 26283 20995
rect 26433 20961 26467 20995
rect 27077 20961 27111 20995
rect 27169 20961 27203 20995
rect 27261 20961 27295 20995
rect 27537 20961 27571 20995
rect 27721 20961 27755 20995
rect 29029 20961 29063 20995
rect 29929 20961 29963 20995
rect 8769 20893 8803 20927
rect 12725 20893 12759 20927
rect 14013 20893 14047 20927
rect 14565 20893 14599 20927
rect 18061 20893 18095 20927
rect 20453 20893 20487 20927
rect 20821 20893 20855 20927
rect 21557 20893 21591 20927
rect 22017 20893 22051 20927
rect 24961 20893 24995 20927
rect 25605 20893 25639 20927
rect 26801 20893 26835 20927
rect 27445 20893 27479 20927
rect 29285 20893 29319 20927
rect 18429 20825 18463 20859
rect 20637 20825 20671 20859
rect 21281 20825 21315 20859
rect 21373 20825 21407 20859
rect 24685 20825 24719 20859
rect 25145 20825 25179 20859
rect 26433 20825 26467 20859
rect 26525 20825 26559 20859
rect 26985 20825 27019 20859
rect 27077 20825 27111 20859
rect 27169 20825 27203 20859
rect 29745 20825 29779 20859
rect 10241 20757 10275 20791
rect 10977 20757 11011 20791
rect 12817 20757 12851 20791
rect 12909 20757 12943 20791
rect 15945 20757 15979 20791
rect 18153 20757 18187 20791
rect 20729 20757 20763 20791
rect 24409 20757 24443 20791
rect 25973 20757 26007 20791
rect 26065 20757 26099 20791
rect 27905 20757 27939 20791
rect 8861 20553 8895 20587
rect 12817 20553 12851 20587
rect 15669 20553 15703 20587
rect 18889 20553 18923 20587
rect 20913 20553 20947 20587
rect 24961 20553 24995 20587
rect 25053 20553 25087 20587
rect 27445 20553 27479 20587
rect 11345 20485 11379 20519
rect 13553 20485 13587 20519
rect 17049 20485 17083 20519
rect 21741 20485 21775 20519
rect 22477 20485 22511 20519
rect 24501 20485 24535 20519
rect 28457 20485 28491 20519
rect 29009 20485 29043 20519
rect 9965 20417 9999 20451
rect 13185 20417 13219 20451
rect 14105 20417 14139 20451
rect 14565 20417 14599 20451
rect 16405 20417 16439 20451
rect 17141 20417 17175 20451
rect 24777 20417 24811 20451
rect 25421 20417 25455 20451
rect 26801 20417 26835 20451
rect 27721 20417 27755 20451
rect 28181 20417 28215 20451
rect 4905 20349 4939 20383
rect 6009 20349 6043 20383
rect 6745 20349 6779 20383
rect 8677 20349 8711 20383
rect 9229 20349 9263 20383
rect 9597 20349 9631 20383
rect 9689 20349 9723 20383
rect 9873 20349 9907 20383
rect 10232 20349 10266 20383
rect 11437 20349 11471 20383
rect 11713 20349 11747 20383
rect 13001 20349 13035 20383
rect 13737 20349 13771 20383
rect 13829 20349 13863 20383
rect 14749 20349 14783 20383
rect 15117 20349 15151 20383
rect 15301 20349 15335 20383
rect 16681 20349 16715 20383
rect 17601 20349 17635 20383
rect 17785 20349 17819 20383
rect 18092 20349 18126 20383
rect 18337 20349 18371 20383
rect 19068 20349 19102 20383
rect 19385 20349 19419 20383
rect 19533 20349 19567 20383
rect 20269 20349 20303 20383
rect 20361 20349 20395 20383
rect 20539 20349 20573 20383
rect 20729 20349 20763 20383
rect 20913 20349 20947 20383
rect 21925 20349 21959 20383
rect 22201 20349 22235 20383
rect 22385 20349 22419 20383
rect 22615 20349 22649 20383
rect 22753 20349 22787 20383
rect 22973 20349 23007 20383
rect 23121 20349 23155 20383
rect 24685 20349 24719 20383
rect 25237 20349 25271 20383
rect 26424 20349 26458 20383
rect 26709 20349 26743 20383
rect 26893 20349 26927 20383
rect 26985 20349 27019 20383
rect 27629 20349 27663 20383
rect 27813 20349 27847 20383
rect 28089 20349 28123 20383
rect 28457 20349 28491 20383
rect 28549 20349 28583 20383
rect 30389 20349 30423 20383
rect 6990 20281 7024 20315
rect 15761 20281 15795 20315
rect 19165 20281 19199 20315
rect 19257 20281 19291 20315
rect 22845 20281 22879 20315
rect 24961 20281 24995 20315
rect 28365 20281 28399 20315
rect 28733 20281 28767 20315
rect 30122 20281 30156 20315
rect 5089 20213 5123 20247
rect 6193 20213 6227 20247
rect 8125 20213 8159 20247
rect 9045 20213 9079 20247
rect 9781 20213 9815 20247
rect 11621 20213 11655 20247
rect 16589 20213 16623 20247
rect 20085 20213 20119 20247
rect 20453 20213 20487 20247
rect 26249 20213 26283 20247
rect 27169 20213 27203 20247
rect 28089 20213 28123 20247
rect 3433 20009 3467 20043
rect 6469 20009 6503 20043
rect 7941 20009 7975 20043
rect 9873 20009 9907 20043
rect 11253 20009 11287 20043
rect 13829 20009 13863 20043
rect 14289 20009 14323 20043
rect 16221 20009 16255 20043
rect 16865 20009 16899 20043
rect 19073 20009 19107 20043
rect 22661 20009 22695 20043
rect 24961 20009 24995 20043
rect 28733 20009 28767 20043
rect 29929 20009 29963 20043
rect 6806 19941 6840 19975
rect 9597 19941 9631 19975
rect 10241 19941 10275 19975
rect 11590 19941 11624 19975
rect 13553 19941 13587 19975
rect 16957 19941 16991 19975
rect 17960 19941 17994 19975
rect 20361 19941 20395 19975
rect 24501 19941 24535 19975
rect 24593 19941 24627 19975
rect 25145 19941 25179 19975
rect 27822 19941 27856 19975
rect 28457 19941 28491 19975
rect 29193 19941 29227 19975
rect 2973 19873 3007 19907
rect 3249 19873 3283 19907
rect 3709 19873 3743 19907
rect 4813 19873 4847 19907
rect 4997 19873 5031 19907
rect 5089 19873 5123 19907
rect 5365 19873 5399 19907
rect 6285 19873 6319 19907
rect 6561 19873 6595 19907
rect 8861 19873 8895 19907
rect 8953 19873 8987 19907
rect 9045 19873 9079 19907
rect 9873 19873 9907 19907
rect 10057 19873 10091 19907
rect 11069 19873 11103 19907
rect 13185 19873 13219 19907
rect 13278 19873 13312 19907
rect 13461 19873 13495 19907
rect 13691 19873 13725 19907
rect 13909 19873 13943 19907
rect 14832 19873 14866 19907
rect 16497 19873 16531 19907
rect 16681 19873 16715 19907
rect 17233 19873 17267 19907
rect 17325 19873 17359 19907
rect 17417 19873 17451 19907
rect 19349 19873 19383 19907
rect 20085 19873 20119 19907
rect 20453 19873 20487 19907
rect 21537 19873 21571 19907
rect 23009 19873 23043 19907
rect 24409 19873 24443 19907
rect 24777 19873 24811 19907
rect 24869 19873 24903 19907
rect 25973 19873 26007 19907
rect 26157 19873 26191 19907
rect 28365 19873 28399 19907
rect 28549 19873 28583 19907
rect 28641 19873 28675 19907
rect 28825 19873 28859 19907
rect 29745 19873 29779 19907
rect 5641 19805 5675 19839
rect 8677 19805 8711 19839
rect 9321 19805 9355 19839
rect 11345 19805 11379 19839
rect 14013 19805 14047 19839
rect 14565 19805 14599 19839
rect 17601 19805 17635 19839
rect 17693 19805 17727 19839
rect 20729 19805 20763 19839
rect 21281 19805 21315 19839
rect 22753 19805 22787 19839
rect 28089 19805 28123 19839
rect 29469 19805 29503 19839
rect 3893 19737 3927 19771
rect 5365 19737 5399 19771
rect 5457 19737 5491 19771
rect 9045 19737 9079 19771
rect 9137 19737 9171 19771
rect 9781 19737 9815 19771
rect 17141 19737 17175 19771
rect 17233 19737 17267 19771
rect 19165 19737 19199 19771
rect 20177 19737 20211 19771
rect 20453 19737 20487 19771
rect 20545 19737 20579 19771
rect 3157 19669 3191 19703
rect 4537 19669 4571 19703
rect 4997 19669 5031 19703
rect 5273 19669 5307 19703
rect 6101 19669 6135 19703
rect 8585 19669 8619 19703
rect 8953 19669 8987 19703
rect 12725 19669 12759 19703
rect 13921 19669 13955 19703
rect 15945 19669 15979 19703
rect 17509 19669 17543 19703
rect 19993 19669 20027 19703
rect 20269 19669 20303 19703
rect 24133 19669 24167 19703
rect 24225 19669 24259 19703
rect 26709 19669 26743 19703
rect 29285 19669 29319 19703
rect 3249 19465 3283 19499
rect 3525 19465 3559 19499
rect 3985 19465 4019 19499
rect 7389 19465 7423 19499
rect 8953 19465 8987 19499
rect 9229 19465 9263 19499
rect 9965 19465 9999 19499
rect 11253 19465 11287 19499
rect 13921 19465 13955 19499
rect 17601 19465 17635 19499
rect 17877 19465 17911 19499
rect 20913 19465 20947 19499
rect 22109 19465 22143 19499
rect 23673 19465 23707 19499
rect 24685 19465 24719 19499
rect 30021 19465 30055 19499
rect 4077 19397 4111 19431
rect 10609 19397 10643 19431
rect 11161 19397 11195 19431
rect 18061 19397 18095 19431
rect 18153 19397 18187 19431
rect 19717 19397 19751 19431
rect 20361 19397 20395 19431
rect 29193 19397 29227 19431
rect 29653 19397 29687 19431
rect 10057 19329 10091 19363
rect 10701 19329 10735 19363
rect 13553 19329 13587 19363
rect 15853 19329 15887 19363
rect 16037 19329 16071 19363
rect 17785 19329 17819 19363
rect 19625 19329 19659 19363
rect 24869 19329 24903 19363
rect 29561 19329 29595 19363
rect 3433 19261 3467 19295
rect 3709 19261 3743 19295
rect 3801 19261 3835 19295
rect 3985 19261 4019 19295
rect 4629 19261 4663 19295
rect 4905 19261 4939 19295
rect 5172 19261 5206 19295
rect 6377 19261 6411 19295
rect 6561 19261 6595 19295
rect 6653 19261 6687 19295
rect 6929 19261 6963 19295
rect 7205 19261 7239 19295
rect 7389 19261 7423 19295
rect 8677 19261 8711 19295
rect 8769 19261 8803 19295
rect 8861 19261 8895 19295
rect 8953 19261 8987 19295
rect 9137 19261 9171 19295
rect 9229 19261 9263 19295
rect 9413 19261 9447 19295
rect 9597 19261 9631 19295
rect 9689 19261 9723 19295
rect 9781 19261 9815 19295
rect 9873 19261 9907 19295
rect 10149 19261 10183 19295
rect 10333 19257 10367 19291
rect 10609 19261 10643 19295
rect 11253 19261 11287 19295
rect 11437 19261 11471 19295
rect 13737 19255 13771 19289
rect 14289 19261 14323 19295
rect 17417 19261 17451 19295
rect 17601 19261 17635 19295
rect 17693 19261 17727 19295
rect 18061 19261 18095 19295
rect 18705 19261 18739 19295
rect 19165 19261 19199 19295
rect 19349 19261 19383 19295
rect 19717 19261 19751 19295
rect 19809 19261 19843 19295
rect 19901 19261 19935 19295
rect 20177 19261 20211 19295
rect 20361 19261 20395 19295
rect 20459 19261 20493 19295
rect 20637 19261 20671 19295
rect 20729 19261 20763 19295
rect 21925 19261 21959 19295
rect 22293 19261 22327 19295
rect 24133 19261 24167 19295
rect 24501 19261 24535 19295
rect 24961 19261 24995 19295
rect 25053 19261 25087 19295
rect 26801 19261 26835 19295
rect 26893 19261 26927 19295
rect 26985 19261 27019 19295
rect 27261 19261 27295 19295
rect 29285 19271 29319 19305
rect 29653 19261 29687 19295
rect 29745 19261 29779 19295
rect 30297 19261 30331 19295
rect 10885 19193 10919 19227
rect 10977 19193 11011 19227
rect 11682 19193 11716 19227
rect 14534 19193 14568 19227
rect 17969 19193 18003 19227
rect 18337 19193 18371 19227
rect 19257 19193 19291 19227
rect 19441 19193 19475 19227
rect 20085 19193 20119 19227
rect 22560 19193 22594 19227
rect 24317 19193 24351 19227
rect 24409 19193 24443 19227
rect 29009 19193 29043 19227
rect 29377 19193 29411 19227
rect 4445 19125 4479 19159
rect 6285 19125 6319 19159
rect 6469 19125 6503 19159
rect 6837 19125 6871 19159
rect 7113 19125 7147 19159
rect 10517 19125 10551 19159
rect 12817 19125 12851 19159
rect 15669 19125 15703 19159
rect 16129 19125 16163 19159
rect 16497 19125 16531 19159
rect 19809 19125 19843 19159
rect 20545 19125 20579 19159
rect 25237 19125 25271 19159
rect 27169 19125 27203 19159
rect 27445 19125 27479 19159
rect 29285 19125 29319 19159
rect 29929 19125 29963 19159
rect 30481 19125 30515 19159
rect 5365 18921 5399 18955
rect 6101 18921 6135 18955
rect 9321 18921 9355 18955
rect 10149 18921 10183 18955
rect 10701 18921 10735 18955
rect 11253 18921 11287 18955
rect 14657 18921 14691 18955
rect 18245 18921 18279 18955
rect 18521 18921 18555 18955
rect 19257 18921 19291 18955
rect 23029 18921 23063 18955
rect 24041 18921 24075 18955
rect 24317 18921 24351 18955
rect 25504 18921 25538 18955
rect 27077 18921 27111 18955
rect 27629 18921 27663 18955
rect 29101 18921 29135 18955
rect 4997 18853 5031 18887
rect 5641 18853 5675 18887
rect 6929 18853 6963 18887
rect 7358 18853 7392 18887
rect 13001 18853 13035 18887
rect 13737 18853 13771 18887
rect 16374 18853 16408 18887
rect 20637 18853 20671 18887
rect 21526 18853 21560 18887
rect 24409 18853 24443 18887
rect 26525 18853 26559 18887
rect 28825 18853 28859 18887
rect 30858 18853 30892 18887
rect 2881 18785 2915 18819
rect 3801 18785 3835 18819
rect 3985 18785 4019 18819
rect 4077 18785 4111 18819
rect 4537 18785 4571 18819
rect 5273 18785 5307 18819
rect 5365 18785 5399 18819
rect 6009 18785 6043 18819
rect 6193 18785 6227 18819
rect 6561 18785 6595 18819
rect 6653 18785 6687 18819
rect 8769 18785 8803 18819
rect 9321 18785 9355 18819
rect 9689 18785 9723 18819
rect 9965 18807 9999 18841
rect 10081 18785 10115 18819
rect 10235 18785 10269 18819
rect 10333 18785 10367 18819
rect 10609 18785 10643 18819
rect 10793 18785 10827 18819
rect 11069 18785 11103 18819
rect 12725 18785 12759 18819
rect 12818 18785 12852 18819
rect 13093 18785 13127 18819
rect 13190 18785 13224 18819
rect 13461 18785 13495 18819
rect 13554 18785 13588 18819
rect 13829 18785 13863 18819
rect 13967 18785 14001 18819
rect 14197 18785 14231 18819
rect 14473 18785 14507 18819
rect 17785 18785 17819 18819
rect 18153 18785 18187 18819
rect 18337 18785 18371 18819
rect 18429 18785 18463 18819
rect 18613 18785 18647 18819
rect 19073 18785 19107 18819
rect 19625 18785 19659 18819
rect 19809 18785 19843 18819
rect 19993 18785 20027 18819
rect 20177 18785 20211 18819
rect 20545 18785 20579 18819
rect 20913 18785 20947 18819
rect 23213 18785 23247 18819
rect 25881 18785 25915 18819
rect 25973 18785 26007 18819
rect 27353 18785 27387 18819
rect 27721 18785 27755 18819
rect 28733 18785 28767 18819
rect 28917 18785 28951 18819
rect 29009 18785 29043 18819
rect 29193 18785 29227 18819
rect 29377 18785 29411 18819
rect 31125 18785 31159 18819
rect 3893 18717 3927 18751
rect 4353 18717 4387 18751
rect 4813 18717 4847 18751
rect 6285 18717 6319 18751
rect 6469 18717 6503 18751
rect 7113 18717 7147 18751
rect 9597 18717 9631 18751
rect 9873 18717 9907 18751
rect 16129 18717 16163 18751
rect 19717 18717 19751 18751
rect 20269 18717 20303 18751
rect 20453 18717 20487 18751
rect 21281 18717 21315 18751
rect 24200 18717 24234 18751
rect 24685 18717 24719 18751
rect 26985 18717 27019 18751
rect 27838 18717 27872 18751
rect 3709 18649 3743 18683
rect 4169 18649 4203 18683
rect 5181 18649 5215 18683
rect 5457 18649 5491 18683
rect 6561 18649 6595 18683
rect 6745 18649 6779 18683
rect 8493 18649 8527 18683
rect 9229 18649 9263 18683
rect 9413 18649 9447 18683
rect 14105 18649 14139 18683
rect 14289 18649 14323 18683
rect 17509 18649 17543 18683
rect 20821 18649 20855 18683
rect 22753 18649 22787 18683
rect 26525 18649 26559 18683
rect 27997 18649 28031 18683
rect 29745 18649 29779 18683
rect 4261 18581 4295 18615
rect 5089 18581 5123 18615
rect 6653 18581 6687 18615
rect 8953 18581 8987 18615
rect 9781 18581 9815 18615
rect 10517 18581 10551 18615
rect 13369 18581 13403 18615
rect 17601 18581 17635 18615
rect 18889 18581 18923 18615
rect 20545 18581 20579 18615
rect 20913 18581 20947 18615
rect 22661 18581 22695 18615
rect 25329 18581 25363 18615
rect 25513 18581 25547 18615
rect 26157 18581 26191 18615
rect 27261 18581 27295 18615
rect 29561 18581 29595 18615
rect 4997 18377 5031 18411
rect 10241 18377 10275 18411
rect 10701 18377 10735 18411
rect 12265 18377 12299 18411
rect 18429 18377 18463 18411
rect 18981 18377 19015 18411
rect 19993 18377 20027 18411
rect 20637 18377 20671 18411
rect 26525 18377 26559 18411
rect 26985 18377 27019 18411
rect 28733 18377 28767 18411
rect 5641 18309 5675 18343
rect 9965 18309 9999 18343
rect 10057 18309 10091 18343
rect 10333 18309 10367 18343
rect 19165 18309 19199 18343
rect 20269 18309 20303 18343
rect 22753 18309 22787 18343
rect 23029 18309 23063 18343
rect 26249 18309 26283 18343
rect 27353 18309 27387 18343
rect 28641 18309 28675 18343
rect 29285 18309 29319 18343
rect 4445 18241 4479 18275
rect 4629 18241 4663 18275
rect 5365 18241 5399 18275
rect 10149 18241 10183 18275
rect 22293 18241 22327 18275
rect 22845 18241 22879 18275
rect 26893 18241 26927 18275
rect 28825 18241 28859 18275
rect 4353 18173 4387 18207
rect 4721 18173 4755 18207
rect 4813 18173 4847 18207
rect 4997 18173 5031 18207
rect 5457 18173 5491 18207
rect 6193 18173 6227 18207
rect 6285 18173 6319 18207
rect 6469 18173 6503 18207
rect 7021 18173 7055 18207
rect 7389 18173 7423 18207
rect 7481 18173 7515 18207
rect 10057 18173 10091 18207
rect 10425 18173 10459 18207
rect 10517 18173 10551 18207
rect 10701 18173 10735 18207
rect 10885 18173 10919 18207
rect 11141 18173 11175 18207
rect 12357 18173 12391 18207
rect 13553 18173 13587 18207
rect 18245 18173 18279 18207
rect 18889 18173 18923 18207
rect 18981 18173 19015 18207
rect 19073 18173 19107 18207
rect 19441 18173 19475 18207
rect 19619 18173 19653 18207
rect 20545 18173 20579 18207
rect 20637 18173 20671 18207
rect 20913 18173 20947 18207
rect 21097 18173 21131 18207
rect 22201 18173 22235 18207
rect 22385 18173 22419 18207
rect 22661 18173 22695 18207
rect 22753 18173 22787 18207
rect 23121 18173 23155 18207
rect 23397 18173 23431 18207
rect 24225 18173 24259 18207
rect 24593 18173 24627 18207
rect 24961 18173 24995 18207
rect 26065 18173 26099 18207
rect 26801 18173 26835 18207
rect 27261 18173 27295 18207
rect 27537 18173 27571 18207
rect 28549 18173 28583 18207
rect 29193 18173 29227 18207
rect 29285 18173 29319 18207
rect 29561 18173 29595 18207
rect 29817 18173 29851 18207
rect 7205 18105 7239 18139
rect 9781 18105 9815 18139
rect 13798 18105 13832 18139
rect 18705 18105 18739 18139
rect 19349 18105 19383 18139
rect 19533 18105 19567 18139
rect 21005 18105 21039 18139
rect 22477 18105 22511 18139
rect 29009 18105 29043 18139
rect 4721 18037 4755 18071
rect 6377 18037 6411 18071
rect 6837 18037 6871 18071
rect 7665 18037 7699 18071
rect 12541 18037 12575 18071
rect 14933 18037 14967 18071
rect 19073 18037 19107 18071
rect 23121 18037 23155 18071
rect 23213 18037 23247 18071
rect 24225 18037 24259 18071
rect 27169 18037 27203 18071
rect 30941 18037 30975 18071
rect 5457 17833 5491 17867
rect 5917 17833 5951 17867
rect 9597 17833 9631 17867
rect 10977 17833 11011 17867
rect 14749 17833 14783 17867
rect 18797 17833 18831 17867
rect 19625 17833 19659 17867
rect 25329 17833 25363 17867
rect 26709 17833 26743 17867
rect 27353 17833 27387 17867
rect 29101 17833 29135 17867
rect 29469 17833 29503 17867
rect 4813 17765 4847 17799
rect 6285 17765 6319 17799
rect 7113 17765 7147 17799
rect 7748 17765 7782 17799
rect 9321 17765 9355 17799
rect 13001 17765 13035 17799
rect 17224 17765 17258 17799
rect 19533 17765 19567 17799
rect 20085 17765 20119 17799
rect 23204 17765 23238 17799
rect 24685 17765 24719 17799
rect 27169 17765 27203 17799
rect 27629 17765 27663 17799
rect 28089 17765 28123 17799
rect 29920 17765 29954 17799
rect 1593 17697 1627 17731
rect 4261 17697 4295 17731
rect 4445 17697 4479 17731
rect 4721 17697 4755 17731
rect 4997 17697 5031 17731
rect 5089 17697 5123 17731
rect 5457 17697 5491 17731
rect 5825 17697 5859 17731
rect 6009 17697 6043 17731
rect 6193 17697 6227 17731
rect 6377 17697 6411 17731
rect 7021 17697 7055 17731
rect 7389 17697 7423 17731
rect 7481 17697 7515 17731
rect 9137 17697 9171 17731
rect 9229 17697 9263 17731
rect 9413 17697 9447 17731
rect 9505 17697 9539 17731
rect 9701 17697 9735 17731
rect 10149 17697 10183 17731
rect 10517 17697 10551 17731
rect 10609 17697 10643 17731
rect 10977 17697 11011 17731
rect 11345 17697 11379 17731
rect 11529 17697 11563 17731
rect 12817 17697 12851 17731
rect 13093 17697 13127 17731
rect 13185 17697 13219 17731
rect 13461 17697 13495 17731
rect 15853 17697 15887 17731
rect 16957 17697 16991 17731
rect 18705 17697 18739 17731
rect 18889 17697 18923 17731
rect 19257 17697 19291 17731
rect 19349 17697 19383 17731
rect 19625 17697 19659 17731
rect 19993 17697 20027 17731
rect 20177 17697 20211 17731
rect 20269 17697 20303 17731
rect 20453 17697 20487 17731
rect 20545 17697 20579 17731
rect 20913 17697 20947 17731
rect 22937 17697 22971 17731
rect 24777 17697 24811 17731
rect 25789 17697 25823 17731
rect 29009 17697 29043 17731
rect 29193 17697 29227 17731
rect 29377 17697 29411 17731
rect 29561 17697 29595 17731
rect 5181 17629 5215 17663
rect 6745 17629 6779 17663
rect 7297 17629 7331 17663
rect 10333 17629 10367 17663
rect 11253 17629 11287 17663
rect 11437 17629 11471 17663
rect 13553 17629 13587 17663
rect 14841 17629 14875 17663
rect 15025 17629 15059 17663
rect 19901 17629 19935 17663
rect 20361 17629 20395 17663
rect 24568 17629 24602 17663
rect 25053 17629 25087 17663
rect 26617 17629 26651 17663
rect 27537 17629 27571 17663
rect 29653 17629 29687 17663
rect 4445 17561 4479 17595
rect 5089 17561 5123 17595
rect 5365 17561 5399 17595
rect 6929 17561 6963 17595
rect 8861 17561 8895 17595
rect 10609 17561 10643 17595
rect 11069 17561 11103 17595
rect 13369 17561 13403 17595
rect 19717 17561 19751 17595
rect 24317 17561 24351 17595
rect 26433 17561 26467 17595
rect 27169 17561 27203 17595
rect 28089 17561 28123 17595
rect 1409 17493 1443 17527
rect 4537 17493 4571 17527
rect 6653 17493 6687 17527
rect 6837 17493 6871 17527
rect 7205 17493 7239 17527
rect 9873 17493 9907 17527
rect 13461 17493 13495 17527
rect 13829 17493 13863 17527
rect 14381 17493 14415 17527
rect 15669 17493 15703 17527
rect 18337 17493 18371 17527
rect 19257 17493 19291 17527
rect 21097 17493 21131 17527
rect 24409 17493 24443 17527
rect 25697 17493 25731 17527
rect 31033 17493 31067 17527
rect 6837 17289 6871 17323
rect 10149 17289 10183 17323
rect 13277 17289 13311 17323
rect 14749 17289 14783 17323
rect 15117 17289 15151 17323
rect 18153 17289 18187 17323
rect 24501 17289 24535 17323
rect 27445 17289 27479 17323
rect 29469 17289 29503 17323
rect 4629 17221 4663 17255
rect 10057 17221 10091 17255
rect 10333 17221 10367 17255
rect 12357 17221 12391 17255
rect 24317 17221 24351 17255
rect 5089 17153 5123 17187
rect 10609 17153 10643 17187
rect 14565 17153 14599 17187
rect 16589 17153 16623 17187
rect 17325 17153 17359 17187
rect 26065 17153 26099 17187
rect 27077 17153 27111 17187
rect 1225 17085 1259 17119
rect 3249 17085 3283 17119
rect 4813 17085 4847 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 7297 17085 7331 17119
rect 7573 17085 7607 17119
rect 8401 17085 8435 17119
rect 9965 17085 9999 17119
rect 10333 17085 10367 17119
rect 10425 17085 10459 17119
rect 10701 17085 10735 17119
rect 10977 17085 11011 17119
rect 12725 17085 12759 17119
rect 13001 17085 13035 17119
rect 13093 17085 13127 17119
rect 13829 17085 13863 17119
rect 14013 17085 14047 17119
rect 14381 17085 14415 17119
rect 16230 17085 16264 17119
rect 16497 17085 16531 17119
rect 17233 17085 17267 17119
rect 17601 17085 17635 17119
rect 17785 17085 17819 17119
rect 18061 17085 18095 17119
rect 18245 17085 18279 17119
rect 18521 17085 18555 17119
rect 18889 17085 18923 17119
rect 19073 17085 19107 17119
rect 19257 17085 19291 17119
rect 19533 17085 19567 17119
rect 19993 17085 20027 17119
rect 20269 17085 20303 17119
rect 21741 17085 21775 17119
rect 26341 17085 26375 17119
rect 26801 17085 26835 17119
rect 26985 17085 27019 17119
rect 28825 17085 28859 17119
rect 29009 17085 29043 17119
rect 29101 17085 29135 17119
rect 29745 17085 29779 17119
rect 1501 17017 1535 17051
rect 3494 17017 3528 17051
rect 5334 17017 5368 17051
rect 8646 17017 8680 17051
rect 10241 17017 10275 17051
rect 11222 17017 11256 17051
rect 12909 17017 12943 17051
rect 18981 17017 19015 17051
rect 20514 17017 20548 17051
rect 21986 17017 22020 17051
rect 24869 17017 24903 17051
rect 27261 17017 27295 17051
rect 28558 17017 28592 17051
rect 29285 17017 29319 17051
rect 2973 16949 3007 16983
rect 4997 16949 5031 16983
rect 6469 16949 6503 16983
rect 7113 16949 7147 16983
rect 7757 16949 7791 16983
rect 9781 16949 9815 16983
rect 10885 16949 10919 16983
rect 17877 16949 17911 16983
rect 18337 16949 18371 16983
rect 18705 16949 18739 16983
rect 19349 16949 19383 16983
rect 20177 16949 20211 16983
rect 21649 16949 21683 16983
rect 23121 16949 23155 16983
rect 24492 16949 24526 16983
rect 26893 16949 26927 16983
rect 29009 16949 29043 16983
rect 29929 16949 29963 16983
rect 2329 16745 2363 16779
rect 4905 16745 4939 16779
rect 7205 16745 7239 16779
rect 10333 16745 10367 16779
rect 10517 16745 10551 16779
rect 13921 16745 13955 16779
rect 14841 16745 14875 16779
rect 15945 16745 15979 16779
rect 17785 16745 17819 16779
rect 23949 16745 23983 16779
rect 25053 16745 25087 16779
rect 27629 16745 27663 16779
rect 28089 16745 28123 16779
rect 28917 16745 28951 16779
rect 29653 16745 29687 16779
rect 31309 16745 31343 16779
rect 19064 16677 19098 16711
rect 21833 16677 21867 16711
rect 21925 16677 21959 16711
rect 22845 16677 22879 16711
rect 22937 16677 22971 16711
rect 24409 16677 24443 16711
rect 25973 16677 26007 16711
rect 27353 16677 27387 16711
rect 30174 16677 30208 16711
rect 1225 16609 1259 16643
rect 2421 16609 2455 16643
rect 2697 16609 2731 16643
rect 3525 16609 3559 16643
rect 3792 16609 3826 16643
rect 7205 16609 7239 16643
rect 7573 16609 7607 16643
rect 7665 16609 7699 16643
rect 10149 16609 10183 16643
rect 10425 16609 10459 16643
rect 10609 16609 10643 16643
rect 10977 16609 11011 16643
rect 12909 16609 12943 16643
rect 13093 16609 13127 16643
rect 13185 16609 13219 16643
rect 13277 16609 13311 16643
rect 13553 16609 13587 16643
rect 13737 16609 13771 16643
rect 14933 16609 14967 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 16672 16609 16706 16643
rect 18061 16609 18095 16643
rect 18153 16609 18187 16643
rect 18245 16609 18279 16643
rect 18429 16609 18463 16643
rect 21649 16609 21683 16643
rect 22017 16609 22051 16643
rect 22753 16609 22787 16643
rect 23121 16609 23155 16643
rect 23213 16609 23247 16643
rect 23673 16609 23707 16643
rect 24225 16609 24259 16643
rect 24317 16609 24351 16643
rect 24593 16609 24627 16643
rect 24777 16609 24811 16643
rect 25232 16609 25266 16643
rect 25329 16609 25363 16643
rect 25421 16609 25455 16643
rect 25549 16609 25583 16643
rect 25697 16609 25731 16643
rect 26617 16609 26651 16643
rect 26709 16609 26743 16643
rect 26893 16609 26927 16643
rect 27261 16609 27295 16643
rect 27629 16615 27663 16649
rect 27997 16609 28031 16643
rect 28273 16609 28307 16643
rect 28917 16609 28951 16643
rect 29285 16609 29319 16643
rect 29469 16609 29503 16643
rect 29561 16609 29595 16643
rect 29745 16609 29779 16643
rect 29929 16609 29963 16643
rect 1317 16541 1351 16575
rect 1593 16541 1627 16575
rect 7481 16541 7515 16575
rect 7849 16541 7883 16575
rect 16405 16541 16439 16575
rect 18797 16541 18831 16575
rect 26801 16541 26835 16575
rect 26985 16541 27019 16575
rect 27169 16541 27203 16575
rect 28825 16541 28859 16575
rect 29193 16541 29227 16575
rect 29377 16541 29411 16575
rect 7297 16473 7331 16507
rect 7573 16473 7607 16507
rect 13461 16473 13495 16507
rect 17877 16473 17911 16507
rect 25789 16473 25823 16507
rect 27261 16473 27295 16507
rect 27537 16473 27571 16507
rect 27813 16473 27847 16507
rect 29009 16473 29043 16507
rect 2605 16405 2639 16439
rect 15669 16405 15703 16439
rect 20177 16405 20211 16439
rect 22201 16405 22235 16439
rect 22569 16405 22603 16439
rect 23857 16405 23891 16439
rect 24225 16405 24259 16439
rect 4721 16201 4755 16235
rect 8033 16201 8067 16235
rect 10149 16201 10183 16235
rect 13369 16201 13403 16235
rect 16129 16201 16163 16235
rect 16773 16201 16807 16235
rect 17969 16201 18003 16235
rect 20821 16201 20855 16235
rect 21097 16201 21131 16235
rect 22293 16201 22327 16235
rect 25513 16201 25547 16235
rect 29009 16201 29043 16235
rect 7941 16133 7975 16167
rect 12633 16133 12667 16167
rect 26709 16133 26743 16167
rect 28549 16133 28583 16167
rect 1317 16065 1351 16099
rect 6561 16065 6595 16099
rect 8769 16065 8803 16099
rect 16037 16065 16071 16099
rect 21741 16065 21775 16099
rect 30389 16065 30423 16099
rect 1041 15997 1075 16031
rect 1225 15997 1259 16031
rect 3341 15997 3375 16031
rect 4997 15997 5031 16031
rect 6828 15997 6862 16031
rect 8033 15997 8067 16031
rect 8217 15997 8251 16031
rect 9036 15997 9070 16031
rect 10241 15997 10275 16031
rect 10497 15997 10531 16031
rect 12081 15997 12115 16031
rect 12357 15997 12391 16031
rect 12449 15997 12483 16031
rect 12725 15997 12759 16031
rect 12818 15997 12852 16031
rect 13001 15997 13035 16031
rect 13231 15997 13265 16031
rect 13829 15997 13863 16031
rect 13922 15997 13956 16031
rect 14335 15997 14369 16031
rect 15209 15997 15243 16031
rect 15347 15997 15381 16031
rect 15485 15997 15519 16031
rect 16313 15997 16347 16031
rect 16405 15997 16439 16031
rect 16497 15997 16531 16031
rect 16681 15997 16715 16031
rect 16957 15997 16991 16031
rect 17233 15997 17267 16031
rect 17693 15997 17727 16031
rect 18153 15997 18187 16031
rect 18429 15997 18463 16031
rect 20085 15997 20119 16031
rect 20177 15997 20211 16031
rect 20545 15997 20579 16031
rect 20637 15997 20671 16031
rect 21465 15997 21499 16031
rect 22472 15997 22506 16031
rect 22661 15997 22695 16031
rect 22844 15997 22878 16031
rect 22937 15997 22971 16031
rect 23213 15997 23247 16031
rect 23581 15997 23615 16031
rect 24133 15997 24167 16031
rect 28089 15997 28123 16031
rect 28273 15997 28307 16031
rect 30122 15997 30156 16031
rect 1133 15929 1167 15963
rect 1593 15929 1627 15963
rect 3586 15929 3620 15963
rect 5242 15929 5276 15963
rect 12265 15929 12299 15963
rect 13093 15929 13127 15963
rect 14105 15929 14139 15963
rect 14197 15929 14231 15963
rect 20315 15929 20349 15963
rect 20453 15929 20487 15963
rect 20913 15929 20947 15963
rect 21129 15929 21163 15963
rect 22569 15929 22603 15963
rect 23305 15929 23339 15963
rect 23397 15929 23431 15963
rect 24389 15929 24423 15963
rect 27822 15929 27856 15963
rect 28733 15929 28767 15963
rect 3065 15861 3099 15895
rect 6377 15861 6411 15895
rect 11621 15861 11655 15895
rect 14473 15861 14507 15895
rect 17141 15861 17175 15895
rect 17509 15861 17543 15895
rect 18337 15861 18371 15895
rect 19901 15861 19935 15895
rect 21281 15861 21315 15895
rect 23029 15861 23063 15895
rect 28457 15861 28491 15895
rect 1501 15657 1535 15691
rect 2237 15657 2271 15691
rect 3801 15657 3835 15691
rect 7389 15657 7423 15691
rect 8033 15657 8067 15691
rect 9505 15657 9539 15691
rect 10701 15657 10735 15691
rect 14289 15657 14323 15691
rect 18521 15657 18555 15691
rect 20269 15657 20303 15691
rect 21649 15657 21683 15691
rect 27169 15657 27203 15691
rect 27997 15657 28031 15691
rect 31309 15657 31343 15691
rect 1777 15589 1811 15623
rect 8370 15589 8404 15623
rect 9781 15589 9815 15623
rect 11222 15589 11256 15623
rect 24041 15589 24075 15623
rect 24133 15589 24167 15623
rect 25982 15589 26016 15623
rect 30174 15589 30208 15623
rect 1685 15521 1719 15555
rect 1869 15521 1903 15555
rect 2145 15521 2179 15555
rect 2421 15521 2455 15555
rect 2513 15521 2547 15555
rect 3617 15521 3651 15555
rect 3893 15521 3927 15555
rect 5089 15521 5123 15555
rect 5365 15521 5399 15555
rect 7297 15521 7331 15555
rect 7481 15521 7515 15555
rect 7573 15521 7607 15555
rect 7849 15521 7883 15555
rect 9597 15521 9631 15555
rect 10517 15521 10551 15555
rect 12996 15521 13030 15555
rect 13093 15521 13127 15555
rect 13185 15521 13219 15555
rect 13313 15521 13347 15555
rect 13461 15521 13495 15555
rect 13553 15521 13587 15555
rect 13737 15521 13771 15555
rect 13829 15521 13863 15555
rect 13921 15521 13955 15555
rect 14197 15521 14231 15555
rect 14473 15521 14507 15555
rect 17601 15521 17635 15555
rect 17785 15521 17819 15555
rect 18153 15521 18187 15555
rect 19145 15521 19179 15555
rect 21373 15521 21407 15555
rect 21465 15521 21499 15555
rect 22293 15521 22327 15555
rect 22477 15521 22511 15555
rect 23857 15521 23891 15555
rect 24225 15521 24259 15555
rect 26249 15521 26283 15555
rect 26985 15521 27019 15555
rect 29110 15521 29144 15555
rect 29469 15521 29503 15555
rect 2329 15453 2363 15487
rect 8125 15453 8159 15487
rect 10977 15453 11011 15487
rect 16129 15453 16163 15487
rect 16405 15453 16439 15487
rect 18337 15453 18371 15487
rect 18889 15453 18923 15487
rect 29377 15453 29411 15487
rect 29929 15453 29963 15487
rect 2053 15385 2087 15419
rect 14105 15385 14139 15419
rect 22661 15385 22695 15419
rect 24409 15385 24443 15419
rect 3433 15317 3467 15351
rect 5273 15317 5307 15351
rect 5549 15317 5583 15351
rect 12357 15317 12391 15351
rect 12817 15317 12851 15351
rect 14657 15317 14691 15351
rect 22293 15317 22327 15351
rect 24869 15317 24903 15351
rect 5089 15113 5123 15147
rect 10793 15113 10827 15147
rect 12265 15113 12299 15147
rect 15209 15113 15243 15147
rect 15485 15113 15519 15147
rect 17693 15113 17727 15147
rect 25237 15113 25271 15147
rect 27261 15113 27295 15147
rect 7849 15045 7883 15079
rect 8585 15045 8619 15079
rect 15025 15045 15059 15079
rect 16957 15045 16991 15079
rect 19349 15045 19383 15079
rect 27169 15045 27203 15079
rect 5457 14977 5491 15011
rect 8125 14977 8159 15011
rect 15209 14977 15243 15011
rect 20361 14977 20395 15011
rect 28641 14977 28675 15011
rect 2881 14909 2915 14943
rect 3065 14909 3099 14943
rect 3341 14909 3375 14943
rect 5713 14909 5747 14943
rect 7305 14909 7339 14943
rect 7573 14909 7607 14943
rect 7757 14909 7791 14943
rect 7849 14909 7883 14943
rect 7941 14909 7975 14943
rect 8677 14909 8711 14943
rect 8769 14909 8803 14943
rect 8965 14909 8999 14943
rect 9137 14909 9171 14943
rect 9413 14909 9447 14943
rect 10885 14909 10919 14943
rect 13553 14909 13587 14943
rect 13646 14909 13680 14943
rect 13829 14909 13863 14943
rect 14059 14909 14093 14943
rect 14381 14909 14415 14943
rect 14474 14909 14508 14943
rect 14657 14909 14691 14943
rect 14846 14909 14880 14943
rect 15117 14909 15151 14943
rect 15577 14909 15611 14943
rect 17049 14909 17083 14943
rect 17142 14909 17176 14943
rect 17514 14909 17548 14943
rect 18705 14909 18739 14943
rect 18853 14909 18887 14943
rect 19211 14909 19245 14943
rect 20085 14909 20119 14943
rect 22753 14909 22787 14943
rect 22845 14909 22879 14943
rect 22937 14909 22971 14943
rect 23121 14909 23155 14943
rect 23213 14909 23247 14943
rect 23857 14909 23891 14943
rect 25789 14909 25823 14943
rect 3617 14841 3651 14875
rect 7665 14841 7699 14875
rect 8401 14841 8435 14875
rect 8861 14841 8895 14875
rect 9658 14841 9692 14875
rect 11130 14841 11164 14875
rect 13921 14841 13955 14875
rect 14749 14841 14783 14875
rect 15822 14841 15856 14875
rect 17325 14841 17359 14875
rect 17417 14841 17451 14875
rect 18981 14841 19015 14875
rect 19073 14841 19107 14875
rect 20606 14841 20640 14875
rect 24102 14841 24136 14875
rect 26056 14841 26090 14875
rect 28396 14841 28430 14875
rect 3065 14773 3099 14807
rect 6837 14773 6871 14807
rect 7481 14773 7515 14807
rect 8677 14773 8711 14807
rect 9321 14773 9355 14807
rect 14197 14773 14231 14807
rect 20269 14773 20303 14807
rect 21741 14773 21775 14807
rect 22569 14773 22603 14807
rect 23397 14773 23431 14807
rect 3433 14569 3467 14603
rect 4445 14569 4479 14603
rect 8953 14569 8987 14603
rect 9413 14569 9447 14603
rect 13001 14569 13035 14603
rect 13645 14569 13679 14603
rect 14289 14569 14323 14603
rect 15669 14569 15703 14603
rect 17509 14569 17543 14603
rect 19165 14569 19199 14603
rect 21281 14569 21315 14603
rect 21925 14569 21959 14603
rect 22109 14569 22143 14603
rect 24317 14569 24351 14603
rect 31309 14569 31343 14603
rect 3157 14501 3191 14535
rect 7818 14501 7852 14535
rect 13369 14501 13403 14535
rect 16374 14501 16408 14535
rect 19502 14501 19536 14535
rect 22385 14501 22419 14535
rect 28825 14501 28859 14535
rect 29101 14501 29135 14535
rect 30174 14501 30208 14535
rect 1133 14433 1167 14467
rect 3249 14433 3283 14467
rect 3617 14433 3651 14467
rect 3801 14433 3835 14467
rect 4353 14433 4387 14467
rect 5825 14433 5859 14467
rect 6092 14433 6126 14467
rect 7573 14433 7607 14467
rect 9229 14433 9263 14467
rect 9505 14433 9539 14467
rect 9873 14433 9907 14467
rect 10517 14433 10551 14467
rect 10701 14433 10735 14467
rect 11161 14433 11195 14467
rect 11437 14433 11471 14467
rect 11621 14433 11655 14467
rect 12449 14433 12483 14467
rect 12633 14433 12667 14467
rect 12725 14433 12759 14467
rect 12817 14433 12851 14467
rect 13093 14433 13127 14467
rect 13277 14433 13311 14467
rect 13461 14433 13495 14467
rect 13737 14433 13771 14467
rect 13921 14433 13955 14467
rect 14013 14433 14047 14467
rect 14105 14433 14139 14467
rect 15485 14433 15519 14467
rect 16129 14433 16163 14467
rect 18981 14433 19015 14467
rect 19257 14433 19291 14467
rect 21649 14433 21683 14467
rect 22017 14433 22051 14467
rect 22293 14433 22327 14467
rect 22477 14433 22511 14467
rect 22661 14433 22695 14467
rect 25441 14433 25475 14467
rect 26617 14433 26651 14467
rect 29009 14433 29043 14467
rect 29193 14433 29227 14467
rect 29377 14433 29411 14467
rect 29653 14433 29687 14467
rect 1409 14365 1443 14399
rect 3893 14365 3927 14399
rect 9781 14365 9815 14399
rect 10149 14365 10183 14399
rect 10609 14365 10643 14399
rect 21557 14365 21591 14399
rect 25697 14365 25731 14399
rect 26709 14365 26743 14399
rect 29929 14365 29963 14399
rect 7205 14297 7239 14331
rect 9597 14297 9631 14331
rect 9873 14297 9907 14331
rect 9965 14297 9999 14331
rect 11437 14297 11471 14331
rect 2881 14229 2915 14263
rect 9505 14229 9539 14263
rect 10241 14229 10275 14263
rect 11345 14229 11379 14263
rect 20637 14229 20671 14263
rect 21741 14229 21775 14263
rect 26985 14229 27019 14263
rect 29561 14229 29595 14263
rect 1409 14025 1443 14059
rect 8401 14025 8435 14059
rect 9781 14025 9815 14059
rect 12725 14025 12759 14059
rect 16037 14025 16071 14059
rect 18245 14025 18279 14059
rect 21189 14025 21223 14059
rect 23581 14025 23615 14059
rect 24225 14025 24259 14059
rect 26065 14025 26099 14059
rect 26801 14025 26835 14059
rect 28641 14025 28675 14059
rect 7021 13957 7055 13991
rect 10885 13957 10919 13991
rect 14381 13957 14415 13991
rect 28825 13957 28859 13991
rect 1133 13889 1167 13923
rect 5641 13889 5675 13923
rect 10241 13889 10275 13923
rect 10425 13889 10459 13923
rect 11069 13889 11103 13923
rect 22201 13889 22235 13923
rect 24593 13889 24627 13923
rect 1041 13821 1075 13855
rect 3985 13821 4019 13855
rect 4169 13821 4203 13855
rect 4261 13821 4295 13855
rect 9597 13821 9631 13855
rect 9781 13821 9815 13855
rect 10057 13821 10091 13855
rect 10149 13821 10183 13855
rect 10333 13821 10367 13855
rect 10609 13821 10643 13855
rect 10701 13821 10735 13855
rect 10793 13821 10827 13855
rect 11345 13821 11379 13855
rect 11601 13821 11635 13855
rect 14197 13821 14231 13855
rect 14657 13821 14691 13855
rect 14913 13821 14947 13855
rect 16865 13821 16899 13855
rect 20637 13821 20671 13855
rect 20913 13821 20947 13855
rect 21005 13821 21039 13855
rect 23949 13821 23983 13855
rect 24041 13821 24075 13855
rect 24225 13821 24259 13855
rect 24317 13821 24351 13855
rect 26709 13821 26743 13855
rect 29193 13821 29227 13855
rect 5908 13753 5942 13787
rect 17132 13753 17166 13787
rect 20821 13753 20855 13787
rect 22446 13753 22480 13787
rect 28457 13753 28491 13787
rect 29469 13753 29503 13787
rect 3801 13685 3835 13719
rect 10701 13685 10735 13719
rect 10793 13685 10827 13719
rect 28667 13685 28701 13719
rect 30941 13685 30975 13719
rect 5181 13481 5215 13515
rect 6009 13481 6043 13515
rect 7941 13481 7975 13515
rect 11253 13481 11287 13515
rect 14105 13481 14139 13515
rect 15577 13481 15611 13515
rect 18889 13481 18923 13515
rect 21925 13481 21959 13515
rect 25329 13481 25363 13515
rect 25605 13481 25639 13515
rect 26525 13481 26559 13515
rect 28457 13481 28491 13515
rect 28825 13481 28859 13515
rect 29469 13481 29503 13515
rect 30297 13481 30331 13515
rect 3065 13413 3099 13447
rect 3709 13413 3743 13447
rect 6193 13413 6227 13447
rect 14442 13413 14476 13447
rect 17776 13413 17810 13447
rect 24685 13413 24719 13447
rect 27997 13413 28031 13447
rect 1133 13345 1167 13379
rect 3157 13345 3191 13379
rect 6101 13345 6135 13379
rect 6817 13345 6851 13379
rect 8289 13345 8323 13379
rect 11069 13345 11103 13379
rect 12992 13345 13026 13379
rect 14197 13345 14231 13379
rect 17509 13345 17543 13379
rect 19533 13345 19567 13379
rect 21465 13345 21499 13379
rect 23049 13345 23083 13379
rect 24501 13345 24535 13379
rect 24961 13345 24995 13379
rect 25237 13345 25271 13379
rect 25421 13345 25455 13379
rect 25697 13345 25731 13379
rect 28273 13345 28307 13379
rect 28549 13345 28583 13379
rect 28733 13345 28767 13379
rect 29009 13345 29043 13379
rect 29101 13345 29135 13379
rect 29285 13345 29319 13379
rect 29377 13345 29411 13379
rect 29561 13345 29595 13379
rect 30205 13345 30239 13379
rect 1409 13277 1443 13311
rect 3433 13277 3467 13311
rect 6561 13277 6595 13311
rect 8033 13277 8067 13311
rect 12725 13277 12759 13311
rect 19441 13277 19475 13311
rect 23305 13277 23339 13311
rect 24317 13277 24351 13311
rect 25145 13277 25179 13311
rect 6377 13209 6411 13243
rect 29009 13209 29043 13243
rect 2881 13141 2915 13175
rect 5825 13141 5859 13175
rect 9413 13141 9447 13175
rect 19901 13141 19935 13175
rect 21373 13141 21407 13175
rect 24777 13141 24811 13175
rect 29101 13141 29135 13175
rect 2881 12937 2915 12971
rect 3985 12937 4019 12971
rect 4445 12937 4479 12971
rect 5273 12937 5307 12971
rect 8217 12937 8251 12971
rect 13369 12937 13403 12971
rect 21833 12937 21867 12971
rect 22385 12937 22419 12971
rect 24777 12937 24811 12971
rect 30849 12937 30883 12971
rect 1041 12869 1075 12903
rect 2697 12869 2731 12903
rect 11897 12869 11931 12903
rect 17693 12869 17727 12903
rect 18337 12869 18371 12903
rect 23213 12869 23247 12903
rect 25513 12869 25547 12903
rect 1501 12801 1535 12835
rect 6837 12801 6871 12835
rect 8861 12801 8895 12835
rect 16129 12801 16163 12835
rect 18245 12801 18279 12835
rect 20361 12801 20395 12835
rect 25145 12801 25179 12835
rect 1409 12733 1443 12767
rect 3617 12733 3651 12767
rect 3709 12733 3743 12767
rect 4353 12733 4387 12767
rect 5181 12733 5215 12767
rect 5365 12733 5399 12767
rect 6009 12733 6043 12767
rect 10517 12733 10551 12767
rect 11989 12733 12023 12767
rect 15853 12733 15887 12767
rect 18337 12733 18371 12767
rect 18521 12733 18555 12767
rect 20085 12733 20119 12767
rect 22661 12733 22695 12767
rect 22937 12733 22971 12767
rect 23305 12733 23339 12767
rect 23489 12733 23523 12767
rect 23673 12733 23707 12767
rect 25053 12733 25087 12767
rect 25237 12733 25271 12767
rect 25329 12733 25363 12767
rect 25513 12733 25547 12767
rect 26157 12733 26191 12767
rect 26893 12733 26927 12767
rect 28641 12733 28675 12767
rect 28825 12733 28859 12767
rect 29101 12733 29135 12767
rect 30941 12733 30975 12767
rect 3065 12665 3099 12699
rect 3433 12665 3467 12699
rect 5825 12665 5859 12699
rect 6377 12665 6411 12699
rect 7104 12665 7138 12699
rect 9106 12665 9140 12699
rect 10762 12665 10796 12699
rect 12256 12665 12290 12699
rect 22201 12665 22235 12699
rect 22401 12665 22435 12699
rect 23029 12665 23063 12699
rect 24593 12665 24627 12699
rect 28733 12665 28767 12699
rect 29377 12665 29411 12699
rect 31033 12665 31067 12699
rect 2865 12597 2899 12631
rect 3801 12597 3835 12631
rect 6101 12597 6135 12631
rect 6193 12597 6227 12631
rect 10241 12597 10275 12631
rect 17601 12597 17635 12631
rect 17877 12597 17911 12631
rect 17969 12597 18003 12631
rect 18061 12597 18095 12631
rect 22569 12597 22603 12631
rect 22845 12597 22879 12631
rect 24793 12597 24827 12631
rect 24961 12597 24995 12631
rect 25973 12597 26007 12631
rect 26985 12597 27019 12631
rect 3157 12393 3191 12427
rect 5181 12393 5215 12427
rect 5641 12393 5675 12427
rect 6929 12393 6963 12427
rect 12357 12393 12391 12427
rect 14473 12393 14507 12427
rect 15945 12393 15979 12427
rect 16957 12393 16991 12427
rect 17877 12393 17911 12427
rect 18061 12393 18095 12427
rect 20085 12393 20119 12427
rect 22661 12393 22695 12427
rect 26433 12393 26467 12427
rect 30757 12393 30791 12427
rect 3709 12325 3743 12359
rect 5273 12325 5307 12359
rect 5478 12325 5512 12359
rect 6193 12325 6227 12359
rect 18245 12325 18279 12359
rect 18950 12325 18984 12359
rect 23305 12325 23339 12359
rect 2329 12257 2363 12291
rect 2513 12257 2547 12291
rect 2789 12257 2823 12291
rect 7113 12257 7147 12291
rect 7297 12257 7331 12291
rect 9045 12257 9079 12291
rect 9229 12257 9263 12291
rect 9597 12257 9631 12291
rect 11233 12257 11267 12291
rect 13093 12257 13127 12291
rect 13360 12257 13394 12291
rect 14565 12257 14599 12291
rect 14832 12257 14866 12291
rect 17049 12257 17083 12291
rect 17417 12257 17451 12291
rect 17509 12257 17543 12291
rect 17693 12257 17727 12291
rect 17969 12257 18003 12291
rect 18337 12257 18371 12291
rect 21281 12257 21315 12291
rect 21548 12257 21582 12291
rect 24317 12257 24351 12291
rect 28457 12257 28491 12291
rect 2421 12189 2455 12223
rect 2697 12189 2731 12223
rect 3433 12189 3467 12223
rect 9413 12189 9447 12223
rect 10977 12189 11011 12223
rect 18153 12189 18187 12223
rect 18705 12189 18739 12223
rect 24593 12189 24627 12223
rect 27905 12189 27939 12223
rect 28181 12189 28215 12223
rect 28365 12189 28399 12223
rect 29009 12189 29043 12223
rect 29285 12189 29319 12223
rect 28825 12121 28859 12155
rect 5457 12053 5491 12087
rect 6101 12053 6135 12087
rect 9689 12053 9723 12087
rect 23397 12053 23431 12087
rect 26065 12053 26099 12087
rect 4629 11849 4663 11883
rect 6745 11849 6779 11883
rect 10425 11849 10459 11883
rect 14841 11849 14875 11883
rect 18521 11849 18555 11883
rect 20545 11849 20579 11883
rect 22845 11849 22879 11883
rect 24501 11849 24535 11883
rect 25513 11849 25547 11883
rect 30113 11849 30147 11883
rect 14105 11781 14139 11815
rect 8125 11713 8159 11747
rect 19165 11713 19199 11747
rect 26985 11713 27019 11747
rect 4721 11645 4755 11679
rect 5089 11645 5123 11679
rect 6009 11645 6043 11679
rect 6285 11645 6319 11679
rect 6469 11645 6503 11679
rect 7481 11645 7515 11679
rect 7665 11645 7699 11679
rect 7941 11645 7975 11679
rect 8401 11645 8435 11679
rect 8585 11645 8619 11679
rect 8677 11645 8711 11679
rect 10701 11645 10735 11679
rect 13829 11645 13863 11679
rect 14933 11645 14967 11679
rect 15301 11645 15335 11679
rect 15577 11645 15611 11679
rect 16129 11645 16163 11679
rect 16221 11645 16255 11679
rect 16773 11645 16807 11679
rect 18889 11645 18923 11679
rect 21465 11645 21499 11679
rect 24685 11645 24719 11679
rect 24961 11645 24995 11679
rect 25145 11645 25179 11679
rect 25605 11645 25639 11679
rect 26893 11645 26927 11679
rect 30021 11645 30055 11679
rect 5365 11577 5399 11611
rect 6929 11577 6963 11611
rect 7757 11577 7791 11611
rect 8493 11577 8527 11611
rect 8953 11577 8987 11611
rect 10609 11577 10643 11611
rect 11897 11577 11931 11611
rect 13553 11577 13587 11611
rect 13737 11577 13771 11611
rect 17049 11577 17083 11611
rect 18797 11577 18831 11611
rect 19432 11577 19466 11611
rect 20821 11577 20855 11611
rect 21189 11577 21223 11611
rect 21732 11577 21766 11611
rect 26801 11577 26835 11611
rect 27261 11577 27295 11611
rect 5825 11509 5859 11543
rect 6561 11509 6595 11543
rect 6729 11509 6763 11543
rect 7573 11509 7607 11543
rect 11805 11509 11839 11543
rect 13921 11509 13955 11543
rect 15485 11509 15519 11543
rect 15761 11509 15795 11543
rect 21005 11509 21039 11543
rect 21097 11509 21131 11543
rect 21373 11509 21407 11543
rect 28733 11509 28767 11543
rect 5089 11305 5123 11339
rect 8946 11305 8980 11339
rect 12909 11305 12943 11339
rect 13445 11305 13479 11339
rect 13829 11305 13863 11339
rect 16497 11305 16531 11339
rect 16773 11305 16807 11339
rect 17509 11305 17543 11339
rect 21557 11305 21591 11339
rect 21649 11305 21683 11339
rect 24317 11305 24351 11339
rect 28549 11305 28583 11339
rect 5365 11237 5399 11271
rect 6101 11237 6135 11271
rect 9045 11237 9079 11271
rect 13645 11237 13679 11271
rect 16681 11237 16715 11271
rect 22017 11237 22051 11271
rect 2881 11169 2915 11203
rect 5457 11169 5491 11203
rect 7665 11169 7699 11203
rect 7849 11169 7883 11203
rect 8769 11169 8803 11203
rect 8861 11169 8895 11203
rect 11161 11169 11195 11203
rect 13001 11169 13035 11203
rect 13185 11169 13219 11203
rect 15577 11169 15611 11203
rect 15761 11169 15795 11203
rect 16313 11169 16347 11203
rect 17693 11169 17727 11203
rect 18061 11169 18095 11203
rect 18245 11169 18279 11203
rect 20085 11169 20119 11203
rect 20361 11169 20395 11203
rect 21465 11169 21499 11203
rect 21925 11169 21959 11203
rect 22109 11169 22143 11203
rect 23204 11169 23238 11203
rect 25237 11169 25271 11203
rect 25421 11169 25455 11203
rect 25789 11169 25823 11203
rect 28181 11169 28215 11203
rect 28641 11169 28675 11203
rect 28917 11169 28951 11203
rect 2789 11101 2823 11135
rect 3341 11101 3375 11135
rect 3617 11101 3651 11135
rect 5825 11101 5859 11135
rect 11437 11101 11471 11135
rect 17969 11101 18003 11135
rect 22937 11101 22971 11135
rect 25329 11101 25363 11135
rect 25697 11101 25731 11135
rect 26433 11101 26467 11135
rect 27905 11101 27939 11135
rect 29101 11101 29135 11135
rect 3249 11033 3283 11067
rect 7573 11033 7607 11067
rect 13277 11033 13311 11067
rect 15945 11033 15979 11067
rect 17877 11033 17911 11067
rect 18153 11033 18187 11067
rect 20269 11033 20303 11067
rect 21281 11033 21315 11067
rect 21833 11033 21867 11067
rect 26157 11033 26191 11067
rect 7665 10965 7699 10999
rect 13185 10965 13219 10999
rect 13461 10965 13495 10999
rect 15313 10965 15347 10999
rect 19901 10965 19935 10999
rect 6193 10761 6227 10795
rect 8217 10761 8251 10795
rect 11621 10761 11655 10795
rect 12173 10761 12207 10795
rect 14105 10761 14139 10795
rect 14841 10761 14875 10795
rect 20545 10761 20579 10795
rect 23489 10761 23523 10795
rect 25697 10761 25731 10795
rect 27445 10761 27479 10795
rect 13829 10693 13863 10727
rect 6469 10625 6503 10659
rect 6745 10625 6779 10659
rect 8861 10625 8895 10659
rect 9321 10625 9355 10659
rect 9689 10625 9723 10659
rect 16405 10625 16439 10659
rect 19073 10625 19107 10659
rect 21189 10625 21223 10659
rect 21649 10625 21683 10659
rect 22017 10625 22051 10659
rect 23949 10625 23983 10659
rect 6101 10557 6135 10591
rect 8585 10557 8619 10591
rect 8953 10557 8987 10591
rect 9413 10557 9447 10591
rect 11437 10557 11471 10591
rect 11621 10557 11655 10591
rect 12081 10557 12115 10591
rect 13553 10557 13587 10591
rect 13921 10557 13955 10591
rect 14105 10557 14139 10591
rect 14933 10557 14967 10591
rect 18521 10557 18555 10591
rect 18797 10557 18831 10591
rect 21281 10557 21315 10591
rect 21741 10557 21775 10591
rect 26065 10557 26099 10591
rect 27537 10557 27571 10591
rect 8493 10489 8527 10523
rect 13829 10489 13863 10523
rect 16681 10489 16715 10523
rect 18429 10489 18463 10523
rect 24225 10489 24259 10523
rect 25973 10489 26007 10523
rect 11161 10421 11195 10455
rect 13645 10421 13679 10455
rect 18153 10421 18187 10455
rect 10517 10217 10551 10251
rect 15393 10217 15427 10251
rect 19809 10217 19843 10251
rect 21281 10217 21315 10251
rect 22937 10217 22971 10251
rect 13277 10149 13311 10183
rect 15669 10149 15703 10183
rect 17877 10149 17911 10183
rect 21449 10149 21483 10183
rect 21649 10149 21683 10183
rect 10425 10081 10459 10115
rect 11253 10081 11287 10115
rect 13645 10081 13679 10115
rect 15577 10081 15611 10115
rect 17141 10081 17175 10115
rect 19717 10081 19751 10115
rect 22845 10081 22879 10115
rect 23581 10081 23615 10115
rect 11529 10013 11563 10047
rect 13921 10013 13955 10047
rect 16773 10013 16807 10047
rect 17233 10013 17267 10047
rect 17601 10013 17635 10047
rect 23489 10013 23523 10047
rect 23949 10013 23983 10047
rect 21465 9877 21499 9911
rect 11989 9673 12023 9707
rect 14105 9673 14139 9707
rect 12357 9605 12391 9639
rect 13829 9537 13863 9571
rect 12081 9469 12115 9503
rect 12265 9469 12299 9503
rect 13737 9469 13771 9503
<< metal1 >>
rect 16298 21836 16304 21888
rect 16356 21876 16362 21888
rect 23934 21876 23940 21888
rect 16356 21848 23940 21876
rect 16356 21836 16362 21848
rect 23934 21836 23940 21848
rect 23992 21876 23998 21888
rect 29362 21876 29368 21888
rect 23992 21848 29368 21876
rect 23992 21836 23998 21848
rect 29362 21836 29368 21848
rect 29420 21836 29426 21888
rect 552 21786 31648 21808
rect 552 21734 4285 21786
rect 4337 21734 4349 21786
rect 4401 21734 4413 21786
rect 4465 21734 4477 21786
rect 4529 21734 4541 21786
rect 4593 21734 12059 21786
rect 12111 21734 12123 21786
rect 12175 21734 12187 21786
rect 12239 21734 12251 21786
rect 12303 21734 12315 21786
rect 12367 21734 19833 21786
rect 19885 21734 19897 21786
rect 19949 21734 19961 21786
rect 20013 21734 20025 21786
rect 20077 21734 20089 21786
rect 20141 21734 27607 21786
rect 27659 21734 27671 21786
rect 27723 21734 27735 21786
rect 27787 21734 27799 21786
rect 27851 21734 27863 21786
rect 27915 21734 31648 21786
rect 552 21712 31648 21734
rect 842 21632 848 21684
rect 900 21632 906 21684
rect 1578 21632 1584 21684
rect 1636 21632 1642 21684
rect 2314 21632 2320 21684
rect 2372 21632 2378 21684
rect 3234 21632 3240 21684
rect 3292 21632 3298 21684
rect 3786 21632 3792 21684
rect 3844 21632 3850 21684
rect 4525 21675 4583 21681
rect 4525 21641 4537 21675
rect 4571 21672 4583 21675
rect 4614 21672 4620 21684
rect 4571 21644 4620 21672
rect 4571 21641 4583 21644
rect 4525 21635 4583 21641
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 5258 21632 5264 21684
rect 5316 21632 5322 21684
rect 5994 21632 6000 21684
rect 6052 21632 6058 21684
rect 6730 21632 6736 21684
rect 6788 21632 6794 21684
rect 7466 21632 7472 21684
rect 7524 21632 7530 21684
rect 8202 21632 8208 21684
rect 8260 21632 8266 21684
rect 8754 21632 8760 21684
rect 8812 21632 8818 21684
rect 9674 21632 9680 21684
rect 9732 21632 9738 21684
rect 10410 21632 10416 21684
rect 10468 21632 10474 21684
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 16298 21672 16304 21684
rect 11256 21644 16304 21672
rect 11256 21604 11284 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 23934 21632 23940 21684
rect 23992 21632 23998 21684
rect 27154 21672 27160 21684
rect 25424 21644 27160 21672
rect 9416 21576 11284 21604
rect 12897 21607 12955 21613
rect 6638 21428 6644 21480
rect 6696 21468 6702 21480
rect 9416 21477 9444 21576
rect 12897 21573 12909 21607
rect 12943 21573 12955 21607
rect 12897 21567 12955 21573
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 6696 21440 9137 21468
rect 6696 21428 6702 21440
rect 9125 21437 9137 21440
rect 9171 21468 9183 21471
rect 9217 21471 9275 21477
rect 9217 21468 9229 21471
rect 9171 21440 9229 21468
rect 9171 21437 9183 21440
rect 9125 21431 9183 21437
rect 9217 21437 9229 21440
rect 9263 21437 9275 21471
rect 9217 21431 9275 21437
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21437 9459 21471
rect 9401 21431 9459 21437
rect 11514 21428 11520 21480
rect 11572 21468 11578 21480
rect 12912 21468 12940 21567
rect 14642 21564 14648 21616
rect 14700 21604 14706 21616
rect 16209 21607 16267 21613
rect 16209 21604 16221 21607
rect 14700 21576 16221 21604
rect 14700 21564 14706 21576
rect 16209 21573 16221 21576
rect 16255 21573 16267 21607
rect 23014 21604 23020 21616
rect 16209 21567 16267 21573
rect 22848 21576 23020 21604
rect 14366 21496 14372 21548
rect 14424 21496 14430 21548
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 16666 21536 16672 21548
rect 14599 21508 16672 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 21729 21539 21787 21545
rect 21729 21536 21741 21539
rect 21008 21508 21741 21536
rect 21008 21480 21036 21508
rect 21729 21505 21741 21508
rect 21775 21505 21787 21539
rect 21729 21499 21787 21505
rect 14645 21471 14703 21477
rect 14645 21468 14657 21471
rect 11572 21440 12848 21468
rect 12912 21440 14657 21468
rect 11572 21428 11578 21440
rect 11422 21360 11428 21412
rect 11480 21400 11486 21412
rect 11762 21403 11820 21409
rect 11762 21400 11774 21403
rect 11480 21372 11774 21400
rect 11480 21360 11486 21372
rect 11762 21369 11774 21372
rect 11808 21369 11820 21403
rect 11762 21363 11820 21369
rect 8754 21292 8760 21344
rect 8812 21332 8818 21344
rect 8941 21335 8999 21341
rect 8941 21332 8953 21335
rect 8812 21304 8953 21332
rect 8812 21292 8818 21304
rect 8941 21301 8953 21304
rect 8987 21301 8999 21335
rect 12820 21332 12848 21440
rect 14645 21437 14657 21440
rect 14691 21437 14703 21471
rect 14645 21431 14703 21437
rect 15841 21471 15899 21477
rect 15841 21437 15853 21471
rect 15887 21468 15899 21471
rect 16298 21468 16304 21480
rect 15887 21440 16304 21468
rect 15887 21437 15899 21440
rect 15841 21431 15899 21437
rect 16298 21428 16304 21440
rect 16356 21428 16362 21480
rect 16393 21471 16451 21477
rect 16393 21437 16405 21471
rect 16439 21437 16451 21471
rect 16393 21431 16451 21437
rect 13814 21360 13820 21412
rect 13872 21360 13878 21412
rect 16408 21400 16436 21431
rect 18230 21428 18236 21480
rect 18288 21468 18294 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 18288 21440 20085 21468
rect 18288 21428 18294 21440
rect 20073 21437 20085 21440
rect 20119 21468 20131 21471
rect 20990 21468 20996 21480
rect 20119 21440 20996 21468
rect 20119 21437 20131 21440
rect 20073 21431 20131 21437
rect 20990 21428 20996 21440
rect 21048 21428 21054 21480
rect 21450 21428 21456 21480
rect 21508 21428 21514 21480
rect 21744 21468 21772 21499
rect 22848 21468 22876 21576
rect 23014 21564 23020 21576
rect 23072 21604 23078 21616
rect 23293 21607 23351 21613
rect 23293 21604 23305 21607
rect 23072 21576 23305 21604
rect 23072 21564 23078 21576
rect 23293 21573 23305 21576
rect 23339 21573 23351 21607
rect 23293 21567 23351 21573
rect 21744 21440 22876 21468
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21437 23535 21471
rect 23952 21468 23980 21632
rect 25424 21616 25452 21644
rect 27154 21632 27160 21644
rect 27212 21672 27218 21684
rect 27709 21675 27767 21681
rect 27709 21672 27721 21675
rect 27212 21644 27721 21672
rect 27212 21632 27218 21644
rect 27709 21641 27721 21644
rect 27755 21641 27767 21675
rect 27709 21635 27767 21641
rect 25406 21564 25412 21616
rect 25464 21564 25470 21616
rect 27338 21564 27344 21616
rect 27396 21604 27402 21616
rect 28997 21607 29055 21613
rect 28997 21604 29009 21607
rect 27396 21576 29009 21604
rect 27396 21564 27402 21576
rect 28997 21573 29009 21576
rect 29043 21573 29055 21607
rect 28997 21567 29055 21573
rect 24596 21508 25544 21536
rect 24596 21477 24624 21508
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23952 21440 24041 21468
rect 23477 21431 23535 21437
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 24581 21471 24639 21477
rect 24581 21437 24593 21471
rect 24627 21437 24639 21471
rect 24581 21431 24639 21437
rect 24673 21471 24731 21477
rect 24673 21437 24685 21471
rect 24719 21437 24731 21471
rect 24673 21431 24731 21437
rect 13924 21372 14688 21400
rect 13924 21332 13952 21372
rect 14660 21344 14688 21372
rect 15856 21372 16436 21400
rect 15856 21344 15884 21372
rect 19058 21360 19064 21412
rect 19116 21400 19122 21412
rect 19806 21403 19864 21409
rect 19806 21400 19818 21403
rect 19116 21372 19818 21400
rect 19116 21360 19122 21372
rect 19806 21369 19818 21372
rect 19852 21369 19864 21403
rect 19806 21363 19864 21369
rect 21996 21403 22054 21409
rect 21996 21369 22008 21403
rect 22042 21400 22054 21403
rect 22186 21400 22192 21412
rect 22042 21372 22192 21400
rect 22042 21369 22054 21372
rect 21996 21363 22054 21369
rect 22186 21360 22192 21372
rect 22244 21360 22250 21412
rect 23492 21400 23520 21431
rect 23845 21403 23903 21409
rect 23845 21400 23857 21403
rect 22664 21372 23857 21400
rect 22664 21344 22692 21372
rect 23845 21369 23857 21372
rect 23891 21369 23903 21403
rect 23845 21363 23903 21369
rect 24688 21344 24716 21431
rect 25222 21428 25228 21480
rect 25280 21428 25286 21480
rect 24854 21360 24860 21412
rect 24912 21360 24918 21412
rect 25516 21344 25544 21508
rect 26878 21496 26884 21548
rect 26936 21536 26942 21548
rect 29273 21539 29331 21545
rect 29273 21536 29285 21539
rect 26936 21508 29285 21536
rect 26936 21496 26942 21508
rect 29273 21505 29285 21508
rect 29319 21505 29331 21539
rect 29273 21499 29331 21505
rect 25777 21471 25835 21477
rect 25777 21437 25789 21471
rect 25823 21437 25835 21471
rect 25777 21431 25835 21437
rect 25792 21400 25820 21431
rect 25866 21428 25872 21480
rect 25924 21428 25930 21480
rect 26786 21428 26792 21480
rect 26844 21428 26850 21480
rect 28534 21428 28540 21480
rect 28592 21428 28598 21480
rect 28994 21428 29000 21480
rect 29052 21468 29058 21480
rect 29181 21471 29239 21477
rect 29181 21468 29193 21471
rect 29052 21440 29193 21468
rect 29052 21428 29058 21440
rect 29181 21437 29193 21440
rect 29227 21437 29239 21471
rect 29181 21431 29239 21437
rect 29546 21428 29552 21480
rect 29604 21428 29610 21480
rect 30006 21428 30012 21480
rect 30064 21428 30070 21480
rect 27246 21400 27252 21412
rect 25792 21372 27252 21400
rect 27246 21360 27252 21372
rect 27304 21360 27310 21412
rect 27801 21403 27859 21409
rect 27801 21369 27813 21403
rect 27847 21400 27859 21403
rect 27985 21403 28043 21409
rect 27985 21400 27997 21403
rect 27847 21372 27997 21400
rect 27847 21369 27859 21372
rect 27801 21363 27859 21369
rect 27985 21369 27997 21372
rect 28031 21400 28043 21403
rect 28074 21400 28080 21412
rect 28031 21372 28080 21400
rect 28031 21369 28043 21372
rect 27985 21363 28043 21369
rect 28074 21360 28080 21372
rect 28132 21360 28138 21412
rect 28169 21403 28227 21409
rect 28169 21369 28181 21403
rect 28215 21400 28227 21403
rect 28215 21372 29868 21400
rect 28215 21369 28227 21372
rect 28169 21363 28227 21369
rect 12820 21304 13952 21332
rect 14093 21335 14151 21341
rect 8941 21295 8999 21301
rect 14093 21301 14105 21335
rect 14139 21332 14151 21335
rect 14366 21332 14372 21344
rect 14139 21304 14372 21332
rect 14139 21301 14151 21304
rect 14093 21295 14151 21301
rect 14366 21292 14372 21304
rect 14424 21292 14430 21344
rect 14642 21292 14648 21344
rect 14700 21292 14706 21344
rect 15010 21292 15016 21344
rect 15068 21292 15074 21344
rect 15749 21335 15807 21341
rect 15749 21301 15761 21335
rect 15795 21332 15807 21335
rect 15838 21332 15844 21344
rect 15795 21304 15844 21332
rect 15795 21301 15807 21304
rect 15749 21295 15807 21301
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 18690 21292 18696 21344
rect 18748 21292 18754 21344
rect 22646 21292 22652 21344
rect 22704 21292 22710 21344
rect 22738 21292 22744 21344
rect 22796 21332 22802 21344
rect 23109 21335 23167 21341
rect 23109 21332 23121 21335
rect 22796 21304 23121 21332
rect 22796 21292 22802 21304
rect 23109 21301 23121 21304
rect 23155 21301 23167 21335
rect 23109 21295 23167 21301
rect 24578 21292 24584 21344
rect 24636 21292 24642 21344
rect 24670 21292 24676 21344
rect 24728 21292 24734 21344
rect 25498 21292 25504 21344
rect 25556 21292 25562 21344
rect 26050 21292 26056 21344
rect 26108 21292 26114 21344
rect 26142 21292 26148 21344
rect 26200 21332 26206 21344
rect 26697 21335 26755 21341
rect 26697 21332 26709 21335
rect 26200 21304 26709 21332
rect 26200 21292 26206 21304
rect 26697 21301 26709 21304
rect 26743 21301 26755 21335
rect 26697 21295 26755 21301
rect 28258 21292 28264 21344
rect 28316 21332 28322 21344
rect 28445 21335 28503 21341
rect 28445 21332 28457 21335
rect 28316 21304 28457 21332
rect 28316 21292 28322 21304
rect 28445 21301 28457 21304
rect 28491 21301 28503 21335
rect 28445 21295 28503 21301
rect 29730 21292 29736 21344
rect 29788 21292 29794 21344
rect 29840 21341 29868 21372
rect 29825 21335 29883 21341
rect 29825 21301 29837 21335
rect 29871 21301 29883 21335
rect 29825 21295 29883 21301
rect 552 21242 31808 21264
rect 552 21190 8172 21242
rect 8224 21190 8236 21242
rect 8288 21190 8300 21242
rect 8352 21190 8364 21242
rect 8416 21190 8428 21242
rect 8480 21190 15946 21242
rect 15998 21190 16010 21242
rect 16062 21190 16074 21242
rect 16126 21190 16138 21242
rect 16190 21190 16202 21242
rect 16254 21190 23720 21242
rect 23772 21190 23784 21242
rect 23836 21190 23848 21242
rect 23900 21190 23912 21242
rect 23964 21190 23976 21242
rect 24028 21190 31494 21242
rect 31546 21190 31558 21242
rect 31610 21190 31622 21242
rect 31674 21190 31686 21242
rect 31738 21190 31750 21242
rect 31802 21190 31808 21242
rect 552 21168 31808 21190
rect 10137 21131 10195 21137
rect 10137 21097 10149 21131
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 10152 21060 10180 21091
rect 11422 21088 11428 21140
rect 11480 21088 11486 21140
rect 12529 21131 12587 21137
rect 12529 21128 12541 21131
rect 12406 21100 12541 21128
rect 12406 21060 12434 21100
rect 12529 21097 12541 21100
rect 12575 21097 12587 21131
rect 12529 21091 12587 21097
rect 13354 21088 13360 21140
rect 13412 21088 13418 21140
rect 14366 21088 14372 21140
rect 14424 21128 14430 21140
rect 15746 21128 15752 21140
rect 14424 21100 15752 21128
rect 14424 21088 14430 21100
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16117 21131 16175 21137
rect 16117 21097 16129 21131
rect 16163 21097 16175 21131
rect 16117 21091 16175 21097
rect 10152 21032 12434 21060
rect 13173 21063 13231 21069
rect 13173 21029 13185 21063
rect 13219 21060 13231 21063
rect 13219 21032 14320 21060
rect 13219 21029 13231 21032
rect 13173 21023 13231 21029
rect 8846 20952 8852 21004
rect 8904 20992 8910 21004
rect 9013 20995 9071 21001
rect 9013 20992 9025 20995
rect 8904 20964 9025 20992
rect 8904 20952 8910 20964
rect 9013 20961 9025 20964
rect 9059 20961 9071 20995
rect 9013 20955 9071 20961
rect 9858 20952 9864 21004
rect 9916 20992 9922 21004
rect 10413 20995 10471 21001
rect 10413 20992 10425 20995
rect 9916 20964 10425 20992
rect 9916 20952 9922 20964
rect 10413 20961 10425 20964
rect 10459 20961 10471 20995
rect 10413 20955 10471 20961
rect 10962 20952 10968 21004
rect 11020 20952 11026 21004
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 11112 20964 11161 20992
rect 11112 20952 11118 20964
rect 11149 20961 11161 20964
rect 11195 20992 11207 20995
rect 11241 20995 11299 21001
rect 11241 20992 11253 20995
rect 11195 20964 11253 20992
rect 11195 20961 11207 20964
rect 11149 20955 11207 20961
rect 11241 20961 11253 20964
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 11882 20952 11888 21004
rect 11940 20952 11946 21004
rect 12437 20995 12495 21001
rect 12437 20961 12449 20995
rect 12483 20961 12495 20995
rect 12437 20955 12495 20961
rect 13909 20995 13967 21001
rect 13909 20961 13921 20995
rect 13955 20992 13967 20995
rect 14182 20992 14188 21004
rect 13955 20964 14188 20992
rect 13955 20961 13967 20964
rect 13909 20955 13967 20961
rect 8754 20884 8760 20936
rect 8812 20884 8818 20936
rect 12452 20856 12480 20955
rect 14182 20952 14188 20964
rect 14240 20952 14246 21004
rect 14292 21001 14320 21032
rect 14384 21001 14412 21088
rect 14820 21063 14878 21069
rect 14820 21029 14832 21063
rect 14866 21060 14878 21063
rect 16132 21060 16160 21091
rect 16666 21088 16672 21140
rect 16724 21088 16730 21140
rect 19058 21088 19064 21140
rect 19116 21088 19122 21140
rect 20993 21131 21051 21137
rect 20993 21097 21005 21131
rect 21039 21128 21051 21131
rect 21174 21128 21180 21140
rect 21039 21100 21180 21128
rect 21039 21097 21051 21100
rect 20993 21091 21051 21097
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 21450 21088 21456 21140
rect 21508 21088 21514 21140
rect 21821 21131 21879 21137
rect 21821 21097 21833 21131
rect 21867 21128 21879 21131
rect 21867 21100 22094 21128
rect 21867 21097 21879 21100
rect 21821 21091 21879 21097
rect 17954 21060 17960 21072
rect 14866 21032 16160 21060
rect 16224 21032 17960 21060
rect 14866 21029 14878 21032
rect 14820 21023 14878 21029
rect 14277 20995 14335 21001
rect 14277 20961 14289 20995
rect 14323 20961 14335 20995
rect 14277 20955 14335 20961
rect 14369 20995 14427 21001
rect 14369 20961 14381 20995
rect 14415 20961 14427 20995
rect 16224 20992 16252 21032
rect 17954 21020 17960 21032
rect 18012 21020 18018 21072
rect 20438 21060 20444 21072
rect 18892 21032 20444 21060
rect 14369 20955 14427 20961
rect 14476 20964 16252 20992
rect 12713 20927 12771 20933
rect 12713 20893 12725 20927
rect 12759 20924 12771 20927
rect 13538 20924 13544 20936
rect 12759 20896 13544 20924
rect 12759 20893 12771 20896
rect 12713 20887 12771 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 14001 20927 14059 20933
rect 14001 20893 14013 20927
rect 14047 20893 14059 20927
rect 14001 20887 14059 20893
rect 14016 20856 14044 20887
rect 14476 20856 14504 20964
rect 16298 20952 16304 21004
rect 16356 20952 16362 21004
rect 16850 20952 16856 21004
rect 16908 20992 16914 21004
rect 17782 20995 17840 21001
rect 17782 20992 17794 20995
rect 16908 20964 17794 20992
rect 16908 20952 16914 20964
rect 17782 20961 17794 20964
rect 17828 20961 17840 20995
rect 17782 20955 17840 20961
rect 18322 20952 18328 21004
rect 18380 20992 18386 21004
rect 18892 21001 18920 21032
rect 20438 21020 20444 21032
rect 20496 21020 20502 21072
rect 21468 21060 21496 21088
rect 22066 21060 22094 21100
rect 22186 21088 22192 21140
rect 22244 21088 22250 21140
rect 24578 21088 24584 21140
rect 24636 21088 24642 21140
rect 24854 21088 24860 21140
rect 24912 21088 24918 21140
rect 25222 21088 25228 21140
rect 25280 21088 25286 21140
rect 25498 21088 25504 21140
rect 25556 21128 25562 21140
rect 25556 21100 28120 21128
rect 25556 21088 25562 21100
rect 23262 21063 23320 21069
rect 23262 21060 23274 21063
rect 20548 21032 21220 21060
rect 21468 21032 21956 21060
rect 22066 21032 23274 21060
rect 18417 20995 18475 21001
rect 18417 20992 18429 20995
rect 18380 20964 18429 20992
rect 18380 20952 18386 20964
rect 18417 20961 18429 20964
rect 18463 20961 18475 20995
rect 18417 20955 18475 20961
rect 18601 20995 18659 21001
rect 18601 20961 18613 20995
rect 18647 20961 18659 20995
rect 18601 20955 18659 20961
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20961 18935 20995
rect 18877 20955 18935 20961
rect 14550 20884 14556 20936
rect 14608 20884 14614 20936
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20924 18107 20927
rect 18230 20924 18236 20936
rect 18095 20896 18236 20924
rect 18095 20893 18107 20896
rect 18049 20887 18107 20893
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 18616 20924 18644 20955
rect 19242 20952 19248 21004
rect 19300 20952 19306 21004
rect 20548 21001 20576 21032
rect 20533 20995 20591 21001
rect 20533 20992 20545 20995
rect 20364 20964 20545 20992
rect 19260 20924 19288 20952
rect 20364 20936 20392 20964
rect 20533 20961 20545 20964
rect 20579 20961 20591 20995
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 20533 20955 20591 20961
rect 20640 20964 20913 20992
rect 18616 20896 19288 20924
rect 20346 20884 20352 20936
rect 20404 20884 20410 20936
rect 20441 20927 20499 20933
rect 20441 20893 20453 20927
rect 20487 20924 20499 20927
rect 20640 20924 20668 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 21085 20995 21143 21001
rect 21085 20961 21097 20995
rect 21131 20961 21143 20995
rect 21192 20996 21220 21032
rect 21928 21001 21956 21032
rect 23262 21029 23274 21032
rect 23308 21029 23320 21063
rect 23262 21023 23320 21029
rect 24596 21060 24624 21088
rect 24596 21032 24808 21060
rect 21269 20996 21327 21001
rect 21192 20995 21327 20996
rect 21192 20968 21281 20995
rect 21085 20955 21143 20961
rect 21269 20961 21281 20968
rect 21315 20961 21327 20995
rect 21637 20995 21695 21001
rect 21637 20992 21649 20995
rect 21269 20955 21327 20961
rect 21376 20964 21649 20992
rect 20487 20896 20668 20924
rect 20487 20893 20499 20896
rect 20441 20887 20499 20893
rect 20806 20884 20812 20936
rect 20864 20884 20870 20936
rect 18417 20859 18475 20865
rect 18417 20856 18429 20859
rect 12452 20828 13952 20856
rect 14016 20828 14504 20856
rect 18064 20828 18429 20856
rect 10226 20748 10232 20800
rect 10284 20748 10290 20800
rect 10870 20748 10876 20800
rect 10928 20788 10934 20800
rect 10965 20791 11023 20797
rect 10965 20788 10977 20791
rect 10928 20760 10977 20788
rect 10928 20748 10934 20760
rect 10965 20757 10977 20760
rect 11011 20757 11023 20791
rect 10965 20751 11023 20757
rect 12802 20748 12808 20800
rect 12860 20748 12866 20800
rect 12894 20748 12900 20800
rect 12952 20748 12958 20800
rect 13924 20788 13952 20828
rect 14550 20788 14556 20800
rect 13924 20760 14556 20788
rect 14550 20748 14556 20760
rect 14608 20748 14614 20800
rect 15933 20791 15991 20797
rect 15933 20757 15945 20791
rect 15979 20788 15991 20791
rect 16574 20788 16580 20800
rect 15979 20760 16580 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16574 20748 16580 20760
rect 16632 20748 16638 20800
rect 16942 20748 16948 20800
rect 17000 20788 17006 20800
rect 18064 20788 18092 20828
rect 18417 20825 18429 20828
rect 18463 20825 18475 20859
rect 18417 20819 18475 20825
rect 20625 20859 20683 20865
rect 20625 20825 20637 20859
rect 20671 20856 20683 20859
rect 21100 20856 21128 20955
rect 21376 20924 21404 20964
rect 21637 20961 21649 20964
rect 21683 20961 21695 20995
rect 21637 20955 21695 20961
rect 21913 20995 21971 21001
rect 21913 20961 21925 20995
rect 21959 20961 21971 20995
rect 21913 20955 21971 20961
rect 22097 20995 22155 21001
rect 22097 20961 22109 20995
rect 22143 20992 22155 20995
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 22143 20964 22385 20992
rect 22143 20961 22155 20964
rect 22097 20955 22155 20961
rect 22373 20961 22385 20964
rect 22419 20961 22431 20995
rect 22373 20955 22431 20961
rect 21284 20896 21404 20924
rect 21545 20927 21603 20933
rect 21284 20865 21312 20896
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21591 20896 22017 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 22005 20893 22017 20896
rect 22051 20893 22063 20927
rect 22388 20924 22416 20955
rect 23014 20952 23020 21004
rect 23072 20952 23078 21004
rect 24596 20992 24624 21032
rect 24780 21001 24808 21032
rect 23124 20964 24624 20992
rect 24673 20995 24731 21001
rect 23124 20924 23152 20964
rect 24673 20961 24685 20995
rect 24719 20961 24731 20995
rect 24673 20955 24731 20961
rect 24765 20995 24823 21001
rect 24765 20961 24777 20995
rect 24811 20961 24823 20995
rect 24765 20955 24823 20961
rect 22388 20896 23152 20924
rect 24688 20924 24716 20955
rect 24688 20896 24808 20924
rect 22005 20887 22063 20893
rect 21269 20859 21327 20865
rect 21269 20856 21281 20859
rect 20671 20828 21281 20856
rect 20671 20825 20683 20828
rect 20625 20819 20683 20825
rect 21269 20825 21281 20828
rect 21315 20825 21327 20859
rect 21269 20819 21327 20825
rect 21361 20859 21419 20865
rect 21361 20825 21373 20859
rect 21407 20825 21419 20859
rect 24670 20856 24676 20868
rect 21361 20819 21419 20825
rect 23952 20828 24676 20856
rect 17000 20760 18092 20788
rect 17000 20748 17006 20760
rect 18138 20748 18144 20800
rect 18196 20748 18202 20800
rect 20530 20748 20536 20800
rect 20588 20788 20594 20800
rect 20717 20791 20775 20797
rect 20717 20788 20729 20791
rect 20588 20760 20729 20788
rect 20588 20748 20594 20760
rect 20717 20757 20729 20760
rect 20763 20788 20775 20791
rect 21376 20788 21404 20819
rect 20763 20760 21404 20788
rect 20763 20757 20775 20760
rect 20717 20751 20775 20757
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 23952 20788 23980 20828
rect 24670 20816 24676 20828
rect 24728 20816 24734 20868
rect 21508 20760 23980 20788
rect 21508 20748 21514 20760
rect 24394 20748 24400 20800
rect 24452 20748 24458 20800
rect 24780 20788 24808 20896
rect 24872 20856 24900 21088
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20992 25191 20995
rect 25240 20992 25268 21088
rect 25332 21032 25820 21060
rect 25332 21001 25360 21032
rect 25179 20964 25268 20992
rect 25317 20995 25375 21001
rect 25179 20961 25191 20964
rect 25133 20955 25191 20961
rect 25317 20961 25329 20995
rect 25363 20961 25375 20995
rect 25317 20955 25375 20961
rect 25406 20952 25412 21004
rect 25464 20992 25470 21004
rect 25792 21001 25820 21032
rect 25501 20995 25559 21001
rect 25501 20992 25513 20995
rect 25464 20964 25513 20992
rect 25464 20952 25470 20964
rect 25501 20961 25513 20964
rect 25547 20961 25559 20995
rect 25501 20955 25559 20961
rect 25685 20995 25743 21001
rect 25685 20961 25697 20995
rect 25731 20961 25743 20995
rect 25685 20955 25743 20961
rect 25777 20995 25835 21001
rect 25777 20961 25789 20995
rect 25823 20992 25835 20995
rect 26237 20995 26295 21001
rect 26237 20992 26249 20995
rect 25823 20964 26249 20992
rect 25823 20961 25835 20964
rect 25777 20955 25835 20961
rect 26237 20961 26249 20964
rect 26283 20961 26295 20995
rect 26237 20955 26295 20961
rect 26421 20995 26479 21001
rect 26421 20961 26433 20995
rect 26467 20992 26479 20995
rect 26620 20992 26648 21100
rect 26697 21063 26755 21069
rect 26697 21029 26709 21063
rect 26743 21060 26755 21063
rect 27617 21063 27675 21069
rect 27617 21060 27629 21063
rect 26743 21032 27629 21060
rect 26743 21029 26755 21032
rect 26697 21023 26755 21029
rect 27617 21029 27629 21032
rect 27663 21029 27675 21063
rect 27617 21023 27675 21029
rect 28092 21004 28120 21100
rect 29362 21088 29368 21140
rect 29420 21128 29426 21140
rect 29457 21131 29515 21137
rect 29457 21128 29469 21131
rect 29420 21100 29469 21128
rect 29420 21088 29426 21100
rect 29457 21097 29469 21100
rect 29503 21097 29515 21131
rect 29730 21128 29736 21140
rect 29457 21091 29515 21097
rect 29564 21100 29736 21128
rect 29564 21069 29592 21100
rect 29730 21088 29736 21100
rect 29788 21088 29794 21140
rect 29549 21063 29607 21069
rect 29549 21029 29561 21063
rect 29595 21029 29607 21063
rect 29549 21023 29607 21029
rect 26467 20964 26648 20992
rect 26467 20961 26479 20964
rect 26421 20955 26479 20961
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 25593 20927 25651 20933
rect 25593 20924 25605 20927
rect 24995 20896 25605 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 25593 20893 25605 20896
rect 25639 20893 25651 20927
rect 25593 20887 25651 20893
rect 25133 20859 25191 20865
rect 25133 20856 25145 20859
rect 24872 20828 25145 20856
rect 25133 20825 25145 20828
rect 25179 20825 25191 20859
rect 25133 20819 25191 20825
rect 25498 20816 25504 20868
rect 25556 20816 25562 20868
rect 25700 20856 25728 20955
rect 26252 20924 26280 20955
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 27157 20995 27215 21001
rect 27157 20992 27169 20995
rect 27120 20964 27169 20992
rect 27120 20952 27126 20964
rect 27157 20961 27169 20964
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 27246 20952 27252 21004
rect 27304 20952 27310 21004
rect 27522 20952 27528 21004
rect 27580 20952 27586 21004
rect 27709 20995 27767 21001
rect 27709 20961 27721 20995
rect 27755 20992 27767 20995
rect 27982 20992 27988 21004
rect 27755 20964 27988 20992
rect 27755 20961 27767 20964
rect 27709 20955 27767 20961
rect 27982 20952 27988 20964
rect 28040 20952 28046 21004
rect 28074 20952 28080 21004
rect 28132 20952 28138 21004
rect 29017 20995 29075 21001
rect 29017 20961 29029 20995
rect 29063 20992 29075 20995
rect 29917 20995 29975 21001
rect 29063 20964 29776 20992
rect 29063 20961 29075 20964
rect 29017 20955 29075 20961
rect 26789 20927 26847 20933
rect 26252 20896 26556 20924
rect 26418 20856 26424 20868
rect 25700 20828 26424 20856
rect 26418 20816 26424 20828
rect 26476 20816 26482 20868
rect 26528 20865 26556 20896
rect 26789 20893 26801 20927
rect 26835 20924 26847 20927
rect 27430 20924 27436 20936
rect 26835 20896 27436 20924
rect 26835 20893 26847 20896
rect 26789 20887 26847 20893
rect 27430 20884 27436 20896
rect 27488 20884 27494 20936
rect 29270 20884 29276 20936
rect 29328 20884 29334 20936
rect 26513 20859 26571 20865
rect 26513 20825 26525 20859
rect 26559 20825 26571 20859
rect 26513 20819 26571 20825
rect 25516 20788 25544 20816
rect 24780 20760 25544 20788
rect 25958 20748 25964 20800
rect 26016 20788 26022 20800
rect 26053 20791 26111 20797
rect 26053 20788 26065 20791
rect 26016 20760 26065 20788
rect 26016 20748 26022 20760
rect 26053 20757 26065 20760
rect 26099 20757 26111 20791
rect 26528 20788 26556 20819
rect 26602 20816 26608 20868
rect 26660 20856 26666 20868
rect 29748 20865 29776 20964
rect 29917 20961 29929 20995
rect 29963 20992 29975 20995
rect 30006 20992 30012 21004
rect 29963 20964 30012 20992
rect 29963 20961 29975 20964
rect 29917 20955 29975 20961
rect 30006 20952 30012 20964
rect 30064 20952 30070 21004
rect 26973 20859 27031 20865
rect 26973 20856 26985 20859
rect 26660 20828 26985 20856
rect 26660 20816 26666 20828
rect 26973 20825 26985 20828
rect 27019 20825 27031 20859
rect 26973 20819 27031 20825
rect 27065 20859 27123 20865
rect 27065 20825 27077 20859
rect 27111 20856 27123 20859
rect 27157 20859 27215 20865
rect 27157 20856 27169 20859
rect 27111 20828 27169 20856
rect 27111 20825 27123 20828
rect 27065 20819 27123 20825
rect 27157 20825 27169 20828
rect 27203 20825 27215 20859
rect 27157 20819 27215 20825
rect 29733 20859 29791 20865
rect 29733 20825 29745 20859
rect 29779 20825 29791 20859
rect 29733 20819 29791 20825
rect 27080 20788 27108 20819
rect 26528 20760 27108 20788
rect 26053 20751 26111 20757
rect 27246 20748 27252 20800
rect 27304 20788 27310 20800
rect 27893 20791 27951 20797
rect 27893 20788 27905 20791
rect 27304 20760 27905 20788
rect 27304 20748 27310 20760
rect 27893 20757 27905 20760
rect 27939 20757 27951 20791
rect 27893 20751 27951 20757
rect 552 20698 31648 20720
rect 552 20646 4285 20698
rect 4337 20646 4349 20698
rect 4401 20646 4413 20698
rect 4465 20646 4477 20698
rect 4529 20646 4541 20698
rect 4593 20646 12059 20698
rect 12111 20646 12123 20698
rect 12175 20646 12187 20698
rect 12239 20646 12251 20698
rect 12303 20646 12315 20698
rect 12367 20646 19833 20698
rect 19885 20646 19897 20698
rect 19949 20646 19961 20698
rect 20013 20646 20025 20698
rect 20077 20646 20089 20698
rect 20141 20646 27607 20698
rect 27659 20646 27671 20698
rect 27723 20646 27735 20698
rect 27787 20646 27799 20698
rect 27851 20646 27863 20698
rect 27915 20646 31648 20698
rect 552 20624 31648 20646
rect 8846 20544 8852 20596
rect 8904 20544 8910 20596
rect 11514 20584 11520 20596
rect 9968 20556 11520 20584
rect 8754 20448 8760 20460
rect 7760 20420 8760 20448
rect 4893 20383 4951 20389
rect 4893 20349 4905 20383
rect 4939 20380 4951 20383
rect 5074 20380 5080 20392
rect 4939 20352 5080 20380
rect 4939 20349 4951 20352
rect 4893 20343 4951 20349
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 5997 20383 6055 20389
rect 5997 20380 6009 20383
rect 5460 20352 6009 20380
rect 5460 20256 5488 20352
rect 5997 20349 6009 20352
rect 6043 20349 6055 20383
rect 5997 20343 6055 20349
rect 6733 20383 6791 20389
rect 6733 20349 6745 20383
rect 6779 20380 6791 20383
rect 7760 20380 7788 20420
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 9968 20457 9996 20556
rect 11514 20544 11520 20556
rect 11572 20544 11578 20596
rect 12802 20544 12808 20596
rect 12860 20544 12866 20596
rect 15470 20584 15476 20596
rect 13648 20556 15476 20584
rect 11333 20519 11391 20525
rect 11333 20485 11345 20519
rect 11379 20516 11391 20519
rect 11379 20488 12434 20516
rect 11379 20485 11391 20488
rect 11333 20479 11391 20485
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20417 10011 20451
rect 12406 20448 12434 20488
rect 13538 20476 13544 20528
rect 13596 20476 13602 20528
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 12406 20420 13185 20448
rect 9953 20411 10011 20417
rect 13173 20417 13185 20420
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 13648 20392 13676 20556
rect 15470 20544 15476 20556
rect 15528 20544 15534 20596
rect 15657 20587 15715 20593
rect 15657 20553 15669 20587
rect 15703 20584 15715 20587
rect 15703 20556 17908 20584
rect 15703 20553 15715 20556
rect 15657 20547 15715 20553
rect 13906 20516 13912 20528
rect 13832 20488 13912 20516
rect 13832 20448 13860 20488
rect 13906 20476 13912 20488
rect 13964 20516 13970 20528
rect 15672 20516 15700 20547
rect 13964 20488 15700 20516
rect 17037 20519 17095 20525
rect 13964 20476 13970 20488
rect 17037 20485 17049 20519
rect 17083 20516 17095 20519
rect 17083 20488 17816 20516
rect 17083 20485 17095 20488
rect 17037 20479 17095 20485
rect 13740 20420 13860 20448
rect 6779 20352 7788 20380
rect 8665 20383 8723 20389
rect 6779 20349 6791 20352
rect 6733 20343 6791 20349
rect 7208 20324 7236 20352
rect 8665 20349 8677 20383
rect 8711 20380 8723 20383
rect 8846 20380 8852 20392
rect 8711 20352 8852 20380
rect 8711 20349 8723 20352
rect 8665 20343 8723 20349
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20380 9275 20383
rect 9398 20380 9404 20392
rect 9263 20352 9404 20380
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20380 9643 20383
rect 9677 20383 9735 20389
rect 9677 20380 9689 20383
rect 9631 20352 9689 20380
rect 9631 20349 9643 20352
rect 9585 20343 9643 20349
rect 9677 20349 9689 20352
rect 9723 20349 9735 20383
rect 9677 20343 9735 20349
rect 9858 20340 9864 20392
rect 9916 20340 9922 20392
rect 10226 20389 10232 20392
rect 10220 20380 10232 20389
rect 10187 20352 10232 20380
rect 10220 20343 10232 20352
rect 10226 20340 10232 20343
rect 10284 20340 10290 20392
rect 11422 20340 11428 20392
rect 11480 20340 11486 20392
rect 11698 20340 11704 20392
rect 11756 20340 11762 20392
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13630 20380 13636 20392
rect 13035 20352 13636 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 13740 20389 13768 20420
rect 14090 20408 14096 20460
rect 14148 20408 14154 20460
rect 14550 20408 14556 20460
rect 14608 20408 14614 20460
rect 15746 20408 15752 20460
rect 15804 20448 15810 20460
rect 16393 20451 16451 20457
rect 16393 20448 16405 20451
rect 15804 20420 16405 20448
rect 15804 20408 15810 20420
rect 16393 20417 16405 20420
rect 16439 20417 16451 20451
rect 16393 20411 16451 20417
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 13725 20383 13783 20389
rect 13725 20349 13737 20383
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20380 14795 20383
rect 15010 20380 15016 20392
rect 14783 20352 15016 20380
rect 14783 20349 14795 20352
rect 14737 20343 14795 20349
rect 6454 20272 6460 20324
rect 6512 20312 6518 20324
rect 6978 20315 7036 20321
rect 6978 20312 6990 20315
rect 6512 20284 6990 20312
rect 6512 20272 6518 20284
rect 6978 20281 6990 20284
rect 7024 20281 7036 20315
rect 6978 20275 7036 20281
rect 7190 20272 7196 20324
rect 7248 20272 7254 20324
rect 13832 20312 13860 20343
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 15102 20340 15108 20392
rect 15160 20340 15166 20392
rect 15286 20340 15292 20392
rect 15344 20340 15350 20392
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 16669 20383 16727 20389
rect 16669 20380 16681 20383
rect 16632 20352 16681 20380
rect 16632 20340 16638 20352
rect 16669 20349 16681 20352
rect 16715 20349 16727 20383
rect 16669 20343 16727 20349
rect 17310 20340 17316 20392
rect 17368 20380 17374 20392
rect 17788 20389 17816 20488
rect 17880 20448 17908 20556
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18877 20587 18935 20593
rect 18877 20584 18889 20587
rect 18012 20556 18889 20584
rect 18012 20544 18018 20556
rect 18877 20553 18889 20556
rect 18923 20553 18935 20587
rect 18877 20547 18935 20553
rect 18966 20544 18972 20596
rect 19024 20584 19030 20596
rect 20622 20584 20628 20596
rect 19024 20556 20628 20584
rect 19024 20544 19030 20556
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 20901 20587 20959 20593
rect 20901 20584 20913 20587
rect 20864 20556 20913 20584
rect 20864 20544 20870 20556
rect 20901 20553 20913 20556
rect 20947 20553 20959 20587
rect 20901 20547 20959 20553
rect 24949 20587 25007 20593
rect 24949 20553 24961 20587
rect 24995 20584 25007 20587
rect 25041 20587 25099 20593
rect 25041 20584 25053 20587
rect 24995 20556 25053 20584
rect 24995 20553 25007 20556
rect 24949 20547 25007 20553
rect 25041 20553 25053 20556
rect 25087 20553 25099 20587
rect 25041 20547 25099 20553
rect 27433 20587 27491 20593
rect 27433 20553 27445 20587
rect 27479 20584 27491 20587
rect 27522 20584 27528 20596
rect 27479 20556 27528 20584
rect 27479 20553 27491 20556
rect 27433 20547 27491 20553
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 30006 20584 30012 20596
rect 28460 20556 30012 20584
rect 21729 20519 21787 20525
rect 21729 20516 21741 20519
rect 18432 20488 21741 20516
rect 17954 20448 17960 20460
rect 17880 20420 17960 20448
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 17589 20383 17647 20389
rect 17589 20380 17601 20383
rect 17368 20352 17601 20380
rect 17368 20340 17374 20352
rect 17589 20349 17601 20352
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 17773 20383 17831 20389
rect 17773 20349 17785 20383
rect 17819 20349 17831 20383
rect 17773 20343 17831 20349
rect 18046 20340 18052 20392
rect 18104 20389 18110 20392
rect 18104 20383 18138 20389
rect 18126 20349 18138 20383
rect 18104 20343 18138 20349
rect 18325 20383 18383 20389
rect 18325 20349 18337 20383
rect 18371 20376 18383 20383
rect 18432 20376 18460 20488
rect 21729 20485 21741 20488
rect 21775 20485 21787 20519
rect 21729 20479 21787 20485
rect 22465 20519 22523 20525
rect 22465 20485 22477 20519
rect 22511 20485 22523 20519
rect 22465 20479 22523 20485
rect 21450 20448 21456 20460
rect 20272 20420 20570 20448
rect 19058 20389 19064 20392
rect 19056 20380 19064 20389
rect 18371 20349 18460 20376
rect 19019 20352 19064 20380
rect 18325 20348 18460 20349
rect 18325 20343 18383 20348
rect 19056 20343 19064 20352
rect 18104 20340 18110 20343
rect 19058 20340 19064 20343
rect 19116 20340 19122 20392
rect 19334 20340 19340 20392
rect 19392 20389 19398 20392
rect 19392 20383 19431 20389
rect 19419 20349 19431 20383
rect 19392 20343 19431 20349
rect 19392 20340 19398 20343
rect 19518 20340 19524 20392
rect 19576 20340 19582 20392
rect 20162 20380 20168 20392
rect 19812 20352 20168 20380
rect 8128 20284 13860 20312
rect 15749 20315 15807 20321
rect 5077 20247 5135 20253
rect 5077 20213 5089 20247
rect 5123 20244 5135 20247
rect 5166 20244 5172 20256
rect 5123 20216 5172 20244
rect 5123 20213 5135 20216
rect 5077 20207 5135 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 5442 20204 5448 20256
rect 5500 20204 5506 20256
rect 6178 20204 6184 20256
rect 6236 20204 6242 20256
rect 8128 20253 8156 20284
rect 15749 20281 15761 20315
rect 15795 20312 15807 20315
rect 18966 20312 18972 20324
rect 15795 20284 18972 20312
rect 15795 20281 15807 20284
rect 15749 20275 15807 20281
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20213 8171 20247
rect 8113 20207 8171 20213
rect 9030 20204 9036 20256
rect 9088 20204 9094 20256
rect 9766 20204 9772 20256
rect 9824 20204 9830 20256
rect 11606 20204 11612 20256
rect 11664 20204 11670 20256
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 15764 20244 15792 20275
rect 18966 20272 18972 20284
rect 19024 20272 19030 20324
rect 19153 20315 19211 20321
rect 19153 20281 19165 20315
rect 19199 20281 19211 20315
rect 19153 20275 19211 20281
rect 19245 20315 19303 20321
rect 19245 20281 19257 20315
rect 19291 20312 19303 20315
rect 19812 20312 19840 20352
rect 20162 20340 20168 20352
rect 20220 20340 20226 20392
rect 20272 20389 20300 20420
rect 20542 20392 20570 20420
rect 20732 20420 21456 20448
rect 20732 20392 20760 20420
rect 21450 20408 21456 20420
rect 21508 20408 21514 20460
rect 22480 20448 22508 20479
rect 24486 20476 24492 20528
rect 24544 20476 24550 20528
rect 24670 20476 24676 20528
rect 24728 20516 24734 20528
rect 28460 20525 28488 20556
rect 30006 20544 30012 20556
rect 30064 20544 30070 20596
rect 28445 20519 28503 20525
rect 28445 20516 28457 20519
rect 24728 20488 24808 20516
rect 24728 20476 24734 20488
rect 24780 20457 24808 20488
rect 25424 20488 26556 20516
rect 25424 20457 25452 20488
rect 22204 20420 22508 20448
rect 24765 20451 24823 20457
rect 20530 20389 20536 20392
rect 20257 20383 20315 20389
rect 20257 20349 20269 20383
rect 20303 20349 20315 20383
rect 20257 20343 20315 20349
rect 20349 20383 20407 20389
rect 20349 20349 20361 20383
rect 20395 20349 20407 20383
rect 20349 20343 20407 20349
rect 20527 20343 20536 20389
rect 20588 20380 20594 20392
rect 20588 20352 20627 20380
rect 20364 20312 20392 20343
rect 20530 20340 20536 20343
rect 20588 20340 20594 20352
rect 20714 20340 20720 20392
rect 20772 20340 20778 20392
rect 20901 20383 20959 20389
rect 20901 20349 20913 20383
rect 20947 20349 20959 20383
rect 20901 20343 20959 20349
rect 20916 20312 20944 20343
rect 21082 20340 21088 20392
rect 21140 20380 21146 20392
rect 21818 20380 21824 20392
rect 21140 20352 21824 20380
rect 21140 20340 21146 20352
rect 21818 20340 21824 20352
rect 21876 20380 21882 20392
rect 22204 20389 22232 20420
rect 24765 20417 24777 20451
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 25409 20451 25467 20457
rect 25409 20417 25421 20451
rect 25455 20417 25467 20451
rect 25409 20411 25467 20417
rect 21913 20383 21971 20389
rect 21913 20380 21925 20383
rect 21876 20352 21925 20380
rect 21876 20340 21882 20352
rect 21913 20349 21925 20352
rect 21959 20349 21971 20383
rect 21913 20343 21971 20349
rect 22189 20383 22247 20389
rect 22189 20349 22201 20383
rect 22235 20349 22247 20383
rect 22189 20343 22247 20349
rect 22370 20340 22376 20392
rect 22428 20340 22434 20392
rect 22462 20340 22468 20392
rect 22520 20380 22526 20392
rect 22603 20383 22661 20389
rect 22603 20380 22615 20383
rect 22520 20352 22615 20380
rect 22520 20340 22526 20352
rect 22603 20349 22615 20352
rect 22649 20349 22661 20383
rect 22603 20343 22661 20349
rect 22738 20340 22744 20392
rect 22796 20340 22802 20392
rect 22922 20340 22928 20392
rect 22980 20389 22986 20392
rect 22980 20383 23019 20389
rect 23007 20349 23019 20383
rect 22980 20343 23019 20349
rect 22980 20340 22986 20343
rect 23106 20340 23112 20392
rect 23164 20380 23170 20392
rect 24673 20383 24731 20389
rect 24673 20380 24685 20383
rect 23164 20352 24685 20380
rect 23164 20340 23170 20352
rect 24673 20349 24685 20352
rect 24719 20380 24731 20383
rect 24854 20380 24860 20392
rect 24719 20352 24860 20380
rect 24719 20349 24731 20352
rect 24673 20343 24731 20349
rect 24854 20340 24860 20352
rect 24912 20340 24918 20392
rect 26418 20389 26424 20392
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 25148 20352 25237 20380
rect 19291 20284 19840 20312
rect 20272 20284 20944 20312
rect 19291 20281 19303 20284
rect 19245 20275 19303 20281
rect 13504 20216 15792 20244
rect 16577 20247 16635 20253
rect 13504 20204 13510 20216
rect 16577 20213 16589 20247
rect 16623 20244 16635 20247
rect 18690 20244 18696 20256
rect 16623 20216 18696 20244
rect 16623 20213 16635 20216
rect 16577 20207 16635 20213
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 19168 20244 19196 20275
rect 20272 20256 20300 20284
rect 22830 20272 22836 20324
rect 22888 20312 22894 20324
rect 23382 20312 23388 20324
rect 22888 20284 23388 20312
rect 22888 20272 22894 20284
rect 23382 20272 23388 20284
rect 23440 20272 23446 20324
rect 24578 20272 24584 20324
rect 24636 20312 24642 20324
rect 24949 20315 25007 20321
rect 24949 20312 24961 20315
rect 24636 20284 24961 20312
rect 24636 20272 24642 20284
rect 24949 20281 24961 20284
rect 24995 20281 25007 20315
rect 24949 20275 25007 20281
rect 19978 20244 19984 20256
rect 19168 20216 19984 20244
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 20070 20204 20076 20256
rect 20128 20204 20134 20256
rect 20254 20204 20260 20256
rect 20312 20204 20318 20256
rect 20438 20204 20444 20256
rect 20496 20204 20502 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 24762 20244 24768 20256
rect 20680 20216 24768 20244
rect 20680 20204 20686 20216
rect 24762 20204 24768 20216
rect 24820 20244 24826 20256
rect 25148 20244 25176 20352
rect 25225 20349 25237 20352
rect 25271 20349 25283 20383
rect 26412 20380 26424 20389
rect 26379 20352 26424 20380
rect 25225 20343 25283 20349
rect 26412 20343 26424 20352
rect 26418 20340 26424 20343
rect 26476 20340 26482 20392
rect 26528 20312 26556 20488
rect 26712 20488 27844 20516
rect 26712 20389 26740 20488
rect 26789 20451 26847 20457
rect 26789 20417 26801 20451
rect 26835 20448 26847 20451
rect 27430 20448 27436 20460
rect 26835 20420 27436 20448
rect 26835 20417 26847 20420
rect 26789 20411 26847 20417
rect 27430 20408 27436 20420
rect 27488 20448 27494 20460
rect 27709 20451 27767 20457
rect 27709 20448 27721 20451
rect 27488 20420 27721 20448
rect 27488 20408 27494 20420
rect 27709 20417 27721 20420
rect 27755 20417 27767 20451
rect 27709 20411 27767 20417
rect 27816 20448 27844 20488
rect 28184 20488 28457 20516
rect 28184 20457 28212 20488
rect 28445 20485 28457 20488
rect 28491 20485 28503 20519
rect 28445 20479 28503 20485
rect 28997 20519 29055 20525
rect 28997 20485 29009 20519
rect 29043 20485 29055 20519
rect 28997 20479 29055 20485
rect 28169 20451 28227 20457
rect 28169 20448 28181 20451
rect 27816 20420 28181 20448
rect 26697 20383 26755 20389
rect 26697 20349 26709 20383
rect 26743 20349 26755 20383
rect 26697 20343 26755 20349
rect 26878 20340 26884 20392
rect 26936 20340 26942 20392
rect 26973 20383 27031 20389
rect 26973 20349 26985 20383
rect 27019 20380 27031 20383
rect 27019 20352 27568 20380
rect 27019 20349 27031 20352
rect 26973 20343 27031 20349
rect 27246 20312 27252 20324
rect 26528 20284 27252 20312
rect 27246 20272 27252 20284
rect 27304 20272 27310 20324
rect 24820 20216 25176 20244
rect 24820 20204 24826 20216
rect 26234 20204 26240 20256
rect 26292 20204 26298 20256
rect 27154 20204 27160 20256
rect 27212 20204 27218 20256
rect 27540 20244 27568 20352
rect 27614 20340 27620 20392
rect 27672 20340 27678 20392
rect 27816 20389 27844 20420
rect 28169 20417 28181 20420
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 28626 20408 28632 20460
rect 28684 20448 28690 20460
rect 29012 20448 29040 20479
rect 28684 20420 29040 20448
rect 28684 20408 28690 20420
rect 27801 20383 27859 20389
rect 27801 20349 27813 20383
rect 27847 20349 27859 20383
rect 27801 20343 27859 20349
rect 28074 20340 28080 20392
rect 28132 20380 28138 20392
rect 28445 20383 28503 20389
rect 28445 20380 28457 20383
rect 28132 20352 28457 20380
rect 28132 20340 28138 20352
rect 28445 20349 28457 20352
rect 28491 20349 28503 20383
rect 28445 20343 28503 20349
rect 28537 20383 28595 20389
rect 28537 20349 28549 20383
rect 28583 20349 28595 20383
rect 28537 20343 28595 20349
rect 28350 20272 28356 20324
rect 28408 20272 28414 20324
rect 27982 20244 27988 20256
rect 27540 20216 27988 20244
rect 27982 20204 27988 20216
rect 28040 20244 28046 20256
rect 28077 20247 28135 20253
rect 28077 20244 28089 20247
rect 28040 20216 28089 20244
rect 28040 20204 28046 20216
rect 28077 20213 28089 20216
rect 28123 20244 28135 20247
rect 28552 20244 28580 20343
rect 29270 20340 29276 20392
rect 29328 20380 29334 20392
rect 30377 20383 30435 20389
rect 30377 20380 30389 20383
rect 29328 20352 30389 20380
rect 29328 20340 29334 20352
rect 30377 20349 30389 20352
rect 30423 20349 30435 20383
rect 30377 20343 30435 20349
rect 28721 20315 28779 20321
rect 28721 20281 28733 20315
rect 28767 20312 28779 20315
rect 28810 20312 28816 20324
rect 28767 20284 28816 20312
rect 28767 20281 28779 20284
rect 28721 20275 28779 20281
rect 28810 20272 28816 20284
rect 28868 20272 28874 20324
rect 29914 20272 29920 20324
rect 29972 20312 29978 20324
rect 30110 20315 30168 20321
rect 30110 20312 30122 20315
rect 29972 20284 30122 20312
rect 29972 20272 29978 20284
rect 30110 20281 30122 20284
rect 30156 20281 30168 20315
rect 30110 20275 30168 20281
rect 28123 20216 28580 20244
rect 28123 20213 28135 20216
rect 28077 20207 28135 20213
rect 552 20154 31808 20176
rect 552 20102 8172 20154
rect 8224 20102 8236 20154
rect 8288 20102 8300 20154
rect 8352 20102 8364 20154
rect 8416 20102 8428 20154
rect 8480 20102 15946 20154
rect 15998 20102 16010 20154
rect 16062 20102 16074 20154
rect 16126 20102 16138 20154
rect 16190 20102 16202 20154
rect 16254 20102 23720 20154
rect 23772 20102 23784 20154
rect 23836 20102 23848 20154
rect 23900 20102 23912 20154
rect 23964 20102 23976 20154
rect 24028 20102 31494 20154
rect 31546 20102 31558 20154
rect 31610 20102 31622 20154
rect 31674 20102 31686 20154
rect 31738 20102 31750 20154
rect 31802 20102 31808 20154
rect 552 20080 31808 20102
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20009 3479 20043
rect 3421 20003 3479 20009
rect 2958 19864 2964 19916
rect 3016 19864 3022 19916
rect 3237 19907 3295 19913
rect 3237 19873 3249 19907
rect 3283 19904 3295 19907
rect 3326 19904 3332 19916
rect 3283 19876 3332 19904
rect 3283 19873 3295 19876
rect 3237 19867 3295 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 3436 19904 3464 20003
rect 6178 20000 6184 20052
rect 6236 20000 6242 20052
rect 6454 20000 6460 20052
rect 6512 20000 6518 20052
rect 7929 20043 7987 20049
rect 7929 20009 7941 20043
rect 7975 20009 7987 20043
rect 7929 20003 7987 20009
rect 5902 19972 5908 19984
rect 5000 19944 5908 19972
rect 5000 19913 5028 19944
rect 5902 19932 5908 19944
rect 5960 19932 5966 19984
rect 6196 19972 6224 20000
rect 6794 19975 6852 19981
rect 6794 19972 6806 19975
rect 6196 19944 6806 19972
rect 6794 19941 6806 19944
rect 6840 19941 6852 19975
rect 7944 19972 7972 20003
rect 9766 20000 9772 20052
rect 9824 20000 9830 20052
rect 9861 20043 9919 20049
rect 9861 20009 9873 20043
rect 9907 20040 9919 20043
rect 10042 20040 10048 20052
rect 9907 20012 10048 20040
rect 9907 20009 9919 20012
rect 9861 20003 9919 20009
rect 10042 20000 10048 20012
rect 10100 20040 10106 20052
rect 10594 20040 10600 20052
rect 10100 20012 10600 20040
rect 10100 20000 10106 20012
rect 10594 20000 10600 20012
rect 10652 20040 10658 20052
rect 11241 20043 11299 20049
rect 10652 20012 11100 20040
rect 10652 20000 10658 20012
rect 9214 19972 9220 19984
rect 7944 19944 9220 19972
rect 6794 19935 6852 19941
rect 9214 19932 9220 19944
rect 9272 19932 9278 19984
rect 9585 19975 9643 19981
rect 9585 19941 9597 19975
rect 9631 19972 9643 19975
rect 9784 19972 9812 20000
rect 9631 19944 9812 19972
rect 9631 19941 9643 19944
rect 9585 19935 9643 19941
rect 9950 19932 9956 19984
rect 10008 19972 10014 19984
rect 10229 19975 10287 19981
rect 10229 19972 10241 19975
rect 10008 19944 10241 19972
rect 10008 19932 10014 19944
rect 10229 19941 10241 19944
rect 10275 19972 10287 19975
rect 10962 19972 10968 19984
rect 10275 19944 10968 19972
rect 10275 19941 10287 19944
rect 10229 19935 10287 19941
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 3697 19907 3755 19913
rect 3697 19904 3709 19907
rect 3436 19876 3709 19904
rect 3697 19873 3709 19876
rect 3743 19873 3755 19907
rect 3697 19867 3755 19873
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19873 4859 19907
rect 4801 19867 4859 19873
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19873 5043 19907
rect 4985 19867 5043 19873
rect 3881 19771 3939 19777
rect 3881 19737 3893 19771
rect 3927 19768 3939 19771
rect 4706 19768 4712 19780
rect 3927 19740 4712 19768
rect 3927 19737 3939 19740
rect 3881 19731 3939 19737
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 4816 19768 4844 19867
rect 5074 19864 5080 19916
rect 5132 19864 5138 19916
rect 5350 19864 5356 19916
rect 5408 19864 5414 19916
rect 6273 19907 6331 19913
rect 6273 19873 6285 19907
rect 6319 19904 6331 19907
rect 6362 19904 6368 19916
rect 6319 19876 6368 19904
rect 6319 19873 6331 19876
rect 6273 19867 6331 19873
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 6549 19907 6607 19913
rect 6549 19873 6561 19907
rect 6595 19904 6607 19907
rect 6638 19904 6644 19916
rect 6595 19876 6644 19904
rect 6595 19873 6607 19876
rect 6549 19867 6607 19873
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 8846 19864 8852 19916
rect 8904 19864 8910 19916
rect 8941 19907 8999 19913
rect 8941 19873 8953 19907
rect 8987 19904 8999 19907
rect 9030 19904 9036 19916
rect 8987 19876 9036 19904
rect 8987 19873 8999 19876
rect 8941 19867 8999 19873
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 9456 19876 9873 19904
rect 9456 19864 9462 19876
rect 5092 19836 5120 19864
rect 5092 19808 5396 19836
rect 5368 19777 5396 19808
rect 5626 19796 5632 19848
rect 5684 19796 5690 19848
rect 8662 19796 8668 19848
rect 8720 19796 8726 19848
rect 5353 19771 5411 19777
rect 4816 19740 5304 19768
rect 5276 19712 5304 19740
rect 5353 19737 5365 19771
rect 5399 19737 5411 19771
rect 5353 19731 5411 19737
rect 5442 19728 5448 19780
rect 5500 19728 5506 19780
rect 8864 19768 8892 19864
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 9692 19780 9720 19876
rect 9861 19873 9873 19876
rect 9907 19873 9919 19907
rect 9861 19867 9919 19873
rect 10045 19907 10103 19913
rect 10045 19873 10057 19907
rect 10091 19904 10103 19907
rect 10410 19904 10416 19916
rect 10091 19876 10416 19904
rect 10091 19873 10103 19876
rect 10045 19867 10103 19873
rect 10410 19864 10416 19876
rect 10468 19864 10474 19916
rect 11072 19913 11100 20012
rect 11241 20009 11253 20043
rect 11287 20009 11299 20043
rect 11241 20003 11299 20009
rect 13817 20043 13875 20049
rect 13817 20009 13829 20043
rect 13863 20009 13875 20043
rect 13817 20003 13875 20009
rect 14277 20043 14335 20049
rect 14277 20009 14289 20043
rect 14323 20040 14335 20043
rect 15102 20040 15108 20052
rect 14323 20012 15108 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 11256 19972 11284 20003
rect 11578 19975 11636 19981
rect 11578 19972 11590 19975
rect 11256 19944 11590 19972
rect 11578 19941 11590 19944
rect 11624 19941 11636 19975
rect 11578 19935 11636 19941
rect 13538 19932 13544 19984
rect 13596 19932 13602 19984
rect 11057 19907 11115 19913
rect 11057 19873 11069 19907
rect 11103 19873 11115 19907
rect 11057 19867 11115 19873
rect 13170 19864 13176 19916
rect 13228 19864 13234 19916
rect 13262 19864 13268 19916
rect 13320 19864 13326 19916
rect 13446 19864 13452 19916
rect 13504 19864 13510 19916
rect 13722 19913 13728 19916
rect 13679 19907 13728 19913
rect 13679 19873 13691 19907
rect 13725 19873 13728 19907
rect 13679 19867 13728 19873
rect 13722 19864 13728 19867
rect 13780 19864 13786 19916
rect 13832 19904 13860 20003
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15470 20000 15476 20052
rect 15528 20040 15534 20052
rect 16209 20043 16267 20049
rect 16209 20040 16221 20043
rect 15528 20012 16221 20040
rect 15528 20000 15534 20012
rect 16209 20009 16221 20012
rect 16255 20040 16267 20043
rect 16666 20040 16672 20052
rect 16255 20012 16672 20040
rect 16255 20009 16267 20012
rect 16209 20003 16267 20009
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 16850 20000 16856 20052
rect 16908 20000 16914 20052
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 18230 20040 18236 20052
rect 17552 20012 18236 20040
rect 17552 20000 17558 20012
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 19061 20043 19119 20049
rect 19061 20009 19073 20043
rect 19107 20040 19119 20043
rect 19334 20040 19340 20052
rect 19107 20012 19340 20040
rect 19107 20009 19119 20012
rect 19061 20003 19119 20009
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 20438 20000 20444 20052
rect 20496 20000 20502 20052
rect 22649 20043 22707 20049
rect 22649 20009 22661 20043
rect 22695 20040 22707 20043
rect 22922 20040 22928 20052
rect 22695 20012 22928 20040
rect 22695 20009 22707 20012
rect 22649 20003 22707 20009
rect 22922 20000 22928 20012
rect 22980 20000 22986 20052
rect 24394 20000 24400 20052
rect 24452 20000 24458 20052
rect 24762 20040 24768 20052
rect 24596 20012 24768 20040
rect 16942 19932 16948 19984
rect 17000 19932 17006 19984
rect 17678 19972 17684 19984
rect 17328 19944 17684 19972
rect 13897 19907 13955 19913
rect 13897 19904 13909 19907
rect 13832 19876 13909 19904
rect 13897 19873 13909 19876
rect 13943 19873 13955 19907
rect 13897 19867 13955 19873
rect 14820 19907 14878 19913
rect 14820 19873 14832 19907
rect 14866 19904 14878 19907
rect 15102 19904 15108 19916
rect 14866 19876 15108 19904
rect 14866 19873 14878 19876
rect 14820 19867 14878 19873
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 16482 19864 16488 19916
rect 16540 19864 16546 19916
rect 17328 19913 17356 19944
rect 17678 19932 17684 19944
rect 17736 19932 17742 19984
rect 17948 19975 18006 19981
rect 17948 19941 17960 19975
rect 17994 19972 18006 19975
rect 20349 19975 20407 19981
rect 17994 19944 19472 19972
rect 17994 19941 18006 19944
rect 17948 19935 18006 19941
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 17313 19907 17371 19913
rect 17313 19904 17325 19907
rect 17267 19876 17325 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 17313 19873 17325 19876
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 17405 19907 17463 19913
rect 17405 19873 17417 19907
rect 17451 19904 17463 19907
rect 19150 19904 19156 19916
rect 17451 19876 19156 19904
rect 17451 19873 17463 19876
rect 17405 19867 17463 19873
rect 11333 19839 11391 19845
rect 11333 19805 11345 19839
rect 11379 19805 11391 19839
rect 11333 19799 11391 19805
rect 9033 19771 9091 19777
rect 9033 19768 9045 19771
rect 8864 19740 9045 19768
rect 9033 19737 9045 19740
rect 9079 19737 9091 19771
rect 9033 19731 9091 19737
rect 9125 19771 9183 19777
rect 9125 19737 9137 19771
rect 9171 19737 9183 19771
rect 9125 19731 9183 19737
rect 3145 19703 3203 19709
rect 3145 19669 3157 19703
rect 3191 19700 3203 19703
rect 3694 19700 3700 19712
rect 3191 19672 3700 19700
rect 3191 19669 3203 19672
rect 3145 19663 3203 19669
rect 3694 19660 3700 19672
rect 3752 19660 3758 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 4525 19703 4583 19709
rect 4525 19700 4537 19703
rect 4212 19672 4537 19700
rect 4212 19660 4218 19672
rect 4525 19669 4537 19672
rect 4571 19669 4583 19703
rect 4525 19663 4583 19669
rect 4614 19660 4620 19712
rect 4672 19700 4678 19712
rect 4985 19703 5043 19709
rect 4985 19700 4997 19703
rect 4672 19672 4997 19700
rect 4672 19660 4678 19672
rect 4985 19669 4997 19672
rect 5031 19669 5043 19703
rect 4985 19663 5043 19669
rect 5258 19660 5264 19712
rect 5316 19660 5322 19712
rect 6086 19660 6092 19712
rect 6144 19660 6150 19712
rect 8570 19660 8576 19712
rect 8628 19660 8634 19712
rect 8941 19703 8999 19709
rect 8941 19669 8953 19703
rect 8987 19700 8999 19703
rect 9140 19700 9168 19731
rect 9674 19728 9680 19780
rect 9732 19728 9738 19780
rect 9766 19728 9772 19780
rect 9824 19728 9830 19780
rect 9858 19728 9864 19780
rect 9916 19728 9922 19780
rect 9876 19700 9904 19728
rect 8987 19672 9904 19700
rect 8987 19669 8999 19672
rect 8941 19663 8999 19669
rect 10778 19660 10784 19712
rect 10836 19700 10842 19712
rect 11348 19700 11376 19799
rect 13998 19796 14004 19848
rect 14056 19796 14062 19848
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19805 14611 19839
rect 16684 19836 16712 19867
rect 17420 19836 17448 19867
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 19242 19864 19248 19916
rect 19300 19904 19306 19916
rect 19337 19907 19395 19913
rect 19337 19904 19349 19907
rect 19300 19876 19349 19904
rect 19300 19864 19306 19876
rect 19337 19873 19349 19876
rect 19383 19873 19395 19907
rect 19337 19867 19395 19873
rect 16684 19808 17448 19836
rect 14553 19799 14611 19805
rect 13170 19728 13176 19780
rect 13228 19768 13234 19780
rect 13814 19768 13820 19780
rect 13228 19740 13820 19768
rect 13228 19728 13234 19740
rect 13814 19728 13820 19740
rect 13872 19768 13878 19780
rect 14292 19768 14320 19796
rect 13872 19740 14320 19768
rect 13872 19728 13878 19740
rect 11514 19700 11520 19712
rect 10836 19672 11520 19700
rect 10836 19660 10842 19672
rect 11514 19660 11520 19672
rect 11572 19660 11578 19712
rect 12710 19660 12716 19712
rect 12768 19660 12774 19712
rect 13722 19660 13728 19712
rect 13780 19700 13786 19712
rect 13909 19703 13967 19709
rect 13909 19700 13921 19703
rect 13780 19672 13921 19700
rect 13780 19660 13786 19672
rect 13909 19669 13921 19672
rect 13955 19669 13967 19703
rect 14568 19700 14596 19799
rect 17129 19771 17187 19777
rect 17129 19737 17141 19771
rect 17175 19737 17187 19771
rect 17129 19731 17187 19737
rect 17221 19771 17279 19777
rect 17221 19737 17233 19771
rect 17267 19768 17279 19771
rect 17420 19768 17448 19808
rect 17494 19796 17500 19848
rect 17552 19796 17558 19848
rect 17586 19796 17592 19848
rect 17644 19796 17650 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 19444 19836 19472 19944
rect 20349 19941 20361 19975
rect 20395 19972 20407 19975
rect 20456 19972 20484 20000
rect 20395 19944 20484 19972
rect 20395 19941 20407 19944
rect 20349 19935 20407 19941
rect 20530 19932 20536 19984
rect 20588 19972 20594 19984
rect 23106 19972 23112 19984
rect 20588 19944 23112 19972
rect 20588 19932 20594 19944
rect 23106 19932 23112 19944
rect 23164 19932 23170 19984
rect 24412 19972 24440 20000
rect 24596 19981 24624 20012
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 24854 20000 24860 20052
rect 24912 20040 24918 20052
rect 24949 20043 25007 20049
rect 24949 20040 24961 20043
rect 24912 20012 24961 20040
rect 24912 20000 24918 20012
rect 24949 20009 24961 20012
rect 24995 20040 25007 20043
rect 25682 20040 25688 20052
rect 24995 20012 25688 20040
rect 24995 20009 25007 20012
rect 24949 20003 25007 20009
rect 25682 20000 25688 20012
rect 25740 20000 25746 20052
rect 26142 20000 26148 20052
rect 26200 20000 26206 20052
rect 27154 20000 27160 20052
rect 27212 20000 27218 20052
rect 27614 20000 27620 20052
rect 27672 20040 27678 20052
rect 27672 20012 28304 20040
rect 27672 20000 27678 20012
rect 24489 19975 24547 19981
rect 24489 19972 24501 19975
rect 24412 19944 24501 19972
rect 24489 19941 24501 19944
rect 24535 19941 24547 19975
rect 24489 19935 24547 19941
rect 24581 19975 24639 19981
rect 24581 19941 24593 19975
rect 24627 19941 24639 19975
rect 25133 19975 25191 19981
rect 25133 19972 25145 19975
rect 24581 19935 24639 19941
rect 24688 19944 25145 19972
rect 20073 19907 20131 19913
rect 20073 19873 20085 19907
rect 20119 19904 20131 19907
rect 20438 19904 20444 19916
rect 20119 19876 20444 19904
rect 20119 19873 20131 19876
rect 20073 19867 20131 19873
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 20542 19876 20852 19904
rect 20542 19836 20570 19876
rect 20824 19848 20852 19876
rect 20898 19864 20904 19916
rect 20956 19904 20962 19916
rect 21525 19907 21583 19913
rect 21525 19904 21537 19907
rect 20956 19876 21537 19904
rect 20956 19864 20962 19876
rect 21525 19873 21537 19876
rect 21571 19873 21583 19907
rect 21525 19867 21583 19873
rect 22094 19864 22100 19916
rect 22152 19904 22158 19916
rect 22997 19907 23055 19913
rect 22997 19904 23009 19907
rect 22152 19876 23009 19904
rect 22152 19864 22158 19876
rect 22997 19873 23009 19876
rect 23043 19873 23055 19907
rect 22997 19867 23055 19873
rect 23290 19864 23296 19916
rect 23348 19904 23354 19916
rect 23348 19876 23796 19904
rect 23348 19864 23354 19876
rect 17681 19799 17739 19805
rect 19168 19808 19472 19836
rect 19536 19808 20570 19836
rect 20717 19839 20775 19845
rect 17267 19740 17448 19768
rect 17512 19768 17540 19796
rect 17696 19768 17724 19799
rect 19168 19777 19196 19808
rect 17512 19740 17724 19768
rect 19153 19771 19211 19777
rect 17267 19737 17279 19740
rect 17221 19731 17279 19737
rect 19153 19737 19165 19771
rect 19199 19737 19211 19771
rect 19153 19731 19211 19737
rect 15838 19700 15844 19712
rect 14568 19672 15844 19700
rect 13909 19663 13967 19669
rect 15838 19660 15844 19672
rect 15896 19660 15902 19712
rect 15930 19660 15936 19712
rect 15988 19660 15994 19712
rect 17144 19700 17172 19731
rect 17497 19703 17555 19709
rect 17497 19700 17509 19703
rect 17144 19672 17509 19700
rect 17497 19669 17509 19672
rect 17543 19700 17555 19703
rect 19536 19700 19564 19808
rect 20717 19805 20729 19839
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 20165 19771 20223 19777
rect 20165 19737 20177 19771
rect 20211 19768 20223 19771
rect 20438 19768 20444 19780
rect 20211 19740 20444 19768
rect 20211 19737 20223 19740
rect 20165 19731 20223 19737
rect 20438 19728 20444 19740
rect 20496 19728 20502 19780
rect 20533 19771 20591 19777
rect 20533 19737 20545 19771
rect 20579 19737 20591 19771
rect 20732 19768 20760 19799
rect 20806 19796 20812 19848
rect 20864 19796 20870 19848
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21269 19839 21327 19845
rect 21269 19836 21281 19839
rect 21048 19808 21281 19836
rect 21048 19796 21054 19808
rect 21269 19805 21281 19808
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 22738 19796 22744 19848
rect 22796 19796 22802 19848
rect 23768 19836 23796 19876
rect 24302 19864 24308 19916
rect 24360 19904 24366 19916
rect 24397 19907 24455 19913
rect 24397 19904 24409 19907
rect 24360 19876 24409 19904
rect 24360 19864 24366 19876
rect 24397 19873 24409 19876
rect 24443 19873 24455 19907
rect 24397 19867 24455 19873
rect 24688 19836 24716 19944
rect 25133 19941 25145 19944
rect 25179 19941 25191 19975
rect 26160 19972 26188 20000
rect 25133 19935 25191 19941
rect 25976 19944 26188 19972
rect 27172 19972 27200 20000
rect 27810 19975 27868 19981
rect 27810 19972 27822 19975
rect 27172 19944 27822 19972
rect 24765 19907 24823 19913
rect 24765 19873 24777 19907
rect 24811 19873 24823 19907
rect 24765 19867 24823 19873
rect 23768 19808 24716 19836
rect 21174 19768 21180 19780
rect 20732 19740 21180 19768
rect 20533 19731 20591 19737
rect 17543 19672 19564 19700
rect 19981 19703 20039 19709
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 19981 19669 19993 19703
rect 20027 19700 20039 19703
rect 20070 19700 20076 19712
rect 20027 19672 20076 19700
rect 20027 19669 20039 19672
rect 19981 19663 20039 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20257 19703 20315 19709
rect 20257 19669 20269 19703
rect 20303 19700 20315 19703
rect 20548 19700 20576 19731
rect 21174 19728 21180 19740
rect 21232 19728 21238 19780
rect 24780 19768 24808 19867
rect 24854 19864 24860 19916
rect 24912 19864 24918 19916
rect 25976 19913 26004 19944
rect 27810 19941 27822 19944
rect 27856 19941 27868 19975
rect 28276 19972 28304 20012
rect 28350 20000 28356 20052
rect 28408 20040 28414 20052
rect 28721 20043 28779 20049
rect 28721 20040 28733 20043
rect 28408 20012 28733 20040
rect 28408 20000 28414 20012
rect 28721 20009 28733 20012
rect 28767 20009 28779 20043
rect 28721 20003 28779 20009
rect 28810 20000 28816 20052
rect 28868 20000 28874 20052
rect 29914 20000 29920 20052
rect 29972 20000 29978 20052
rect 28445 19975 28503 19981
rect 28276 19944 28396 19972
rect 27810 19935 27868 19941
rect 28368 19916 28396 19944
rect 28445 19941 28457 19975
rect 28491 19972 28503 19975
rect 28828 19972 28856 20000
rect 28491 19944 28856 19972
rect 29181 19975 29239 19981
rect 28491 19941 28503 19944
rect 28445 19935 28503 19941
rect 29181 19941 29193 19975
rect 29227 19972 29239 19975
rect 29362 19972 29368 19984
rect 29227 19944 29368 19972
rect 29227 19941 29239 19944
rect 29181 19935 29239 19941
rect 29362 19932 29368 19944
rect 29420 19972 29426 19984
rect 29638 19972 29644 19984
rect 29420 19944 29644 19972
rect 29420 19932 29426 19944
rect 29638 19932 29644 19944
rect 29696 19932 29702 19984
rect 25961 19907 26019 19913
rect 25961 19873 25973 19907
rect 26007 19873 26019 19907
rect 25961 19867 26019 19873
rect 26050 19864 26056 19916
rect 26108 19904 26114 19916
rect 26145 19907 26203 19913
rect 26145 19904 26157 19907
rect 26108 19876 26157 19904
rect 26108 19864 26114 19876
rect 26145 19873 26157 19876
rect 26191 19873 26203 19907
rect 28258 19904 28264 19916
rect 26145 19867 26203 19873
rect 26252 19876 28264 19904
rect 24872 19836 24900 19864
rect 26252 19836 26280 19876
rect 28258 19864 28264 19876
rect 28316 19864 28322 19916
rect 28350 19864 28356 19916
rect 28408 19864 28414 19916
rect 28537 19907 28595 19913
rect 28537 19873 28549 19907
rect 28583 19873 28595 19907
rect 28537 19867 28595 19873
rect 28629 19907 28687 19913
rect 28629 19873 28641 19907
rect 28675 19873 28687 19907
rect 28629 19867 28687 19873
rect 28813 19907 28871 19913
rect 28813 19873 28825 19907
rect 28859 19904 28871 19907
rect 29086 19904 29092 19916
rect 28859 19876 29092 19904
rect 28859 19873 28871 19876
rect 28813 19867 28871 19873
rect 24872 19808 26280 19836
rect 28077 19839 28135 19845
rect 28077 19805 28089 19839
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 23676 19740 24808 19768
rect 23676 19712 23704 19740
rect 20622 19700 20628 19712
rect 20303 19672 20628 19700
rect 20303 19669 20315 19672
rect 20257 19663 20315 19669
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 24118 19660 24124 19712
rect 24176 19660 24182 19712
rect 24210 19660 24216 19712
rect 24268 19660 24274 19712
rect 26694 19660 26700 19712
rect 26752 19660 26758 19712
rect 28092 19700 28120 19799
rect 28552 19768 28580 19867
rect 28644 19836 28672 19867
rect 29086 19864 29092 19876
rect 29144 19864 29150 19916
rect 29733 19907 29791 19913
rect 29733 19873 29745 19907
rect 29779 19873 29791 19907
rect 29733 19867 29791 19873
rect 29457 19839 29515 19845
rect 29457 19836 29469 19839
rect 28644 19808 29469 19836
rect 29457 19805 29469 19808
rect 29503 19805 29515 19839
rect 29457 19799 29515 19805
rect 29362 19768 29368 19780
rect 28552 19740 29368 19768
rect 29362 19728 29368 19740
rect 29420 19768 29426 19780
rect 29748 19768 29776 19867
rect 29420 19740 29776 19768
rect 29420 19728 29426 19740
rect 29270 19700 29276 19712
rect 28092 19672 29276 19700
rect 29270 19660 29276 19672
rect 29328 19660 29334 19712
rect 552 19610 31648 19632
rect 552 19558 4285 19610
rect 4337 19558 4349 19610
rect 4401 19558 4413 19610
rect 4465 19558 4477 19610
rect 4529 19558 4541 19610
rect 4593 19558 12059 19610
rect 12111 19558 12123 19610
rect 12175 19558 12187 19610
rect 12239 19558 12251 19610
rect 12303 19558 12315 19610
rect 12367 19558 19833 19610
rect 19885 19558 19897 19610
rect 19949 19558 19961 19610
rect 20013 19558 20025 19610
rect 20077 19558 20089 19610
rect 20141 19558 27607 19610
rect 27659 19558 27671 19610
rect 27723 19558 27735 19610
rect 27787 19558 27799 19610
rect 27851 19558 27863 19610
rect 27915 19558 31648 19610
rect 552 19536 31648 19558
rect 2958 19456 2964 19508
rect 3016 19496 3022 19508
rect 3237 19499 3295 19505
rect 3237 19496 3249 19499
rect 3016 19468 3249 19496
rect 3016 19456 3022 19468
rect 3237 19465 3249 19468
rect 3283 19465 3295 19499
rect 3237 19459 3295 19465
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 3513 19499 3571 19505
rect 3513 19496 3525 19499
rect 3384 19468 3525 19496
rect 3384 19456 3390 19468
rect 3513 19465 3525 19468
rect 3559 19465 3571 19499
rect 3513 19459 3571 19465
rect 3973 19499 4031 19505
rect 3973 19465 3985 19499
rect 4019 19496 4031 19499
rect 4614 19496 4620 19508
rect 4019 19468 4620 19496
rect 4019 19465 4031 19468
rect 3973 19459 4031 19465
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 5626 19456 5632 19508
rect 5684 19496 5690 19508
rect 7377 19499 7435 19505
rect 7377 19496 7389 19499
rect 5684 19468 7389 19496
rect 5684 19456 5690 19468
rect 7377 19465 7389 19468
rect 7423 19465 7435 19499
rect 7377 19459 7435 19465
rect 8662 19456 8668 19508
rect 8720 19496 8726 19508
rect 8941 19499 8999 19505
rect 8941 19496 8953 19499
rect 8720 19468 8953 19496
rect 8720 19456 8726 19468
rect 8941 19465 8953 19468
rect 8987 19465 8999 19499
rect 8941 19459 8999 19465
rect 9217 19499 9275 19505
rect 9217 19465 9229 19499
rect 9263 19496 9275 19499
rect 9306 19496 9312 19508
rect 9263 19468 9312 19496
rect 9263 19465 9275 19468
rect 9217 19459 9275 19465
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 9953 19499 10011 19505
rect 9953 19496 9965 19499
rect 9824 19468 9965 19496
rect 9824 19456 9830 19468
rect 9953 19465 9965 19468
rect 9999 19496 10011 19499
rect 11054 19496 11060 19508
rect 9999 19468 11060 19496
rect 9999 19465 10011 19468
rect 9953 19459 10011 19465
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11238 19456 11244 19508
rect 11296 19456 11302 19508
rect 11422 19456 11428 19508
rect 11480 19456 11486 19508
rect 12710 19456 12716 19508
rect 12768 19456 12774 19508
rect 13909 19499 13967 19505
rect 13909 19465 13921 19499
rect 13955 19496 13967 19499
rect 13998 19496 14004 19508
rect 13955 19468 14004 19496
rect 13955 19465 13967 19468
rect 13909 19459 13967 19465
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 16482 19496 16488 19508
rect 14200 19468 16488 19496
rect 3602 19388 3608 19440
rect 3660 19428 3666 19440
rect 4065 19431 4123 19437
rect 4065 19428 4077 19431
rect 3660 19400 4077 19428
rect 3660 19388 3666 19400
rect 4065 19397 4077 19400
rect 4111 19397 4123 19431
rect 4065 19391 4123 19397
rect 5902 19388 5908 19440
rect 5960 19428 5966 19440
rect 9674 19428 9680 19440
rect 5960 19400 7328 19428
rect 5960 19388 5966 19400
rect 3620 19332 4936 19360
rect 3421 19295 3479 19301
rect 3421 19261 3433 19295
rect 3467 19292 3479 19295
rect 3620 19292 3648 19332
rect 3467 19264 3648 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 3694 19252 3700 19304
rect 3752 19252 3758 19304
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 3973 19295 4031 19301
rect 3835 19264 3924 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 3896 19156 3924 19264
rect 3973 19261 3985 19295
rect 4019 19261 4031 19295
rect 3973 19255 4031 19261
rect 3988 19224 4016 19255
rect 4154 19252 4160 19304
rect 4212 19252 4218 19304
rect 4617 19295 4675 19301
rect 4617 19261 4629 19295
rect 4663 19292 4675 19295
rect 4798 19292 4804 19304
rect 4663 19264 4804 19292
rect 4663 19261 4675 19264
rect 4617 19255 4675 19261
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 4908 19301 4936 19332
rect 6472 19332 7052 19360
rect 6472 19304 6500 19332
rect 4893 19295 4951 19301
rect 4893 19261 4905 19295
rect 4939 19292 4951 19295
rect 4982 19292 4988 19304
rect 4939 19264 4988 19292
rect 4939 19261 4951 19264
rect 4893 19255 4951 19261
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 5166 19301 5172 19304
rect 5160 19292 5172 19301
rect 5127 19264 5172 19292
rect 5160 19255 5172 19264
rect 5166 19252 5172 19255
rect 5224 19252 5230 19304
rect 6086 19252 6092 19304
rect 6144 19292 6150 19304
rect 6365 19295 6423 19301
rect 6365 19292 6377 19295
rect 6144 19264 6377 19292
rect 6144 19252 6150 19264
rect 6365 19261 6377 19264
rect 6411 19261 6423 19295
rect 6365 19255 6423 19261
rect 6454 19252 6460 19304
rect 6512 19252 6518 19304
rect 6549 19295 6607 19301
rect 6549 19261 6561 19295
rect 6595 19292 6607 19295
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 6595 19264 6653 19292
rect 6595 19261 6607 19264
rect 6549 19255 6607 19261
rect 6641 19261 6653 19264
rect 6687 19292 6699 19295
rect 6730 19292 6736 19304
rect 6687 19264 6736 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 6914 19252 6920 19304
rect 6972 19252 6978 19304
rect 7024 19292 7052 19332
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7024 19264 7205 19292
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7300 19292 7328 19400
rect 7484 19400 9680 19428
rect 7484 19372 7512 19400
rect 9674 19388 9680 19400
rect 9732 19428 9738 19440
rect 10597 19431 10655 19437
rect 9732 19400 10180 19428
rect 9732 19388 9738 19400
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 8680 19332 9260 19360
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 7300 19264 7389 19292
rect 7193 19255 7251 19261
rect 7377 19261 7389 19264
rect 7423 19292 7435 19295
rect 8018 19292 8024 19304
rect 7423 19264 8024 19292
rect 7423 19261 7435 19264
rect 7377 19255 7435 19261
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 8570 19252 8576 19304
rect 8628 19252 8634 19304
rect 8680 19301 8708 19332
rect 8665 19295 8723 19301
rect 8665 19261 8677 19295
rect 8711 19261 8723 19295
rect 8665 19255 8723 19261
rect 8754 19252 8760 19304
rect 8812 19252 8818 19304
rect 8846 19252 8852 19304
rect 8904 19252 8910 19304
rect 9232 19301 9260 19332
rect 9416 19332 9996 19360
rect 9416 19304 9444 19332
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19261 8999 19295
rect 8941 19255 8999 19261
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19261 9183 19295
rect 9125 19255 9183 19261
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19292 9275 19295
rect 9306 19292 9312 19304
rect 9263 19264 9312 19292
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 4172 19224 4200 19252
rect 5258 19224 5264 19236
rect 3988 19196 4200 19224
rect 4264 19196 5264 19224
rect 4264 19156 4292 19196
rect 5258 19184 5264 19196
rect 5316 19184 5322 19236
rect 8588 19224 8616 19252
rect 8956 19224 8984 19255
rect 6380 19196 7236 19224
rect 8588 19196 8984 19224
rect 9140 19224 9168 19255
rect 9306 19252 9312 19264
rect 9364 19252 9370 19304
rect 9398 19252 9404 19304
rect 9456 19252 9462 19304
rect 9582 19252 9588 19304
rect 9640 19252 9646 19304
rect 9674 19252 9680 19304
rect 9732 19252 9738 19304
rect 9766 19252 9772 19304
rect 9824 19252 9830 19304
rect 9858 19252 9864 19304
rect 9916 19252 9922 19304
rect 9490 19224 9496 19236
rect 9140 19196 9496 19224
rect 3896 19128 4292 19156
rect 4338 19116 4344 19168
rect 4396 19156 4402 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4396 19128 4445 19156
rect 4396 19116 4402 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4433 19119 4491 19125
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 6380 19156 6408 19196
rect 6319 19128 6408 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 6454 19116 6460 19168
rect 6512 19116 6518 19168
rect 6822 19116 6828 19168
rect 6880 19116 6886 19168
rect 7098 19116 7104 19168
rect 7156 19116 7162 19168
rect 7208 19156 7236 19196
rect 9490 19184 9496 19196
rect 9548 19184 9554 19236
rect 8938 19156 8944 19168
rect 7208 19128 8944 19156
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9858 19116 9864 19168
rect 9916 19156 9922 19168
rect 9968 19156 9996 19332
rect 10042 19320 10048 19372
rect 10100 19320 10106 19372
rect 10152 19360 10180 19400
rect 10597 19397 10609 19431
rect 10643 19428 10655 19431
rect 11149 19431 11207 19437
rect 11149 19428 11161 19431
rect 10643 19400 11161 19428
rect 10643 19397 10655 19400
rect 10597 19391 10655 19397
rect 11149 19397 11161 19400
rect 11195 19428 11207 19431
rect 11440 19428 11468 19456
rect 11195 19400 11468 19428
rect 11195 19397 11207 19400
rect 11149 19391 11207 19397
rect 10689 19363 10747 19369
rect 10152 19332 10640 19360
rect 10152 19301 10180 19332
rect 10612 19301 10640 19332
rect 10689 19329 10701 19363
rect 10735 19360 10747 19363
rect 11054 19360 11060 19372
rect 10735 19332 11060 19360
rect 10735 19329 10747 19332
rect 10689 19323 10747 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 12728 19360 12756 19456
rect 13262 19388 13268 19440
rect 13320 19428 13326 19440
rect 13320 19400 13768 19428
rect 13320 19388 13326 19400
rect 13541 19363 13599 19369
rect 13541 19360 13553 19363
rect 12728 19332 13553 19360
rect 13541 19329 13553 19332
rect 13587 19329 13599 19363
rect 13541 19323 13599 19329
rect 13740 19360 13768 19400
rect 14200 19360 14228 19468
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 17586 19456 17592 19508
rect 17644 19456 17650 19508
rect 17865 19499 17923 19505
rect 17865 19465 17877 19499
rect 17911 19496 17923 19499
rect 19242 19496 19248 19508
rect 17911 19468 19248 19496
rect 17911 19465 17923 19468
rect 17865 19459 17923 19465
rect 18156 19437 18184 19468
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20070 19456 20076 19508
rect 20128 19456 20134 19508
rect 20162 19456 20168 19508
rect 20220 19496 20226 19508
rect 20220 19468 20570 19496
rect 20220 19456 20226 19468
rect 18049 19431 18107 19437
rect 18049 19428 18061 19431
rect 17926 19400 18061 19428
rect 15746 19360 15752 19372
rect 13740 19332 14228 19360
rect 15672 19332 15752 19360
rect 10137 19295 10195 19301
rect 10137 19261 10149 19295
rect 10183 19261 10195 19295
rect 10137 19255 10195 19261
rect 10321 19291 10379 19297
rect 10321 19257 10333 19291
rect 10367 19270 10379 19291
rect 10597 19295 10655 19301
rect 10367 19257 10450 19270
rect 10321 19251 10450 19257
rect 10597 19261 10609 19295
rect 10643 19292 10655 19295
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 10643 19264 11253 19292
rect 10643 19261 10655 19264
rect 10597 19255 10655 19261
rect 11241 19261 11253 19264
rect 11287 19261 11299 19295
rect 11241 19255 11299 19261
rect 11425 19295 11483 19301
rect 11425 19261 11437 19295
rect 11471 19292 11483 19295
rect 11514 19292 11520 19304
rect 11471 19264 11520 19292
rect 11471 19261 11483 19264
rect 11425 19255 11483 19261
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 13740 19295 13768 19332
rect 14277 19295 14335 19301
rect 13725 19289 13783 19295
rect 13725 19255 13737 19289
rect 13771 19255 13783 19289
rect 14277 19261 14289 19295
rect 14323 19292 14335 19295
rect 14323 19264 14780 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 10336 19242 10450 19251
rect 13725 19249 13783 19255
rect 10422 19156 10450 19242
rect 14752 19236 14780 19264
rect 10870 19184 10876 19236
rect 10928 19184 10934 19236
rect 10962 19184 10968 19236
rect 11020 19184 11026 19236
rect 11670 19227 11728 19233
rect 11670 19193 11682 19227
rect 11716 19193 11728 19227
rect 11670 19187 11728 19193
rect 9916 19128 10450 19156
rect 10505 19159 10563 19165
rect 9916 19116 9922 19128
rect 10505 19125 10517 19159
rect 10551 19156 10563 19159
rect 11685 19156 11713 19187
rect 13814 19184 13820 19236
rect 13872 19224 13878 19236
rect 14522 19227 14580 19233
rect 14522 19224 14534 19227
rect 13872 19196 14534 19224
rect 13872 19184 13878 19196
rect 14522 19193 14534 19196
rect 14568 19193 14580 19227
rect 14522 19187 14580 19193
rect 14734 19184 14740 19236
rect 14792 19184 14798 19236
rect 15672 19224 15700 19332
rect 15746 19320 15752 19332
rect 15804 19360 15810 19372
rect 15841 19363 15899 19369
rect 15841 19360 15853 19363
rect 15804 19332 15853 19360
rect 15804 19320 15810 19332
rect 15841 19329 15853 19332
rect 15887 19329 15899 19363
rect 15841 19323 15899 19329
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16025 19363 16083 19369
rect 16025 19360 16037 19363
rect 15988 19332 16037 19360
rect 15988 19320 15994 19332
rect 16025 19329 16037 19332
rect 16071 19329 16083 19363
rect 17770 19360 17776 19372
rect 16025 19323 16083 19329
rect 17420 19332 17776 19360
rect 17420 19301 17448 19332
rect 17770 19320 17776 19332
rect 17828 19360 17834 19372
rect 17926 19360 17954 19400
rect 18049 19397 18061 19400
rect 18095 19397 18107 19431
rect 18049 19391 18107 19397
rect 18141 19431 18199 19437
rect 18141 19397 18153 19431
rect 18187 19397 18199 19431
rect 18141 19391 18199 19397
rect 19058 19388 19064 19440
rect 19116 19428 19122 19440
rect 19705 19431 19763 19437
rect 19116 19400 19656 19428
rect 19116 19388 19122 19400
rect 17828 19332 17954 19360
rect 17828 19320 17834 19332
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 19628 19369 19656 19400
rect 19705 19397 19717 19431
rect 19751 19428 19763 19431
rect 20088 19428 20116 19456
rect 20349 19431 20407 19437
rect 20349 19428 20361 19431
rect 19751 19400 19932 19428
rect 20088 19400 20361 19428
rect 19751 19397 19763 19400
rect 19705 19391 19763 19397
rect 19613 19363 19671 19369
rect 18288 19332 19380 19360
rect 18288 19320 18294 19332
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 15028 19196 15700 19224
rect 17604 19224 17632 19255
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17736 19264 18061 19292
rect 17736 19252 17742 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18506 19252 18512 19304
rect 18564 19292 18570 19304
rect 18693 19295 18751 19301
rect 18693 19292 18705 19295
rect 18564 19264 18705 19292
rect 18564 19252 18570 19264
rect 18693 19261 18705 19264
rect 18739 19261 18751 19295
rect 18693 19255 18751 19261
rect 19150 19252 19156 19304
rect 19208 19252 19214 19304
rect 19352 19301 19380 19332
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 19613 19323 19671 19329
rect 19904 19304 19932 19400
rect 20349 19397 20361 19400
rect 20395 19397 20407 19431
rect 20349 19391 20407 19397
rect 20088 19332 20300 19360
rect 19337 19295 19395 19301
rect 19337 19261 19349 19295
rect 19383 19292 19395 19295
rect 19383 19264 19656 19292
rect 19383 19261 19395 19264
rect 19337 19255 19395 19261
rect 17604 19196 17816 19224
rect 15028 19168 15056 19196
rect 10551 19128 11713 19156
rect 12805 19159 12863 19165
rect 10551 19125 10563 19128
rect 10505 19119 10563 19125
rect 12805 19125 12817 19159
rect 12851 19156 12863 19159
rect 13538 19156 13544 19168
rect 12851 19128 13544 19156
rect 12851 19125 12863 19128
rect 12805 19119 12863 19125
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 15010 19116 15016 19168
rect 15068 19116 15074 19168
rect 15657 19159 15715 19165
rect 15657 19125 15669 19159
rect 15703 19156 15715 19159
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 15703 19128 16129 19156
rect 15703 19125 15715 19128
rect 15657 19119 15715 19125
rect 16117 19125 16129 19128
rect 16163 19125 16175 19159
rect 16117 19119 16175 19125
rect 16485 19159 16543 19165
rect 16485 19125 16497 19159
rect 16531 19156 16543 19159
rect 17126 19156 17132 19168
rect 16531 19128 17132 19156
rect 16531 19125 16543 19128
rect 16485 19119 16543 19125
rect 17126 19116 17132 19128
rect 17184 19116 17190 19168
rect 17788 19156 17816 19196
rect 17954 19184 17960 19236
rect 18012 19184 18018 19236
rect 18322 19184 18328 19236
rect 18380 19184 18386 19236
rect 19245 19227 19303 19233
rect 19245 19193 19257 19227
rect 19291 19224 19303 19227
rect 19429 19227 19487 19233
rect 19429 19224 19441 19227
rect 19291 19196 19441 19224
rect 19291 19193 19303 19196
rect 19245 19187 19303 19193
rect 19429 19193 19441 19196
rect 19475 19193 19487 19227
rect 19628 19224 19656 19264
rect 19702 19252 19708 19304
rect 19760 19292 19766 19304
rect 19797 19295 19855 19301
rect 19797 19292 19809 19295
rect 19760 19264 19809 19292
rect 19760 19252 19766 19264
rect 19797 19261 19809 19264
rect 19843 19261 19855 19295
rect 19797 19255 19855 19261
rect 19886 19252 19892 19304
rect 19944 19252 19950 19304
rect 20088 19292 20116 19332
rect 20272 19304 20300 19332
rect 19996 19264 20116 19292
rect 19996 19224 20024 19264
rect 20162 19252 20168 19304
rect 20220 19252 20226 19304
rect 20254 19252 20260 19304
rect 20312 19292 20318 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 20312 19264 20361 19292
rect 20312 19252 20318 19264
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 20349 19255 20407 19261
rect 20447 19295 20505 19301
rect 20447 19261 20459 19295
rect 20493 19292 20505 19295
rect 20542 19292 20570 19468
rect 20898 19456 20904 19508
rect 20956 19456 20962 19508
rect 20990 19456 20996 19508
rect 21048 19456 21054 19508
rect 22094 19456 22100 19508
rect 22152 19456 22158 19508
rect 23658 19456 23664 19508
rect 23716 19456 23722 19508
rect 24670 19456 24676 19508
rect 24728 19456 24734 19508
rect 24762 19456 24768 19508
rect 24820 19496 24826 19508
rect 27246 19496 27252 19508
rect 24820 19468 27252 19496
rect 24820 19456 24826 19468
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 28994 19456 29000 19508
rect 29052 19496 29058 19508
rect 30009 19499 30067 19505
rect 30009 19496 30021 19499
rect 29052 19468 30021 19496
rect 29052 19456 29058 19468
rect 30009 19465 30021 19468
rect 30055 19465 30067 19499
rect 30009 19459 30067 19465
rect 20806 19388 20812 19440
rect 20864 19388 20870 19440
rect 21008 19428 21036 19456
rect 21008 19400 22094 19428
rect 20824 19360 20852 19388
rect 20640 19332 21956 19360
rect 20640 19301 20668 19332
rect 20898 19302 20904 19304
rect 20732 19301 20904 19302
rect 20493 19264 20570 19292
rect 20625 19295 20683 19301
rect 20493 19261 20505 19264
rect 20447 19255 20505 19261
rect 20625 19261 20637 19295
rect 20671 19261 20683 19295
rect 20625 19255 20683 19261
rect 20717 19295 20904 19301
rect 20717 19261 20729 19295
rect 20763 19274 20904 19295
rect 20763 19261 20775 19274
rect 20717 19255 20775 19261
rect 20898 19252 20904 19274
rect 20956 19252 20962 19304
rect 21928 19301 21956 19332
rect 21913 19295 21971 19301
rect 21913 19261 21925 19295
rect 21959 19261 21971 19295
rect 21913 19255 21971 19261
rect 22066 19292 22094 19400
rect 29086 19388 29092 19440
rect 29144 19428 29150 19440
rect 29181 19431 29239 19437
rect 29181 19428 29193 19431
rect 29144 19400 29193 19428
rect 29144 19388 29150 19400
rect 29181 19397 29193 19400
rect 29227 19428 29239 19431
rect 29641 19431 29699 19437
rect 29641 19428 29653 19431
rect 29227 19400 29653 19428
rect 29227 19397 29239 19400
rect 29181 19391 29239 19397
rect 29641 19397 29653 19400
rect 29687 19397 29699 19431
rect 29641 19391 29699 19397
rect 24857 19363 24915 19369
rect 24857 19329 24869 19363
rect 24903 19360 24915 19363
rect 26050 19360 26056 19372
rect 24903 19332 26056 19360
rect 24903 19329 24915 19332
rect 24857 19323 24915 19329
rect 26050 19320 26056 19332
rect 26108 19320 26114 19372
rect 26804 19332 27108 19360
rect 22281 19295 22339 19301
rect 22281 19292 22293 19295
rect 22066 19264 22293 19292
rect 19628 19196 20024 19224
rect 20073 19227 20131 19233
rect 19429 19187 19487 19193
rect 20073 19193 20085 19227
rect 20119 19224 20131 19227
rect 20119 19196 20386 19224
rect 20119 19193 20131 19196
rect 20073 19187 20131 19193
rect 18138 19156 18144 19168
rect 17788 19128 18144 19156
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 19797 19159 19855 19165
rect 19797 19156 19809 19159
rect 19208 19128 19809 19156
rect 19208 19116 19214 19128
rect 19797 19125 19809 19128
rect 19843 19125 19855 19159
rect 19797 19119 19855 19125
rect 19886 19116 19892 19168
rect 19944 19156 19950 19168
rect 20162 19156 20168 19168
rect 19944 19128 20168 19156
rect 19944 19116 19950 19128
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 20358 19156 20386 19196
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 20358 19128 20545 19156
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 22066 19156 22094 19264
rect 22281 19261 22293 19264
rect 22327 19261 22339 19295
rect 22281 19255 22339 19261
rect 23750 19252 23756 19304
rect 23808 19252 23814 19304
rect 24118 19252 24124 19304
rect 24176 19252 24182 19304
rect 24486 19252 24492 19304
rect 24544 19252 24550 19304
rect 24946 19252 24952 19304
rect 25004 19252 25010 19304
rect 25038 19252 25044 19304
rect 25096 19252 25102 19304
rect 26694 19252 26700 19304
rect 26752 19252 26758 19304
rect 26804 19301 26832 19332
rect 26789 19295 26847 19301
rect 26789 19261 26801 19295
rect 26835 19261 26847 19295
rect 26789 19255 26847 19261
rect 26881 19295 26939 19301
rect 26881 19261 26893 19295
rect 26927 19261 26939 19295
rect 26881 19255 26939 19261
rect 26973 19295 27031 19301
rect 26973 19261 26985 19295
rect 27019 19261 27031 19295
rect 27080 19292 27108 19332
rect 29362 19320 29368 19372
rect 29420 19360 29426 19372
rect 29549 19363 29607 19369
rect 29549 19360 29561 19363
rect 29420 19346 29561 19360
rect 29420 19332 29460 19346
rect 29420 19320 29426 19332
rect 29273 19305 29331 19311
rect 27249 19295 27307 19301
rect 27249 19292 27261 19295
rect 27080 19264 27261 19292
rect 26973 19255 27031 19261
rect 27249 19261 27261 19264
rect 27295 19292 27307 19295
rect 27338 19292 27344 19304
rect 27295 19264 27344 19292
rect 27295 19261 27307 19264
rect 27249 19255 27307 19261
rect 22548 19227 22606 19233
rect 22548 19193 22560 19227
rect 22594 19224 22606 19227
rect 23014 19224 23020 19236
rect 22594 19196 23020 19224
rect 22594 19193 22606 19196
rect 22548 19187 22606 19193
rect 23014 19184 23020 19196
rect 23072 19184 23078 19236
rect 23768 19224 23796 19252
rect 24302 19224 24308 19236
rect 23768 19196 24308 19224
rect 24302 19184 24308 19196
rect 24360 19184 24366 19236
rect 24397 19227 24455 19233
rect 24397 19193 24409 19227
rect 24443 19224 24455 19227
rect 26712 19224 26740 19252
rect 24443 19196 26740 19224
rect 24443 19193 24455 19196
rect 24397 19187 24455 19193
rect 22278 19156 22284 19168
rect 22066 19128 22284 19156
rect 20533 19119 20591 19125
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 25222 19116 25228 19168
rect 25280 19116 25286 19168
rect 25774 19116 25780 19168
rect 25832 19156 25838 19168
rect 26804 19156 26832 19255
rect 26896 19168 26924 19255
rect 26988 19168 27016 19255
rect 27338 19252 27344 19264
rect 27396 19252 27402 19304
rect 28534 19292 28540 19304
rect 28184 19264 28540 19292
rect 27062 19184 27068 19236
rect 27120 19224 27126 19236
rect 28184 19224 28212 19264
rect 28534 19252 28540 19264
rect 28592 19292 28598 19304
rect 29273 19302 29285 19305
rect 29196 19292 29285 19302
rect 28592 19274 29285 19292
rect 28592 19264 29224 19274
rect 29273 19271 29285 19274
rect 29319 19271 29331 19305
rect 29454 19294 29460 19332
rect 29512 19332 29561 19346
rect 29512 19294 29518 19332
rect 29549 19329 29561 19332
rect 29595 19329 29607 19363
rect 29656 19360 29684 19391
rect 29656 19332 29776 19360
rect 29549 19323 29607 19329
rect 29748 19301 29776 19332
rect 29641 19295 29699 19301
rect 29641 19292 29653 19295
rect 29564 19282 29653 19292
rect 29273 19265 29331 19271
rect 28592 19252 28598 19264
rect 27120 19196 28212 19224
rect 27120 19184 27126 19196
rect 28994 19184 29000 19236
rect 29052 19184 29058 19236
rect 29104 19168 29132 19264
rect 29362 19184 29368 19236
rect 29420 19184 29426 19236
rect 29546 19230 29552 19282
rect 29604 19264 29653 19282
rect 29604 19230 29610 19264
rect 29641 19261 29653 19264
rect 29687 19261 29699 19295
rect 29641 19255 29699 19261
rect 29733 19295 29791 19301
rect 29733 19261 29745 19295
rect 29779 19261 29791 19295
rect 29733 19255 29791 19261
rect 30285 19295 30343 19301
rect 30285 19261 30297 19295
rect 30331 19261 30343 19295
rect 30285 19255 30343 19261
rect 30300 19224 30328 19255
rect 29656 19196 30328 19224
rect 25832 19128 26832 19156
rect 25832 19116 25838 19128
rect 26878 19116 26884 19168
rect 26936 19116 26942 19168
rect 26970 19116 26976 19168
rect 27028 19116 27034 19168
rect 27154 19116 27160 19168
rect 27212 19116 27218 19168
rect 27430 19116 27436 19168
rect 27488 19116 27494 19168
rect 29086 19116 29092 19168
rect 29144 19116 29150 19168
rect 29273 19159 29331 19165
rect 29273 19125 29285 19159
rect 29319 19156 29331 19159
rect 29454 19156 29460 19168
rect 29319 19128 29460 19156
rect 29319 19125 29331 19128
rect 29273 19119 29331 19125
rect 29454 19116 29460 19128
rect 29512 19116 29518 19168
rect 29546 19116 29552 19168
rect 29604 19156 29610 19168
rect 29656 19156 29684 19196
rect 29604 19128 29684 19156
rect 29604 19116 29610 19128
rect 29914 19116 29920 19168
rect 29972 19116 29978 19168
rect 30466 19116 30472 19168
rect 30524 19116 30530 19168
rect 552 19066 31808 19088
rect 552 19014 8172 19066
rect 8224 19014 8236 19066
rect 8288 19014 8300 19066
rect 8352 19014 8364 19066
rect 8416 19014 8428 19066
rect 8480 19014 15946 19066
rect 15998 19014 16010 19066
rect 16062 19014 16074 19066
rect 16126 19014 16138 19066
rect 16190 19014 16202 19066
rect 16254 19014 23720 19066
rect 23772 19014 23784 19066
rect 23836 19014 23848 19066
rect 23900 19014 23912 19066
rect 23964 19014 23976 19066
rect 24028 19014 31494 19066
rect 31546 19014 31558 19066
rect 31610 19014 31622 19066
rect 31674 19014 31686 19066
rect 31738 19014 31750 19066
rect 31802 19014 31808 19066
rect 552 18992 31808 19014
rect 5353 18955 5411 18961
rect 5353 18952 5365 18955
rect 3712 18924 5365 18952
rect 2406 18776 2412 18828
rect 2464 18816 2470 18828
rect 2869 18819 2927 18825
rect 2869 18816 2881 18819
rect 2464 18788 2881 18816
rect 2464 18776 2470 18788
rect 2869 18785 2881 18788
rect 2915 18785 2927 18819
rect 2869 18779 2927 18785
rect 3712 18806 3740 18924
rect 5353 18921 5365 18924
rect 5399 18952 5411 18955
rect 5442 18952 5448 18964
rect 5399 18924 5448 18952
rect 5399 18921 5411 18924
rect 5353 18915 5411 18921
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 6089 18955 6147 18961
rect 6089 18921 6101 18955
rect 6135 18952 6147 18955
rect 6135 18924 6960 18952
rect 6135 18921 6147 18924
rect 6089 18915 6147 18921
rect 4985 18887 5043 18893
rect 4985 18884 4997 18887
rect 4264 18856 4997 18884
rect 3789 18819 3847 18825
rect 3789 18806 3801 18819
rect 3712 18785 3801 18806
rect 3835 18785 3847 18819
rect 3712 18779 3847 18785
rect 2884 18612 2912 18779
rect 3712 18778 3823 18779
rect 3970 18776 3976 18828
rect 4028 18776 4034 18828
rect 4062 18776 4068 18828
rect 4120 18776 4126 18828
rect 3881 18751 3939 18757
rect 3881 18717 3893 18751
rect 3927 18748 3939 18751
rect 4264 18748 4292 18856
rect 4985 18853 4997 18856
rect 5031 18853 5043 18887
rect 4985 18847 5043 18853
rect 5626 18844 5632 18896
rect 5684 18844 5690 18896
rect 6932 18893 6960 18924
rect 7098 18912 7104 18964
rect 7156 18912 7162 18964
rect 9309 18955 9367 18961
rect 9309 18921 9321 18955
rect 9355 18952 9367 18955
rect 9398 18952 9404 18964
rect 9355 18924 9404 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 9398 18912 9404 18924
rect 9456 18912 9462 18964
rect 10137 18955 10195 18961
rect 10137 18952 10149 18955
rect 9661 18924 10149 18952
rect 6917 18887 6975 18893
rect 6917 18853 6929 18887
rect 6963 18853 6975 18887
rect 7116 18884 7144 18912
rect 7346 18887 7404 18893
rect 7346 18884 7358 18887
rect 7116 18856 7358 18884
rect 6917 18847 6975 18853
rect 7346 18853 7358 18856
rect 7392 18853 7404 18887
rect 7346 18847 7404 18853
rect 9030 18844 9036 18896
rect 9088 18844 9094 18896
rect 9661 18884 9689 18924
rect 10137 18921 10149 18924
rect 10183 18921 10195 18955
rect 10137 18915 10195 18921
rect 10689 18955 10747 18961
rect 10689 18921 10701 18955
rect 10735 18952 10747 18955
rect 10962 18952 10968 18964
rect 10735 18924 10968 18952
rect 10735 18921 10747 18924
rect 10689 18915 10747 18921
rect 10962 18912 10968 18924
rect 11020 18912 11026 18964
rect 11241 18955 11299 18961
rect 11241 18921 11253 18955
rect 11287 18952 11299 18955
rect 13814 18952 13820 18964
rect 11287 18924 13820 18952
rect 11287 18921 11299 18924
rect 11241 18915 11299 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 14642 18912 14648 18964
rect 14700 18912 14706 18964
rect 17770 18912 17776 18964
rect 17828 18912 17834 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18233 18955 18291 18961
rect 18233 18952 18245 18955
rect 18012 18924 18245 18952
rect 18012 18912 18018 18924
rect 18233 18921 18245 18924
rect 18279 18921 18291 18955
rect 18233 18915 18291 18921
rect 18322 18912 18328 18964
rect 18380 18952 18386 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 18380 18924 18521 18952
rect 18380 18912 18386 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 19245 18955 19303 18961
rect 19245 18921 19257 18955
rect 19291 18952 19303 18955
rect 19291 18924 21036 18952
rect 19291 18921 19303 18924
rect 19245 18915 19303 18921
rect 9600 18856 9689 18884
rect 12989 18887 13047 18893
rect 4525 18819 4583 18825
rect 4525 18785 4537 18819
rect 4571 18816 4583 18819
rect 4706 18816 4712 18828
rect 4571 18788 4712 18816
rect 4571 18785 4583 18788
rect 4525 18779 4583 18785
rect 4706 18776 4712 18788
rect 4764 18816 4770 18828
rect 5166 18816 5172 18828
rect 4764 18788 5172 18816
rect 4764 18776 4770 18788
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 5261 18819 5319 18825
rect 5261 18785 5273 18819
rect 5307 18816 5319 18819
rect 5350 18816 5356 18828
rect 5307 18788 5356 18816
rect 5307 18785 5319 18788
rect 5261 18779 5319 18785
rect 3927 18720 4292 18748
rect 4341 18751 4399 18757
rect 3927 18717 3939 18720
rect 3881 18711 3939 18717
rect 4341 18717 4353 18751
rect 4387 18748 4399 18751
rect 4614 18748 4620 18760
rect 4387 18720 4620 18748
rect 4387 18717 4399 18720
rect 4341 18711 4399 18717
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 4798 18708 4804 18760
rect 4856 18708 4862 18760
rect 5074 18708 5080 18760
rect 5132 18748 5138 18760
rect 5276 18748 5304 18779
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 5994 18776 6000 18828
rect 6052 18776 6058 18828
rect 6178 18776 6184 18828
rect 6236 18776 6242 18828
rect 6546 18776 6552 18828
rect 6604 18816 6610 18828
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 6604 18788 6653 18816
rect 6604 18776 6610 18788
rect 6641 18785 6653 18788
rect 6687 18785 6699 18819
rect 6641 18779 6699 18785
rect 8757 18819 8815 18825
rect 8757 18785 8769 18819
rect 8803 18785 8815 18819
rect 9048 18816 9076 18844
rect 9309 18819 9367 18825
rect 9309 18816 9321 18819
rect 9048 18788 9321 18816
rect 8757 18779 8815 18785
rect 9309 18785 9321 18788
rect 9355 18816 9367 18819
rect 9398 18816 9404 18828
rect 9355 18788 9404 18816
rect 9355 18785 9367 18788
rect 9309 18779 9367 18785
rect 5132 18720 5304 18748
rect 5132 18708 5138 18720
rect 6270 18708 6276 18760
rect 6328 18708 6334 18760
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 7098 18708 7104 18760
rect 7156 18708 7162 18760
rect 8772 18748 8800 18779
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 9600 18757 9628 18856
rect 12989 18853 13001 18887
rect 13035 18884 13047 18887
rect 13354 18884 13360 18896
rect 13035 18856 13360 18884
rect 13035 18853 13047 18856
rect 9674 18776 9680 18828
rect 9732 18776 9738 18828
rect 9858 18798 9864 18850
rect 9916 18838 9922 18850
rect 12989 18847 13047 18853
rect 9953 18841 10011 18847
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 13725 18887 13783 18893
rect 13725 18853 13737 18887
rect 13771 18884 13783 18887
rect 14550 18884 14556 18896
rect 13771 18856 14556 18884
rect 13771 18853 13783 18856
rect 13725 18847 13783 18853
rect 14550 18844 14556 18856
rect 14608 18844 14614 18896
rect 15194 18844 15200 18896
rect 15252 18884 15258 18896
rect 16362 18887 16420 18893
rect 16362 18884 16374 18887
rect 15252 18856 16374 18884
rect 15252 18844 15258 18856
rect 16362 18853 16374 18856
rect 16408 18853 16420 18887
rect 16362 18847 16420 18853
rect 9953 18838 9965 18841
rect 9916 18810 9965 18838
rect 9916 18798 9922 18810
rect 9953 18807 9965 18810
rect 9999 18807 10011 18841
rect 10069 18819 10127 18825
rect 10069 18816 10081 18819
rect 9953 18801 10011 18807
rect 10060 18785 10081 18816
rect 10115 18806 10127 18819
rect 10223 18819 10281 18825
rect 10115 18785 10180 18806
rect 10060 18778 10180 18785
rect 10223 18785 10235 18819
rect 10269 18785 10281 18819
rect 10223 18779 10281 18785
rect 9585 18751 9643 18757
rect 8772 18720 9444 18748
rect 3697 18683 3755 18689
rect 3697 18649 3709 18683
rect 3743 18680 3755 18683
rect 4157 18683 4215 18689
rect 4157 18680 4169 18683
rect 3743 18652 4169 18680
rect 3743 18649 3755 18652
rect 3697 18643 3755 18649
rect 4157 18649 4169 18652
rect 4203 18649 4215 18683
rect 5169 18683 5227 18689
rect 5169 18680 5181 18683
rect 4157 18643 4215 18649
rect 4264 18652 5181 18680
rect 4062 18612 4068 18624
rect 2884 18584 4068 18612
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 4264 18621 4292 18652
rect 4724 18624 4752 18652
rect 5169 18649 5181 18652
rect 5215 18649 5227 18683
rect 5169 18643 5227 18649
rect 5258 18640 5264 18692
rect 5316 18680 5322 18692
rect 5445 18683 5503 18689
rect 5445 18680 5457 18683
rect 5316 18652 5457 18680
rect 5316 18640 5322 18652
rect 5445 18649 5457 18652
rect 5491 18649 5503 18683
rect 5445 18643 5503 18649
rect 6549 18683 6607 18689
rect 6549 18649 6561 18683
rect 6595 18680 6607 18683
rect 6730 18680 6736 18692
rect 6595 18652 6736 18680
rect 6595 18649 6607 18652
rect 6549 18643 6607 18649
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 6822 18640 6828 18692
rect 6880 18680 6886 18692
rect 7116 18680 7144 18708
rect 6880 18652 7144 18680
rect 6880 18640 6886 18652
rect 8478 18640 8484 18692
rect 8536 18640 8542 18692
rect 9214 18640 9220 18692
rect 9272 18640 9278 18692
rect 9416 18689 9444 18720
rect 9585 18717 9597 18751
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 9950 18748 9956 18760
rect 9907 18720 9956 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 9401 18683 9459 18689
rect 9401 18649 9413 18683
rect 9447 18680 9459 18683
rect 9490 18680 9496 18692
rect 9447 18652 9496 18680
rect 9447 18649 9459 18652
rect 9401 18643 9459 18649
rect 9490 18640 9496 18652
rect 9548 18680 9554 18692
rect 10152 18680 10180 18778
rect 9548 18652 9674 18680
rect 9548 18640 9554 18652
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18581 4307 18615
rect 4249 18575 4307 18581
rect 4706 18572 4712 18624
rect 4764 18572 4770 18624
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 5077 18615 5135 18621
rect 5077 18612 5089 18615
rect 4948 18584 5089 18612
rect 4948 18572 4954 18584
rect 5077 18581 5089 18584
rect 5123 18581 5135 18615
rect 5077 18575 5135 18581
rect 6362 18572 6368 18624
rect 6420 18612 6426 18624
rect 6641 18615 6699 18621
rect 6641 18612 6653 18615
rect 6420 18584 6653 18612
rect 6420 18572 6426 18584
rect 6641 18581 6653 18584
rect 6687 18581 6699 18615
rect 6641 18575 6699 18581
rect 8941 18615 8999 18621
rect 8941 18581 8953 18615
rect 8987 18612 8999 18615
rect 9030 18612 9036 18624
rect 8987 18584 9036 18612
rect 8987 18581 8999 18584
rect 8941 18575 8999 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9646 18612 9674 18652
rect 10060 18652 10180 18680
rect 10238 18680 10266 18779
rect 10318 18776 10324 18828
rect 10376 18776 10382 18828
rect 10594 18776 10600 18828
rect 10652 18776 10658 18828
rect 10781 18819 10839 18825
rect 10781 18785 10793 18819
rect 10827 18785 10839 18819
rect 10781 18779 10839 18785
rect 10796 18748 10824 18779
rect 11054 18776 11060 18828
rect 11112 18776 11118 18828
rect 11698 18776 11704 18828
rect 11756 18776 11762 18828
rect 12713 18819 12771 18825
rect 12713 18785 12725 18819
rect 12759 18785 12771 18819
rect 12713 18779 12771 18785
rect 11716 18748 11744 18776
rect 10796 18720 11744 18748
rect 12728 18748 12756 18779
rect 12802 18776 12808 18828
rect 12860 18776 12866 18828
rect 13078 18776 13084 18828
rect 13136 18776 13142 18828
rect 13170 18776 13176 18828
rect 13228 18825 13234 18828
rect 13228 18816 13236 18825
rect 13228 18788 13273 18816
rect 13228 18779 13236 18788
rect 13228 18776 13234 18779
rect 13446 18776 13452 18828
rect 13504 18776 13510 18828
rect 13538 18776 13544 18828
rect 13596 18776 13602 18828
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18785 13875 18819
rect 13817 18779 13875 18785
rect 12986 18748 12992 18760
rect 12728 18720 12992 18748
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 10238 18652 10364 18680
rect 10060 18624 10088 18652
rect 10336 18624 10364 18652
rect 11146 18640 11152 18692
rect 11204 18680 11210 18692
rect 13832 18680 13860 18779
rect 13906 18776 13912 18828
rect 13964 18825 13970 18828
rect 13964 18819 14013 18825
rect 13964 18785 13967 18819
rect 14001 18816 14013 18819
rect 14001 18788 14136 18816
rect 14001 18785 14013 18788
rect 13964 18779 14013 18785
rect 13964 18776 13970 18779
rect 14108 18748 14136 18788
rect 14182 18776 14188 18828
rect 14240 18776 14246 18828
rect 17788 18825 17816 18912
rect 18340 18856 19472 18884
rect 14461 18819 14519 18825
rect 14461 18785 14473 18819
rect 14507 18816 14519 18819
rect 17773 18819 17831 18825
rect 14507 18788 17724 18816
rect 14507 18785 14519 18788
rect 14461 18779 14519 18785
rect 14108 18720 14688 18748
rect 14660 18692 14688 18720
rect 14734 18708 14740 18760
rect 14792 18748 14798 18760
rect 16117 18751 16175 18757
rect 16117 18748 16129 18751
rect 14792 18720 16129 18748
rect 14792 18708 14798 18720
rect 16117 18717 16129 18720
rect 16163 18717 16175 18751
rect 17696 18748 17724 18788
rect 17773 18785 17785 18819
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18816 18199 18819
rect 18230 18816 18236 18828
rect 18187 18788 18236 18816
rect 18187 18785 18199 18788
rect 18141 18779 18199 18785
rect 18230 18776 18236 18788
rect 18288 18776 18294 18828
rect 18340 18825 18368 18856
rect 19444 18828 19472 18856
rect 20070 18844 20076 18896
rect 20128 18884 20134 18896
rect 20625 18887 20683 18893
rect 20625 18884 20637 18887
rect 20128 18856 20637 18884
rect 20128 18844 20134 18856
rect 20625 18853 20637 18856
rect 20671 18853 20683 18887
rect 21008 18884 21036 18924
rect 23014 18912 23020 18964
rect 23072 18912 23078 18964
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 24029 18955 24087 18961
rect 24029 18952 24041 18955
rect 23532 18924 24041 18952
rect 23532 18912 23538 18924
rect 24029 18921 24041 18924
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 24305 18955 24363 18961
rect 24305 18921 24317 18955
rect 24351 18952 24363 18955
rect 24946 18952 24952 18964
rect 24351 18924 24952 18952
rect 24351 18921 24363 18924
rect 24305 18915 24363 18921
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 25492 18955 25550 18961
rect 25492 18921 25504 18955
rect 25538 18952 25550 18955
rect 26142 18952 26148 18964
rect 25538 18924 26148 18952
rect 25538 18921 25550 18924
rect 25492 18915 25550 18921
rect 26142 18912 26148 18924
rect 26200 18912 26206 18964
rect 26878 18912 26884 18964
rect 26936 18952 26942 18964
rect 27065 18955 27123 18961
rect 27065 18952 27077 18955
rect 26936 18924 27077 18952
rect 26936 18912 26942 18924
rect 27065 18921 27077 18924
rect 27111 18921 27123 18955
rect 27065 18915 27123 18921
rect 21514 18887 21572 18893
rect 21514 18884 21526 18887
rect 21008 18856 21526 18884
rect 20625 18847 20683 18853
rect 21514 18853 21526 18856
rect 21560 18853 21572 18887
rect 21514 18847 21572 18853
rect 24394 18844 24400 18896
rect 24452 18884 24458 18896
rect 25038 18884 25044 18896
rect 24452 18856 25044 18884
rect 24452 18844 24458 18856
rect 25038 18844 25044 18856
rect 25096 18844 25102 18896
rect 26513 18887 26571 18893
rect 26513 18884 26525 18887
rect 25884 18856 26525 18884
rect 25884 18828 25912 18856
rect 26513 18853 26525 18856
rect 26559 18853 26571 18887
rect 26513 18847 26571 18853
rect 18325 18819 18383 18825
rect 18325 18785 18337 18819
rect 18371 18785 18383 18819
rect 18325 18779 18383 18785
rect 18417 18819 18475 18825
rect 18417 18785 18429 18819
rect 18463 18816 18475 18819
rect 18506 18816 18512 18828
rect 18463 18788 18512 18816
rect 18463 18785 18475 18788
rect 18417 18779 18475 18785
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18966 18816 18972 18828
rect 18647 18788 18972 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18966 18776 18972 18788
rect 19024 18816 19030 18828
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 19024 18788 19073 18816
rect 19024 18776 19030 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 19150 18776 19156 18828
rect 19208 18816 19214 18828
rect 19208 18788 19380 18816
rect 19208 18776 19214 18788
rect 19242 18748 19248 18760
rect 17696 18720 19248 18748
rect 16117 18711 16175 18717
rect 19242 18708 19248 18720
rect 19300 18708 19306 18760
rect 19352 18748 19380 18788
rect 19426 18776 19432 18828
rect 19484 18776 19490 18828
rect 19613 18819 19671 18825
rect 19613 18785 19625 18819
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 19628 18748 19656 18779
rect 19794 18776 19800 18828
rect 19852 18776 19858 18828
rect 19886 18776 19892 18828
rect 19944 18816 19950 18828
rect 19981 18819 20039 18825
rect 19981 18816 19993 18819
rect 19944 18788 19993 18816
rect 19944 18776 19950 18788
rect 19981 18785 19993 18788
rect 20027 18785 20039 18819
rect 19981 18779 20039 18785
rect 20165 18819 20223 18825
rect 20165 18785 20177 18819
rect 20211 18816 20223 18819
rect 20533 18819 20591 18825
rect 20533 18816 20545 18819
rect 20211 18788 20545 18816
rect 20211 18785 20223 18788
rect 20165 18779 20223 18785
rect 20533 18785 20545 18788
rect 20579 18816 20591 18819
rect 20901 18819 20959 18825
rect 20901 18816 20913 18819
rect 20579 18788 20913 18816
rect 20579 18785 20591 18788
rect 20533 18779 20591 18785
rect 20901 18785 20913 18788
rect 20947 18816 20959 18819
rect 20990 18816 20996 18828
rect 20947 18788 20996 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 20990 18776 20996 18788
rect 21048 18816 21054 18828
rect 23201 18819 23259 18825
rect 21048 18788 23060 18816
rect 21048 18776 21054 18788
rect 19352 18720 19656 18748
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18748 19763 18751
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 19751 18720 20269 18748
rect 19751 18717 19763 18720
rect 19705 18711 19763 18717
rect 20257 18717 20269 18720
rect 20303 18717 20315 18751
rect 20257 18711 20315 18717
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18748 20499 18751
rect 21269 18751 21327 18757
rect 20487 18720 20944 18748
rect 20487 18717 20499 18720
rect 20441 18711 20499 18717
rect 11204 18652 13860 18680
rect 14093 18683 14151 18689
rect 11204 18640 11210 18652
rect 14093 18649 14105 18683
rect 14139 18680 14151 18683
rect 14277 18683 14335 18689
rect 14277 18680 14289 18683
rect 14139 18652 14289 18680
rect 14139 18649 14151 18652
rect 14093 18643 14151 18649
rect 14277 18649 14289 18652
rect 14323 18649 14335 18683
rect 14277 18643 14335 18649
rect 14642 18640 14648 18692
rect 14700 18640 14706 18692
rect 17497 18683 17555 18689
rect 17497 18649 17509 18683
rect 17543 18680 17555 18683
rect 19518 18680 19524 18692
rect 17543 18652 19524 18680
rect 17543 18649 17555 18652
rect 17497 18643 17555 18649
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 20806 18680 20812 18692
rect 20548 18652 20812 18680
rect 9769 18615 9827 18621
rect 9769 18612 9781 18615
rect 9646 18584 9781 18612
rect 9769 18581 9781 18584
rect 9815 18581 9827 18615
rect 9769 18575 9827 18581
rect 10042 18572 10048 18624
rect 10100 18572 10106 18624
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 10505 18615 10563 18621
rect 10505 18581 10517 18615
rect 10551 18612 10563 18615
rect 10870 18612 10876 18624
rect 10551 18584 10876 18612
rect 10551 18581 10563 18584
rect 10505 18575 10563 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 13354 18572 13360 18624
rect 13412 18572 13418 18624
rect 13446 18572 13452 18624
rect 13504 18612 13510 18624
rect 15010 18612 15016 18624
rect 13504 18584 15016 18612
rect 13504 18572 13510 18584
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 17586 18572 17592 18624
rect 17644 18572 17650 18624
rect 18874 18572 18880 18624
rect 18932 18572 18938 18624
rect 19058 18572 19064 18624
rect 19116 18612 19122 18624
rect 19886 18612 19892 18624
rect 19116 18584 19892 18612
rect 19116 18572 19122 18584
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 20548 18621 20576 18652
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 20916 18624 20944 18720
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 22646 18748 22652 18760
rect 21269 18711 21327 18717
rect 22296 18720 22652 18748
rect 20533 18615 20591 18621
rect 20533 18581 20545 18615
rect 20579 18581 20591 18615
rect 20533 18575 20591 18581
rect 20898 18572 20904 18624
rect 20956 18572 20962 18624
rect 20990 18572 20996 18624
rect 21048 18612 21054 18624
rect 21291 18612 21319 18711
rect 22296 18612 22324 18720
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 23032 18692 23060 18788
rect 23201 18785 23213 18819
rect 23247 18785 23259 18819
rect 25866 18816 25872 18828
rect 23201 18779 23259 18785
rect 24688 18788 25872 18816
rect 23216 18692 23244 18779
rect 24688 18760 24716 18788
rect 25866 18776 25872 18788
rect 25924 18776 25930 18828
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18816 26019 18819
rect 26050 18816 26056 18828
rect 26007 18788 26056 18816
rect 26007 18785 26019 18788
rect 25961 18779 26019 18785
rect 26050 18776 26056 18788
rect 26108 18776 26114 18828
rect 26528 18816 26556 18847
rect 26970 18844 26976 18896
rect 27028 18844 27034 18896
rect 27080 18884 27108 18915
rect 27430 18912 27436 18964
rect 27488 18952 27494 18964
rect 27617 18955 27675 18961
rect 27617 18952 27629 18955
rect 27488 18924 27629 18952
rect 27488 18912 27494 18924
rect 27617 18921 27629 18924
rect 27663 18921 27675 18955
rect 27617 18915 27675 18921
rect 28994 18912 29000 18964
rect 29052 18952 29058 18964
rect 29089 18955 29147 18961
rect 29089 18952 29101 18955
rect 29052 18924 29101 18952
rect 29052 18912 29058 18924
rect 29089 18921 29101 18924
rect 29135 18921 29147 18955
rect 29089 18915 29147 18921
rect 29362 18912 29368 18964
rect 29420 18912 29426 18964
rect 30466 18912 30472 18964
rect 30524 18912 30530 18964
rect 28813 18887 28871 18893
rect 27080 18856 27752 18884
rect 26988 18816 27016 18844
rect 27341 18819 27399 18825
rect 27341 18816 27353 18819
rect 26528 18788 27353 18816
rect 27341 18785 27353 18788
rect 27387 18785 27399 18819
rect 27341 18779 27399 18785
rect 27430 18776 27436 18828
rect 27488 18776 27494 18828
rect 27724 18825 27752 18856
rect 28813 18853 28825 18887
rect 28859 18884 28871 18887
rect 29380 18884 29408 18912
rect 28859 18856 29408 18884
rect 30484 18884 30512 18912
rect 30846 18887 30904 18893
rect 30846 18884 30858 18887
rect 30484 18856 30858 18884
rect 28859 18853 28871 18856
rect 28813 18847 28871 18853
rect 30846 18853 30858 18856
rect 30892 18853 30904 18887
rect 30846 18847 30904 18853
rect 27709 18819 27767 18825
rect 27709 18785 27721 18819
rect 27755 18816 27767 18819
rect 27982 18816 27988 18828
rect 27755 18788 27988 18816
rect 27755 18785 27767 18788
rect 27709 18779 27767 18785
rect 27982 18776 27988 18788
rect 28040 18776 28046 18828
rect 28718 18776 28724 18828
rect 28776 18776 28782 18828
rect 28902 18776 28908 18828
rect 28960 18776 28966 18828
rect 28994 18776 29000 18828
rect 29052 18776 29058 18828
rect 29178 18776 29184 18828
rect 29236 18816 29242 18828
rect 29365 18819 29423 18825
rect 29365 18816 29377 18819
rect 29236 18788 29377 18816
rect 29236 18776 29242 18788
rect 29365 18785 29377 18788
rect 29411 18785 29423 18819
rect 29365 18779 29423 18785
rect 29454 18776 29460 18828
rect 29512 18816 29518 18828
rect 31113 18819 31171 18825
rect 31113 18816 31125 18819
rect 29512 18788 31125 18816
rect 29512 18776 29518 18788
rect 31113 18785 31125 18788
rect 31159 18785 31171 18819
rect 31113 18779 31171 18785
rect 23566 18708 23572 18760
rect 23624 18748 23630 18760
rect 24188 18751 24246 18757
rect 24188 18748 24200 18751
rect 23624 18720 24200 18748
rect 23624 18708 23630 18720
rect 24188 18717 24200 18720
rect 24234 18717 24246 18751
rect 24188 18711 24246 18717
rect 24670 18708 24676 18760
rect 24728 18708 24734 18760
rect 26973 18751 27031 18757
rect 26973 18748 26985 18751
rect 24872 18720 26985 18748
rect 22554 18640 22560 18692
rect 22612 18680 22618 18692
rect 22741 18683 22799 18689
rect 22741 18680 22753 18683
rect 22612 18652 22753 18680
rect 22612 18640 22618 18652
rect 22741 18649 22753 18652
rect 22787 18649 22799 18683
rect 22741 18643 22799 18649
rect 23014 18640 23020 18692
rect 23072 18640 23078 18692
rect 23198 18640 23204 18692
rect 23256 18680 23262 18692
rect 23842 18680 23848 18692
rect 23256 18652 23848 18680
rect 23256 18640 23262 18652
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 24872 18680 24900 18720
rect 26973 18717 26985 18720
rect 27019 18717 27031 18751
rect 27448 18748 27476 18776
rect 26973 18711 27031 18717
rect 27172 18720 27476 18748
rect 27826 18751 27884 18757
rect 23952 18652 24900 18680
rect 21048 18584 22324 18612
rect 22649 18615 22707 18621
rect 21048 18572 21054 18584
rect 22649 18581 22661 18615
rect 22695 18612 22707 18615
rect 23952 18612 23980 18652
rect 25038 18640 25044 18692
rect 25096 18680 25102 18692
rect 26050 18680 26056 18692
rect 25096 18652 26056 18680
rect 25096 18640 25102 18652
rect 26050 18640 26056 18652
rect 26108 18680 26114 18692
rect 26513 18683 26571 18689
rect 26513 18680 26525 18683
rect 26108 18652 26525 18680
rect 26108 18640 26114 18652
rect 26513 18649 26525 18652
rect 26559 18680 26571 18683
rect 27172 18680 27200 18720
rect 27826 18717 27838 18751
rect 27872 18748 27884 18751
rect 27872 18720 29776 18748
rect 27872 18717 27884 18720
rect 27826 18711 27884 18717
rect 26559 18652 27200 18680
rect 26559 18649 26571 18652
rect 26513 18643 26571 18649
rect 27430 18640 27436 18692
rect 27488 18680 27494 18692
rect 27985 18683 28043 18689
rect 27985 18680 27997 18683
rect 27488 18652 27997 18680
rect 27488 18640 27494 18652
rect 27985 18649 27997 18652
rect 28031 18649 28043 18683
rect 27985 18643 28043 18649
rect 28350 18640 28356 18692
rect 28408 18680 28414 18692
rect 28810 18680 28816 18692
rect 28408 18652 28816 18680
rect 28408 18640 28414 18652
rect 28810 18640 28816 18652
rect 28868 18680 28874 18692
rect 28994 18680 29000 18692
rect 28868 18652 29000 18680
rect 28868 18640 28874 18652
rect 28994 18640 29000 18652
rect 29052 18640 29058 18692
rect 29748 18689 29776 18720
rect 29733 18683 29791 18689
rect 29733 18649 29745 18683
rect 29779 18649 29791 18683
rect 29733 18643 29791 18649
rect 22695 18584 23980 18612
rect 22695 18581 22707 18584
rect 22649 18575 22707 18581
rect 24486 18572 24492 18624
rect 24544 18612 24550 18624
rect 25317 18615 25375 18621
rect 25317 18612 25329 18615
rect 24544 18584 25329 18612
rect 24544 18572 24550 18584
rect 25317 18581 25329 18584
rect 25363 18612 25375 18615
rect 25406 18612 25412 18624
rect 25363 18584 25412 18612
rect 25363 18581 25375 18584
rect 25317 18575 25375 18581
rect 25406 18572 25412 18584
rect 25464 18572 25470 18624
rect 25501 18615 25559 18621
rect 25501 18581 25513 18615
rect 25547 18612 25559 18615
rect 25774 18612 25780 18624
rect 25547 18584 25780 18612
rect 25547 18581 25559 18584
rect 25501 18575 25559 18581
rect 25774 18572 25780 18584
rect 25832 18572 25838 18624
rect 25866 18572 25872 18624
rect 25924 18612 25930 18624
rect 26145 18615 26203 18621
rect 26145 18612 26157 18615
rect 25924 18584 26157 18612
rect 25924 18572 25930 18584
rect 26145 18581 26157 18584
rect 26191 18581 26203 18615
rect 26145 18575 26203 18581
rect 27246 18572 27252 18624
rect 27304 18572 27310 18624
rect 29546 18572 29552 18624
rect 29604 18572 29610 18624
rect 552 18522 31648 18544
rect 552 18470 4285 18522
rect 4337 18470 4349 18522
rect 4401 18470 4413 18522
rect 4465 18470 4477 18522
rect 4529 18470 4541 18522
rect 4593 18470 12059 18522
rect 12111 18470 12123 18522
rect 12175 18470 12187 18522
rect 12239 18470 12251 18522
rect 12303 18470 12315 18522
rect 12367 18470 19833 18522
rect 19885 18470 19897 18522
rect 19949 18470 19961 18522
rect 20013 18470 20025 18522
rect 20077 18470 20089 18522
rect 20141 18470 27607 18522
rect 27659 18470 27671 18522
rect 27723 18470 27735 18522
rect 27787 18470 27799 18522
rect 27851 18470 27863 18522
rect 27915 18470 31648 18522
rect 552 18448 31648 18470
rect 4246 18368 4252 18420
rect 4304 18408 4310 18420
rect 4985 18411 5043 18417
rect 4985 18408 4997 18411
rect 4304 18380 4997 18408
rect 4304 18368 4310 18380
rect 4985 18377 4997 18380
rect 5031 18377 5043 18411
rect 9306 18408 9312 18420
rect 4985 18371 5043 18377
rect 5276 18380 9312 18408
rect 4430 18232 4436 18284
rect 4488 18232 4494 18284
rect 4617 18275 4675 18281
rect 4617 18241 4629 18275
rect 4663 18272 4675 18275
rect 5276 18272 5304 18380
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 9398 18368 9404 18420
rect 9456 18368 9462 18420
rect 9766 18368 9772 18420
rect 9824 18408 9830 18420
rect 10226 18408 10232 18420
rect 9824 18380 10232 18408
rect 9824 18368 9830 18380
rect 5629 18343 5687 18349
rect 5629 18309 5641 18343
rect 5675 18340 5687 18343
rect 9416 18340 9444 18368
rect 9858 18340 9864 18352
rect 5675 18312 8294 18340
rect 9416 18312 9864 18340
rect 5675 18309 5687 18312
rect 5629 18303 5687 18309
rect 4663 18244 4844 18272
rect 4663 18241 4675 18244
rect 4617 18235 4675 18241
rect 4062 18164 4068 18216
rect 4120 18164 4126 18216
rect 4338 18164 4344 18216
rect 4396 18164 4402 18216
rect 4816 18213 4844 18244
rect 5000 18244 5304 18272
rect 5353 18275 5411 18281
rect 4709 18207 4767 18213
rect 4709 18173 4721 18207
rect 4755 18173 4767 18207
rect 4709 18167 4767 18173
rect 4801 18207 4859 18213
rect 4801 18173 4813 18207
rect 4847 18204 4859 18207
rect 4890 18204 4896 18216
rect 4847 18176 4896 18204
rect 4847 18173 4859 18176
rect 4801 18167 4859 18173
rect 4080 18136 4108 18164
rect 4724 18136 4752 18167
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 5000 18213 5028 18244
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 5902 18272 5908 18284
rect 5399 18244 5908 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 6086 18232 6092 18284
rect 6144 18272 6150 18284
rect 6914 18272 6920 18284
rect 6144 18244 6920 18272
rect 6144 18232 6150 18244
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7926 18272 7932 18284
rect 7392 18244 7932 18272
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18173 5043 18207
rect 4985 18167 5043 18173
rect 5442 18164 5448 18216
rect 5500 18164 5506 18216
rect 6181 18207 6239 18213
rect 6181 18173 6193 18207
rect 6227 18204 6239 18207
rect 6273 18207 6331 18213
rect 6273 18204 6285 18207
rect 6227 18176 6285 18204
rect 6227 18173 6239 18176
rect 6181 18167 6239 18173
rect 6273 18173 6285 18176
rect 6319 18173 6331 18207
rect 6273 18167 6331 18173
rect 6454 18164 6460 18216
rect 6512 18164 6518 18216
rect 7392 18213 7420 18244
rect 7926 18232 7932 18244
rect 7984 18232 7990 18284
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18204 7067 18207
rect 7377 18207 7435 18213
rect 7377 18204 7389 18207
rect 7055 18176 7389 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 7377 18173 7389 18176
rect 7423 18173 7435 18207
rect 7377 18167 7435 18173
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7558 18204 7564 18216
rect 7515 18176 7564 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 8266 18204 8294 18312
rect 9858 18300 9864 18312
rect 9916 18300 9922 18352
rect 9968 18349 9996 18380
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 10502 18368 10508 18420
rect 10560 18408 10566 18420
rect 10689 18411 10747 18417
rect 10689 18408 10701 18411
rect 10560 18380 10701 18408
rect 10560 18368 10566 18380
rect 10689 18377 10701 18380
rect 10735 18377 10747 18411
rect 12253 18411 12311 18417
rect 10689 18371 10747 18377
rect 10796 18380 11836 18408
rect 9953 18343 10011 18349
rect 9953 18309 9965 18343
rect 9999 18309 10011 18343
rect 9953 18303 10011 18309
rect 10045 18343 10103 18349
rect 10045 18309 10057 18343
rect 10091 18340 10103 18343
rect 10318 18340 10324 18352
rect 10091 18312 10324 18340
rect 10091 18309 10103 18312
rect 10045 18303 10103 18309
rect 10318 18300 10324 18312
rect 10376 18340 10382 18352
rect 10796 18340 10824 18380
rect 10376 18312 10824 18340
rect 10376 18300 10382 18312
rect 10870 18300 10876 18352
rect 10928 18300 10934 18352
rect 11808 18340 11836 18380
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 13078 18408 13084 18420
rect 12299 18380 13084 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 16298 18408 16304 18420
rect 13188 18380 16304 18408
rect 11808 18312 12388 18340
rect 9876 18204 9904 18300
rect 10134 18232 10140 18284
rect 10192 18232 10198 18284
rect 10594 18272 10600 18284
rect 10428 18244 10600 18272
rect 10042 18204 10048 18216
rect 8266 18176 9720 18204
rect 9876 18176 10048 18204
rect 5074 18136 5080 18148
rect 4080 18108 5080 18136
rect 5074 18096 5080 18108
rect 5132 18096 5138 18148
rect 5166 18096 5172 18148
rect 5224 18136 5230 18148
rect 7193 18139 7251 18145
rect 7193 18136 7205 18139
rect 5224 18108 7205 18136
rect 5224 18096 5230 18108
rect 7193 18105 7205 18108
rect 7239 18105 7251 18139
rect 7193 18099 7251 18105
rect 9582 18096 9588 18148
rect 9640 18096 9646 18148
rect 4706 18028 4712 18080
rect 4764 18028 4770 18080
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 5258 18068 5264 18080
rect 4856 18040 5264 18068
rect 4856 18028 4862 18040
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6365 18071 6423 18077
rect 6365 18068 6377 18071
rect 6328 18040 6377 18068
rect 6328 18028 6334 18040
rect 6365 18037 6377 18040
rect 6411 18037 6423 18071
rect 6365 18031 6423 18037
rect 6825 18071 6883 18077
rect 6825 18037 6837 18071
rect 6871 18068 6883 18071
rect 7006 18068 7012 18080
rect 6871 18040 7012 18068
rect 6871 18037 6883 18040
rect 6825 18031 6883 18037
rect 7006 18028 7012 18040
rect 7064 18068 7070 18080
rect 7466 18068 7472 18080
rect 7064 18040 7472 18068
rect 7064 18028 7070 18040
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18068 7711 18071
rect 7742 18068 7748 18080
rect 7699 18040 7748 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 8018 18028 8024 18080
rect 8076 18068 8082 18080
rect 9600 18068 9628 18096
rect 8076 18040 9628 18068
rect 9692 18068 9720 18176
rect 10042 18164 10048 18176
rect 10100 18204 10106 18216
rect 10428 18213 10456 18244
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 10778 18232 10784 18284
rect 10836 18232 10842 18284
rect 10888 18272 10916 18300
rect 10888 18244 11008 18272
rect 10413 18207 10471 18213
rect 10413 18204 10425 18207
rect 10100 18176 10425 18204
rect 10100 18164 10106 18176
rect 10413 18173 10425 18176
rect 10459 18173 10471 18207
rect 10413 18167 10471 18173
rect 10505 18207 10563 18213
rect 10505 18173 10517 18207
rect 10551 18200 10563 18207
rect 10551 18173 10640 18200
rect 10505 18172 10640 18173
rect 10505 18167 10563 18172
rect 9766 18096 9772 18148
rect 9824 18096 9830 18148
rect 10612 18136 10640 18172
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 10796 18204 10824 18232
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 10796 18176 10885 18204
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10980 18204 11008 18244
rect 12360 18213 12388 18312
rect 12434 18300 12440 18352
rect 12492 18340 12498 18352
rect 13188 18340 13216 18380
rect 16298 18368 16304 18380
rect 16356 18368 16362 18420
rect 17678 18368 17684 18420
rect 17736 18408 17742 18420
rect 18417 18411 18475 18417
rect 18417 18408 18429 18411
rect 17736 18380 18429 18408
rect 17736 18368 17742 18380
rect 18417 18377 18429 18380
rect 18463 18377 18475 18411
rect 18417 18371 18475 18377
rect 12492 18312 13216 18340
rect 12492 18300 12498 18312
rect 16666 18300 16672 18352
rect 16724 18340 16730 18352
rect 18230 18340 18236 18352
rect 16724 18312 18236 18340
rect 16724 18300 16730 18312
rect 18230 18300 18236 18312
rect 18288 18300 18294 18352
rect 14734 18232 14740 18284
rect 14792 18232 14798 18284
rect 18432 18272 18460 18371
rect 18966 18368 18972 18420
rect 19024 18368 19030 18420
rect 19242 18368 19248 18420
rect 19300 18368 19306 18420
rect 19702 18368 19708 18420
rect 19760 18408 19766 18420
rect 19981 18411 20039 18417
rect 19981 18408 19993 18411
rect 19760 18380 19993 18408
rect 19760 18368 19766 18380
rect 19981 18377 19993 18380
rect 20027 18377 20039 18411
rect 19981 18371 20039 18377
rect 20625 18411 20683 18417
rect 20625 18377 20637 18411
rect 20671 18408 20683 18411
rect 26513 18411 26571 18417
rect 26513 18408 26525 18411
rect 20671 18380 26525 18408
rect 20671 18377 20683 18380
rect 20625 18371 20683 18377
rect 26513 18377 26525 18380
rect 26559 18377 26571 18411
rect 26513 18371 26571 18377
rect 26878 18368 26884 18420
rect 26936 18368 26942 18420
rect 26973 18411 27031 18417
rect 26973 18377 26985 18411
rect 27019 18408 27031 18411
rect 27246 18408 27252 18420
rect 27019 18380 27252 18408
rect 27019 18377 27031 18380
rect 26973 18371 27031 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27430 18368 27436 18420
rect 27488 18368 27494 18420
rect 28718 18408 28724 18420
rect 28552 18380 28724 18408
rect 18984 18340 19012 18368
rect 19153 18343 19211 18349
rect 19153 18340 19165 18343
rect 18984 18312 19165 18340
rect 19153 18309 19165 18312
rect 19199 18309 19211 18343
rect 19153 18303 19211 18309
rect 19260 18272 19288 18368
rect 20254 18300 20260 18352
rect 20312 18300 20318 18352
rect 20806 18300 20812 18352
rect 20864 18340 20870 18352
rect 22646 18340 22652 18352
rect 20864 18312 22652 18340
rect 20864 18300 20870 18312
rect 19334 18272 19340 18284
rect 18432 18244 19012 18272
rect 19260 18244 19340 18272
rect 11129 18207 11187 18213
rect 11129 18204 11141 18207
rect 10980 18176 11141 18204
rect 10873 18167 10931 18173
rect 11129 18173 11141 18176
rect 11175 18173 11187 18207
rect 11129 18167 11187 18173
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 14752 18204 14780 18232
rect 18984 18213 19012 18244
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19444 18244 21128 18272
rect 13587 18176 14780 18204
rect 18233 18207 18291 18213
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 18233 18173 18245 18207
rect 18279 18173 18291 18207
rect 18233 18167 18291 18173
rect 18877 18207 18935 18213
rect 18877 18173 18889 18207
rect 18923 18173 18935 18207
rect 18877 18167 18935 18173
rect 18969 18207 19027 18213
rect 18969 18173 18981 18207
rect 19015 18204 19027 18207
rect 19061 18207 19119 18213
rect 19061 18204 19073 18207
rect 19015 18176 19073 18204
rect 19015 18173 19027 18176
rect 18969 18167 19027 18173
rect 19061 18173 19073 18176
rect 19107 18204 19119 18207
rect 19242 18204 19248 18216
rect 19107 18176 19248 18204
rect 19107 18173 19119 18176
rect 19061 18167 19119 18173
rect 10962 18136 10968 18148
rect 10612 18108 10968 18136
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 11514 18096 11520 18148
rect 11572 18096 11578 18148
rect 13786 18139 13844 18145
rect 13786 18136 13798 18139
rect 12544 18108 13798 18136
rect 11532 18068 11560 18096
rect 12544 18077 12572 18108
rect 13786 18105 13798 18108
rect 13832 18105 13844 18139
rect 13786 18099 13844 18105
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 17310 18136 17316 18148
rect 14608 18108 17316 18136
rect 14608 18096 14614 18108
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 9692 18040 11560 18068
rect 12529 18071 12587 18077
rect 8076 18028 8082 18040
rect 12529 18037 12541 18071
rect 12575 18037 12587 18071
rect 12529 18031 12587 18037
rect 14918 18028 14924 18080
rect 14976 18028 14982 18080
rect 18248 18068 18276 18167
rect 18690 18096 18696 18148
rect 18748 18096 18754 18148
rect 18892 18136 18920 18167
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 19444 18213 19472 18244
rect 20272 18216 20300 18244
rect 19429 18207 19487 18213
rect 19429 18173 19441 18207
rect 19475 18173 19487 18207
rect 19429 18167 19487 18173
rect 19607 18207 19665 18213
rect 19607 18173 19619 18207
rect 19653 18204 19665 18207
rect 19702 18204 19708 18216
rect 19653 18176 19708 18204
rect 19653 18173 19665 18176
rect 19607 18167 19665 18173
rect 19702 18164 19708 18176
rect 19760 18164 19766 18216
rect 20254 18164 20260 18216
rect 20312 18164 20318 18216
rect 20530 18164 20536 18216
rect 20588 18164 20594 18216
rect 20625 18207 20683 18213
rect 20625 18173 20637 18207
rect 20671 18204 20683 18207
rect 20806 18204 20812 18216
rect 20671 18176 20812 18204
rect 20671 18173 20683 18176
rect 20625 18167 20683 18173
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 20898 18164 20904 18216
rect 20956 18164 20962 18216
rect 21100 18213 21128 18244
rect 21085 18207 21143 18213
rect 21085 18173 21097 18207
rect 21131 18204 21143 18207
rect 22094 18204 22100 18216
rect 21131 18176 22100 18204
rect 21131 18173 21143 18176
rect 21085 18167 21143 18173
rect 22094 18164 22100 18176
rect 22152 18164 22158 18216
rect 22204 18213 22232 18312
rect 22646 18300 22652 18312
rect 22704 18300 22710 18352
rect 22741 18343 22799 18349
rect 22741 18309 22753 18343
rect 22787 18340 22799 18343
rect 23017 18343 23075 18349
rect 23017 18340 23029 18343
rect 22787 18312 23029 18340
rect 22787 18309 22799 18312
rect 22741 18303 22799 18309
rect 23017 18309 23029 18312
rect 23063 18340 23075 18343
rect 23063 18312 23152 18340
rect 23063 18309 23075 18312
rect 23017 18303 23075 18309
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18272 22339 18275
rect 22833 18275 22891 18281
rect 22833 18272 22845 18275
rect 22327 18244 22845 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 22833 18241 22845 18244
rect 22879 18241 22891 18275
rect 23124 18272 23152 18312
rect 24946 18300 24952 18352
rect 25004 18340 25010 18352
rect 26237 18343 26295 18349
rect 26237 18340 26249 18343
rect 25004 18312 26249 18340
rect 25004 18300 25010 18312
rect 26237 18309 26249 18312
rect 26283 18340 26295 18343
rect 26896 18340 26924 18368
rect 26283 18312 26924 18340
rect 26283 18309 26295 18312
rect 26237 18303 26295 18309
rect 27338 18300 27344 18352
rect 27396 18300 27402 18352
rect 23198 18272 23204 18284
rect 23124 18244 23204 18272
rect 22833 18235 22891 18241
rect 23198 18232 23204 18244
rect 23256 18232 23262 18284
rect 23842 18232 23848 18284
rect 23900 18272 23906 18284
rect 26881 18275 26939 18281
rect 23900 18244 26464 18272
rect 23900 18232 23906 18244
rect 26436 18216 26464 18244
rect 26881 18241 26893 18275
rect 26927 18272 26939 18275
rect 27448 18272 27476 18368
rect 26927 18244 27476 18272
rect 28552 18272 28580 18380
rect 28718 18368 28724 18380
rect 28776 18408 28782 18420
rect 29454 18408 29460 18420
rect 28776 18380 29460 18408
rect 28776 18368 28782 18380
rect 29454 18368 29460 18380
rect 29512 18368 29518 18420
rect 29546 18368 29552 18420
rect 29604 18368 29610 18420
rect 28629 18343 28687 18349
rect 28629 18309 28641 18343
rect 28675 18340 28687 18343
rect 29178 18340 29184 18352
rect 28675 18312 29184 18340
rect 28675 18309 28687 18312
rect 28629 18303 28687 18309
rect 29178 18300 29184 18312
rect 29236 18340 29242 18352
rect 29273 18343 29331 18349
rect 29273 18340 29285 18343
rect 29236 18312 29285 18340
rect 29236 18300 29242 18312
rect 29273 18309 29285 18312
rect 29319 18309 29331 18343
rect 29273 18303 29331 18309
rect 28813 18275 28871 18281
rect 28552 18244 28764 18272
rect 26927 18241 26939 18244
rect 26881 18235 26939 18241
rect 22189 18207 22247 18213
rect 22189 18173 22201 18207
rect 22235 18173 22247 18207
rect 22189 18167 22247 18173
rect 22373 18207 22431 18213
rect 22373 18173 22385 18207
rect 22419 18204 22431 18207
rect 22554 18204 22560 18216
rect 22419 18176 22560 18204
rect 22419 18173 22431 18176
rect 22373 18167 22431 18173
rect 22554 18164 22560 18176
rect 22612 18164 22618 18216
rect 22646 18164 22652 18216
rect 22704 18164 22710 18216
rect 22741 18207 22799 18213
rect 22741 18173 22753 18207
rect 22787 18204 22799 18207
rect 23014 18204 23020 18216
rect 22787 18176 23020 18204
rect 22787 18173 22799 18176
rect 22741 18167 22799 18173
rect 23014 18164 23020 18176
rect 23072 18204 23078 18216
rect 23109 18207 23167 18213
rect 23109 18204 23121 18207
rect 23072 18176 23121 18204
rect 23072 18164 23078 18176
rect 23109 18173 23121 18176
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18200 23443 18207
rect 23566 18200 23572 18216
rect 23431 18173 23572 18200
rect 23385 18172 23572 18173
rect 23385 18167 23443 18172
rect 23566 18164 23572 18172
rect 23624 18164 23630 18216
rect 24213 18207 24271 18213
rect 24213 18173 24225 18207
rect 24259 18204 24271 18207
rect 24394 18204 24400 18216
rect 24259 18176 24400 18204
rect 24259 18173 24271 18176
rect 24213 18167 24271 18173
rect 24394 18164 24400 18176
rect 24452 18164 24458 18216
rect 24581 18207 24639 18213
rect 24581 18173 24593 18207
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 19337 18139 19395 18145
rect 18892 18108 19104 18136
rect 18966 18068 18972 18080
rect 18248 18040 18972 18068
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 19076 18077 19104 18108
rect 19337 18105 19349 18139
rect 19383 18136 19395 18139
rect 19521 18139 19579 18145
rect 19521 18136 19533 18139
rect 19383 18108 19533 18136
rect 19383 18105 19395 18108
rect 19337 18099 19395 18105
rect 19521 18105 19533 18108
rect 19567 18105 19579 18139
rect 19521 18099 19579 18105
rect 20993 18139 21051 18145
rect 20993 18105 21005 18139
rect 21039 18136 21051 18139
rect 22465 18139 22523 18145
rect 22465 18136 22477 18139
rect 21039 18108 22477 18136
rect 21039 18105 21051 18108
rect 20993 18099 21051 18105
rect 22465 18105 22477 18108
rect 22511 18105 22523 18139
rect 22465 18099 22523 18105
rect 23124 18108 23612 18136
rect 19061 18071 19119 18077
rect 19061 18037 19073 18071
rect 19107 18068 19119 18071
rect 19426 18068 19432 18080
rect 19107 18040 19432 18068
rect 19107 18037 19119 18040
rect 19061 18031 19119 18037
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 23124 18077 23152 18108
rect 23584 18080 23612 18108
rect 24302 18096 24308 18148
rect 24360 18096 24366 18148
rect 24596 18136 24624 18167
rect 24946 18164 24952 18216
rect 25004 18164 25010 18216
rect 26053 18207 26111 18213
rect 26053 18173 26065 18207
rect 26099 18204 26111 18207
rect 26142 18204 26148 18216
rect 26099 18176 26148 18204
rect 26099 18173 26111 18176
rect 26053 18167 26111 18173
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 26418 18164 26424 18216
rect 26476 18164 26482 18216
rect 26786 18164 26792 18216
rect 26844 18164 26850 18216
rect 27154 18164 27160 18216
rect 27212 18204 27218 18216
rect 27249 18207 27307 18213
rect 27249 18204 27261 18207
rect 27212 18176 27261 18204
rect 27212 18164 27218 18176
rect 27249 18173 27261 18176
rect 27295 18204 27307 18207
rect 27525 18207 27583 18213
rect 27525 18204 27537 18207
rect 27295 18176 27537 18204
rect 27295 18173 27307 18176
rect 27249 18167 27307 18173
rect 27525 18173 27537 18176
rect 27571 18173 27583 18207
rect 27525 18167 27583 18173
rect 28534 18164 28540 18216
rect 28592 18164 28598 18216
rect 28736 18204 28764 18244
rect 28813 18241 28825 18275
rect 28859 18272 28871 18275
rect 29454 18272 29460 18284
rect 28859 18244 29460 18272
rect 28859 18241 28871 18244
rect 28813 18235 28871 18241
rect 29454 18232 29460 18244
rect 29512 18232 29518 18284
rect 29564 18272 29592 18368
rect 29564 18244 29684 18272
rect 29181 18207 29239 18213
rect 29181 18204 29193 18207
rect 28736 18176 29193 18204
rect 29181 18173 29193 18176
rect 29227 18173 29239 18207
rect 29181 18167 29239 18173
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18173 29331 18207
rect 29273 18167 29331 18173
rect 24670 18136 24676 18148
rect 24596 18108 24676 18136
rect 24670 18096 24676 18108
rect 24728 18136 24734 18148
rect 24728 18108 24992 18136
rect 24728 18096 24734 18108
rect 23109 18071 23167 18077
rect 23109 18037 23121 18071
rect 23155 18037 23167 18071
rect 23109 18031 23167 18037
rect 23198 18028 23204 18080
rect 23256 18028 23262 18080
rect 23566 18028 23572 18080
rect 23624 18028 23630 18080
rect 24213 18071 24271 18077
rect 24213 18037 24225 18071
rect 24259 18068 24271 18071
rect 24320 18068 24348 18096
rect 24964 18080 24992 18108
rect 27172 18108 28948 18136
rect 24259 18040 24348 18068
rect 24259 18037 24271 18040
rect 24213 18031 24271 18037
rect 24946 18028 24952 18080
rect 25004 18028 25010 18080
rect 27172 18077 27200 18108
rect 27157 18071 27215 18077
rect 27157 18037 27169 18071
rect 27203 18037 27215 18071
rect 28920 18068 28948 18108
rect 28994 18096 29000 18148
rect 29052 18096 29058 18148
rect 29086 18096 29092 18148
rect 29144 18136 29150 18148
rect 29288 18136 29316 18167
rect 29362 18164 29368 18216
rect 29420 18204 29426 18216
rect 29549 18207 29607 18213
rect 29549 18204 29561 18207
rect 29420 18176 29561 18204
rect 29420 18164 29426 18176
rect 29549 18173 29561 18176
rect 29595 18173 29607 18207
rect 29656 18204 29684 18244
rect 29805 18207 29863 18213
rect 29805 18204 29817 18207
rect 29656 18176 29817 18204
rect 29549 18167 29607 18173
rect 29805 18173 29817 18176
rect 29851 18173 29863 18207
rect 29805 18167 29863 18173
rect 29144 18108 29316 18136
rect 29144 18096 29150 18108
rect 30929 18071 30987 18077
rect 30929 18068 30941 18071
rect 28920 18040 30941 18068
rect 27157 18031 27215 18037
rect 30929 18037 30941 18040
rect 30975 18037 30987 18071
rect 30929 18031 30987 18037
rect 552 17978 31808 18000
rect 552 17926 8172 17978
rect 8224 17926 8236 17978
rect 8288 17926 8300 17978
rect 8352 17926 8364 17978
rect 8416 17926 8428 17978
rect 8480 17926 15946 17978
rect 15998 17926 16010 17978
rect 16062 17926 16074 17978
rect 16126 17926 16138 17978
rect 16190 17926 16202 17978
rect 16254 17926 23720 17978
rect 23772 17926 23784 17978
rect 23836 17926 23848 17978
rect 23900 17926 23912 17978
rect 23964 17926 23976 17978
rect 24028 17926 31494 17978
rect 31546 17926 31558 17978
rect 31610 17926 31622 17978
rect 31674 17926 31686 17978
rect 31738 17926 31750 17978
rect 31802 17926 31808 17978
rect 552 17904 31808 17926
rect 4246 17824 4252 17876
rect 4304 17864 4310 17876
rect 4304 17836 4844 17864
rect 4304 17824 4310 17836
rect 4816 17805 4844 17836
rect 4890 17824 4896 17876
rect 4948 17824 4954 17876
rect 4982 17824 4988 17876
rect 5040 17864 5046 17876
rect 5166 17864 5172 17876
rect 5040 17836 5172 17864
rect 5040 17824 5046 17836
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 5445 17867 5503 17873
rect 5445 17833 5457 17867
rect 5491 17864 5503 17867
rect 5905 17867 5963 17873
rect 5491 17836 5856 17864
rect 5491 17833 5503 17836
rect 5445 17827 5503 17833
rect 4801 17799 4859 17805
rect 4264 17768 4568 17796
rect 4264 17737 4292 17768
rect 4540 17740 4568 17768
rect 4801 17765 4813 17799
rect 4847 17765 4859 17799
rect 4801 17759 4859 17765
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17697 1639 17731
rect 1581 17691 1639 17697
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17697 4307 17731
rect 4249 17691 4307 17697
rect 1210 17484 1216 17536
rect 1268 17524 1274 17536
rect 1397 17527 1455 17533
rect 1397 17524 1409 17527
rect 1268 17496 1409 17524
rect 1268 17484 1274 17496
rect 1397 17493 1409 17496
rect 1443 17493 1455 17527
rect 1596 17524 1624 17691
rect 4338 17688 4344 17740
rect 4396 17728 4402 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4396 17700 4445 17728
rect 4396 17688 4402 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 4522 17688 4528 17740
rect 4580 17688 4586 17740
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 4908 17728 4936 17824
rect 5460 17796 5488 17827
rect 5000 17768 5488 17796
rect 5000 17740 5028 17768
rect 4755 17700 4936 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 4982 17688 4988 17740
rect 5040 17688 5046 17740
rect 5074 17688 5080 17740
rect 5132 17688 5138 17740
rect 5258 17688 5264 17740
rect 5316 17728 5322 17740
rect 5828 17737 5856 17836
rect 5905 17833 5917 17867
rect 5951 17864 5963 17867
rect 9585 17867 9643 17873
rect 5951 17836 7972 17864
rect 5951 17833 5963 17836
rect 5905 17827 5963 17833
rect 6273 17799 6331 17805
rect 6273 17765 6285 17799
rect 6319 17796 6331 17799
rect 7101 17799 7159 17805
rect 7101 17796 7113 17799
rect 6319 17768 7113 17796
rect 6319 17765 6331 17768
rect 6273 17759 6331 17765
rect 7101 17765 7113 17768
rect 7147 17765 7159 17799
rect 7101 17759 7159 17765
rect 7190 17756 7196 17808
rect 7248 17796 7254 17808
rect 7742 17805 7748 17808
rect 7248 17768 7512 17796
rect 7248 17756 7254 17768
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 5316 17700 5457 17728
rect 5316 17688 5322 17700
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 5445 17691 5503 17697
rect 5813 17731 5871 17737
rect 5813 17697 5825 17731
rect 5859 17697 5871 17731
rect 5813 17691 5871 17697
rect 5902 17688 5908 17740
rect 5960 17728 5966 17740
rect 5997 17731 6055 17737
rect 5997 17728 6009 17731
rect 5960 17700 6009 17728
rect 5960 17688 5966 17700
rect 5997 17697 6009 17700
rect 6043 17697 6055 17731
rect 5997 17691 6055 17697
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 6181 17731 6239 17737
rect 6181 17728 6193 17731
rect 6144 17700 6193 17728
rect 6144 17688 6150 17700
rect 6181 17697 6193 17700
rect 6227 17697 6239 17731
rect 6181 17691 6239 17697
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17728 6423 17731
rect 6411 17700 6960 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 5169 17663 5227 17669
rect 5169 17660 5181 17663
rect 4448 17632 5181 17660
rect 4448 17601 4476 17632
rect 5169 17629 5181 17632
rect 5215 17629 5227 17663
rect 5169 17623 5227 17629
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 6730 17620 6736 17672
rect 6788 17620 6794 17672
rect 6932 17660 6960 17700
rect 7006 17688 7012 17740
rect 7064 17728 7070 17740
rect 7374 17728 7380 17740
rect 7064 17700 7380 17728
rect 7064 17688 7070 17700
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7484 17737 7512 17768
rect 7736 17759 7748 17805
rect 7800 17796 7806 17808
rect 7800 17768 7836 17796
rect 7742 17756 7748 17759
rect 7800 17756 7806 17768
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17697 7527 17731
rect 7944 17728 7972 17836
rect 9585 17833 9597 17867
rect 9631 17864 9643 17867
rect 9766 17864 9772 17876
rect 9631 17836 9772 17864
rect 9631 17833 9643 17836
rect 9585 17827 9643 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 10134 17824 10140 17876
rect 10192 17824 10198 17876
rect 10686 17864 10692 17876
rect 10244 17836 10692 17864
rect 9309 17799 9367 17805
rect 9309 17765 9321 17799
rect 9355 17796 9367 17799
rect 10152 17796 10180 17824
rect 10244 17808 10272 17836
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 10965 17867 11023 17873
rect 10965 17833 10977 17867
rect 11011 17864 11023 17867
rect 11054 17864 11060 17876
rect 11011 17836 11060 17864
rect 11011 17833 11023 17836
rect 10965 17827 11023 17833
rect 9355 17768 10180 17796
rect 9355 17765 9367 17768
rect 9309 17759 9367 17765
rect 10226 17756 10232 17808
rect 10284 17756 10290 17808
rect 10410 17756 10416 17808
rect 10468 17756 10474 17808
rect 10980 17796 11008 17827
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 12802 17864 12808 17876
rect 12406 17836 12808 17864
rect 12406 17796 12434 17836
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 13354 17824 13360 17876
rect 13412 17824 13418 17876
rect 14737 17867 14795 17873
rect 14737 17833 14749 17867
rect 14783 17864 14795 17867
rect 14918 17864 14924 17876
rect 14783 17836 14924 17864
rect 14783 17833 14795 17836
rect 14737 17827 14795 17833
rect 14918 17824 14924 17836
rect 14976 17824 14982 17876
rect 17034 17824 17040 17876
rect 17092 17864 17098 17876
rect 17494 17864 17500 17876
rect 17092 17836 17500 17864
rect 17092 17824 17098 17836
rect 17494 17824 17500 17836
rect 17552 17864 17558 17876
rect 18598 17864 18604 17876
rect 17552 17836 18604 17864
rect 17552 17824 17558 17836
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 18785 17867 18843 17873
rect 18785 17864 18797 17867
rect 18748 17836 18797 17864
rect 18748 17824 18754 17836
rect 18785 17833 18797 17836
rect 18831 17833 18843 17867
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 18785 17827 18843 17833
rect 19306 17836 19625 17864
rect 10520 17768 11008 17796
rect 11072 17768 12434 17796
rect 12989 17799 13047 17805
rect 9125 17731 9183 17737
rect 7944 17700 8524 17728
rect 7469 17691 7527 17697
rect 7190 17660 7196 17672
rect 6932 17632 7196 17660
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7484 17660 7512 17691
rect 7285 17623 7343 17629
rect 7392 17632 7512 17660
rect 8496 17660 8524 17700
rect 9125 17697 9137 17731
rect 9171 17728 9183 17731
rect 9217 17731 9275 17737
rect 9217 17728 9229 17731
rect 9171 17700 9229 17728
rect 9171 17697 9183 17700
rect 9125 17691 9183 17697
rect 9217 17697 9229 17700
rect 9263 17697 9275 17731
rect 9217 17691 9275 17697
rect 9398 17688 9404 17740
rect 9456 17688 9462 17740
rect 9493 17731 9551 17737
rect 9493 17697 9505 17731
rect 9539 17728 9551 17731
rect 9582 17728 9588 17740
rect 9539 17700 9588 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 9689 17731 9747 17737
rect 9689 17697 9701 17731
rect 9735 17728 9747 17731
rect 9950 17728 9956 17740
rect 9735 17700 9956 17728
rect 9735 17697 9747 17700
rect 9689 17691 9747 17697
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10428 17728 10456 17756
rect 10520 17737 10548 17768
rect 10183 17700 10456 17728
rect 10505 17731 10563 17737
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 10505 17697 10517 17731
rect 10551 17697 10563 17731
rect 10505 17691 10563 17697
rect 10594 17688 10600 17740
rect 10652 17728 10658 17740
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 10652 17700 10977 17728
rect 10652 17688 10658 17700
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 10321 17663 10379 17669
rect 10321 17660 10333 17663
rect 8496 17632 10333 17660
rect 4433 17595 4491 17601
rect 4433 17561 4445 17595
rect 4479 17561 4491 17595
rect 4433 17555 4491 17561
rect 5077 17595 5135 17601
rect 5077 17561 5089 17595
rect 5123 17592 5135 17595
rect 5353 17595 5411 17601
rect 5353 17592 5365 17595
rect 5123 17564 5365 17592
rect 5123 17561 5135 17564
rect 5077 17555 5135 17561
rect 5353 17561 5365 17564
rect 5399 17592 5411 17595
rect 5442 17592 5448 17604
rect 5399 17564 5448 17592
rect 5399 17561 5411 17564
rect 5353 17555 5411 17561
rect 5442 17552 5448 17564
rect 5500 17552 5506 17604
rect 6472 17592 6500 17620
rect 6472 17564 6859 17592
rect 6831 17536 6859 17564
rect 6914 17552 6920 17604
rect 6972 17552 6978 17604
rect 7098 17552 7104 17604
rect 7156 17592 7162 17604
rect 7300 17592 7328 17623
rect 7156 17564 7328 17592
rect 7156 17552 7162 17564
rect 4525 17527 4583 17533
rect 4525 17524 4537 17527
rect 1596 17496 4537 17524
rect 1397 17487 1455 17493
rect 4525 17493 4537 17496
rect 4571 17524 4583 17527
rect 6454 17524 6460 17536
rect 4571 17496 6460 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 6638 17484 6644 17536
rect 6696 17484 6702 17536
rect 6822 17484 6828 17536
rect 6880 17484 6886 17536
rect 6932 17524 6960 17552
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 6932 17496 7205 17524
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7392 17524 7420 17632
rect 10321 17629 10333 17632
rect 10367 17629 10379 17663
rect 11072 17660 11100 17768
rect 12989 17765 13001 17799
rect 13035 17796 13047 17799
rect 13035 17768 13308 17796
rect 13035 17765 13047 17768
rect 12989 17759 13047 17765
rect 13280 17740 13308 17768
rect 11330 17728 11336 17740
rect 10321 17623 10379 17629
rect 10520 17632 11100 17660
rect 11164 17700 11336 17728
rect 8849 17595 8907 17601
rect 8849 17561 8861 17595
rect 8895 17592 8907 17595
rect 10520 17592 10548 17632
rect 8895 17564 10548 17592
rect 10597 17595 10655 17601
rect 8895 17561 8907 17564
rect 8849 17555 8907 17561
rect 10597 17561 10609 17595
rect 10643 17592 10655 17595
rect 10686 17592 10692 17604
rect 10643 17564 10692 17592
rect 10643 17561 10655 17564
rect 10597 17555 10655 17561
rect 10686 17552 10692 17564
rect 10744 17592 10750 17604
rect 11057 17595 11115 17601
rect 11057 17592 11069 17595
rect 10744 17564 11069 17592
rect 10744 17552 10750 17564
rect 11057 17561 11069 17564
rect 11103 17561 11115 17595
rect 11057 17555 11115 17561
rect 7742 17524 7748 17536
rect 7392 17496 7748 17524
rect 7193 17487 7251 17493
rect 7742 17484 7748 17496
rect 7800 17484 7806 17536
rect 9398 17484 9404 17536
rect 9456 17524 9462 17536
rect 9766 17524 9772 17536
rect 9456 17496 9772 17524
rect 9456 17484 9462 17496
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 10226 17524 10232 17536
rect 9916 17496 10232 17524
rect 9916 17484 9922 17496
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 10410 17484 10416 17536
rect 10468 17524 10474 17536
rect 11164 17524 11192 17700
rect 11330 17688 11336 17700
rect 11388 17688 11394 17740
rect 11514 17688 11520 17740
rect 11572 17688 11578 17740
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 11756 17700 12817 17728
rect 11756 17688 11762 17700
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 13081 17731 13139 17737
rect 13081 17697 13093 17731
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 11425 17663 11483 17669
rect 11425 17660 11437 17663
rect 11287 17632 11437 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11425 17629 11437 17632
rect 11471 17629 11483 17663
rect 11532 17660 11560 17688
rect 12434 17660 12440 17672
rect 11532 17632 12440 17660
rect 11425 17623 11483 17629
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 12894 17620 12900 17672
rect 12952 17660 12958 17672
rect 13096 17660 13124 17691
rect 13170 17688 13176 17740
rect 13228 17688 13234 17740
rect 13262 17688 13268 17740
rect 13320 17688 13326 17740
rect 13372 17728 13400 17824
rect 17212 17799 17270 17805
rect 15856 17768 17173 17796
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 13372 17700 13461 17728
rect 13449 17697 13461 17700
rect 13495 17697 13507 17731
rect 13449 17691 13507 17697
rect 13722 17688 13728 17740
rect 13780 17688 13786 17740
rect 15856 17737 15884 17768
rect 15841 17731 15899 17737
rect 15841 17697 15853 17731
rect 15887 17697 15899 17731
rect 15841 17691 15899 17697
rect 16945 17731 17003 17737
rect 16945 17697 16957 17731
rect 16991 17728 17003 17731
rect 17034 17728 17040 17740
rect 16991 17700 17040 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 17145 17728 17173 17768
rect 17212 17765 17224 17799
rect 17258 17796 17270 17799
rect 17586 17796 17592 17808
rect 17258 17768 17592 17796
rect 17258 17765 17270 17768
rect 17212 17759 17270 17765
rect 17586 17756 17592 17768
rect 17644 17756 17650 17808
rect 19306 17796 19334 17836
rect 19613 17833 19625 17836
rect 19659 17864 19671 17867
rect 19702 17864 19708 17876
rect 19659 17836 19708 17864
rect 19659 17833 19671 17836
rect 19613 17827 19671 17833
rect 19702 17824 19708 17836
rect 19760 17824 19766 17876
rect 22830 17824 22836 17876
rect 22888 17864 22894 17876
rect 25317 17867 25375 17873
rect 25317 17864 25329 17867
rect 22888 17836 25329 17864
rect 22888 17824 22894 17836
rect 25317 17833 25329 17836
rect 25363 17833 25375 17867
rect 26050 17864 26056 17876
rect 25317 17827 25375 17833
rect 25792 17836 26056 17864
rect 23198 17805 23204 17808
rect 19521 17799 19579 17805
rect 18156 17768 19380 17796
rect 18156 17728 18184 17768
rect 17145 17700 18184 17728
rect 18693 17731 18751 17737
rect 18693 17697 18705 17731
rect 18739 17697 18751 17731
rect 18693 17691 18751 17697
rect 12952 17632 13124 17660
rect 12952 17620 12958 17632
rect 13538 17620 13544 17672
rect 13596 17620 13602 17672
rect 13357 17595 13415 17601
rect 13357 17561 13369 17595
rect 13403 17592 13415 17595
rect 13740 17592 13768 17688
rect 14826 17620 14832 17672
rect 14884 17620 14890 17672
rect 15010 17620 15016 17672
rect 15068 17620 15074 17672
rect 18506 17620 18512 17672
rect 18564 17660 18570 17672
rect 18708 17660 18736 17691
rect 18874 17688 18880 17740
rect 18932 17688 18938 17740
rect 19242 17688 19248 17740
rect 19300 17688 19306 17740
rect 19352 17737 19380 17768
rect 19521 17765 19533 17799
rect 19567 17796 19579 17799
rect 20073 17799 20131 17805
rect 20073 17796 20085 17799
rect 19567 17768 20085 17796
rect 19567 17765 19579 17768
rect 19521 17759 19579 17765
rect 20073 17765 20085 17768
rect 20119 17765 20131 17799
rect 23192 17796 23204 17805
rect 20073 17759 20131 17765
rect 20180 17768 20576 17796
rect 23159 17768 23204 17796
rect 19337 17731 19395 17737
rect 19337 17697 19349 17731
rect 19383 17697 19395 17731
rect 19337 17691 19395 17697
rect 19610 17688 19616 17740
rect 19668 17688 19674 17740
rect 20180 17737 20208 17768
rect 19981 17731 20039 17737
rect 19981 17728 19993 17731
rect 19812 17700 19993 17728
rect 18564 17632 18736 17660
rect 19260 17660 19288 17688
rect 19628 17660 19656 17688
rect 19260 17632 19656 17660
rect 18564 17620 18570 17632
rect 13403 17564 13768 17592
rect 13403 17561 13415 17564
rect 13357 17555 13415 17561
rect 15102 17552 15108 17604
rect 15160 17592 15166 17604
rect 19518 17592 19524 17604
rect 15160 17564 15792 17592
rect 15160 17552 15166 17564
rect 10468 17496 11192 17524
rect 10468 17484 10474 17496
rect 13446 17484 13452 17536
rect 13504 17484 13510 17536
rect 13814 17484 13820 17536
rect 13872 17484 13878 17536
rect 14366 17484 14372 17536
rect 14424 17484 14430 17536
rect 15654 17484 15660 17536
rect 15712 17484 15718 17536
rect 15764 17524 15792 17564
rect 17880 17564 19524 17592
rect 17880 17524 17908 17564
rect 19518 17552 19524 17564
rect 19576 17552 19582 17604
rect 19705 17595 19763 17601
rect 19705 17561 19717 17595
rect 19751 17561 19763 17595
rect 19812 17592 19840 17700
rect 19981 17697 19993 17700
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 20165 17731 20223 17737
rect 20165 17697 20177 17731
rect 20211 17697 20223 17731
rect 20165 17691 20223 17697
rect 20254 17688 20260 17740
rect 20312 17688 20318 17740
rect 20548 17737 20576 17768
rect 23192 17759 23204 17768
rect 23198 17756 23204 17759
rect 23256 17756 23262 17808
rect 24673 17799 24731 17805
rect 24673 17765 24685 17799
rect 24719 17796 24731 17799
rect 24854 17796 24860 17808
rect 24719 17768 24860 17796
rect 24719 17765 24731 17768
rect 24673 17759 24731 17765
rect 24854 17756 24860 17768
rect 24912 17756 24918 17808
rect 20441 17731 20499 17737
rect 20441 17697 20453 17731
rect 20487 17697 20499 17731
rect 20441 17691 20499 17697
rect 20533 17731 20591 17737
rect 20533 17697 20545 17731
rect 20579 17697 20591 17731
rect 20533 17691 20591 17697
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 19935 17632 20361 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 20349 17629 20361 17632
rect 20395 17629 20407 17663
rect 20456 17660 20484 17691
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20772 17700 20913 17728
rect 20772 17688 20778 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 22922 17688 22928 17740
rect 22980 17688 22986 17740
rect 25792 17737 25820 17836
rect 26050 17824 26056 17836
rect 26108 17864 26114 17876
rect 26697 17867 26755 17873
rect 26697 17864 26709 17867
rect 26108 17836 26709 17864
rect 26108 17824 26114 17836
rect 26697 17833 26709 17836
rect 26743 17833 26755 17867
rect 26697 17827 26755 17833
rect 26786 17824 26792 17876
rect 26844 17864 26850 17876
rect 27341 17867 27399 17873
rect 27341 17864 27353 17867
rect 26844 17836 27353 17864
rect 26844 17824 26850 17836
rect 27341 17833 27353 17836
rect 27387 17833 27399 17867
rect 27341 17827 27399 17833
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 29089 17867 29147 17873
rect 29089 17864 29101 17867
rect 29052 17836 29101 17864
rect 29052 17824 29058 17836
rect 29089 17833 29101 17836
rect 29135 17833 29147 17867
rect 29089 17827 29147 17833
rect 29454 17824 29460 17876
rect 29512 17824 29518 17876
rect 25866 17756 25872 17808
rect 25924 17796 25930 17808
rect 29914 17805 29920 17808
rect 27157 17799 27215 17805
rect 27157 17796 27169 17799
rect 25924 17768 27169 17796
rect 25924 17756 25930 17768
rect 27157 17765 27169 17768
rect 27203 17796 27215 17799
rect 27617 17799 27675 17805
rect 27617 17796 27629 17799
rect 27203 17768 27629 17796
rect 27203 17765 27215 17768
rect 27157 17759 27215 17765
rect 27617 17765 27629 17768
rect 27663 17765 27675 17799
rect 27617 17759 27675 17765
rect 28077 17799 28135 17805
rect 28077 17765 28089 17799
rect 28123 17765 28135 17799
rect 29908 17796 29920 17805
rect 28077 17759 28135 17765
rect 29104 17768 29408 17796
rect 29875 17768 29920 17796
rect 24765 17731 24823 17737
rect 24765 17697 24777 17731
rect 24811 17728 24823 17731
rect 25777 17731 25835 17737
rect 25777 17728 25789 17731
rect 24811 17700 25789 17728
rect 24811 17697 24823 17700
rect 24765 17691 24823 17697
rect 25777 17697 25789 17700
rect 25823 17728 25835 17731
rect 28092 17728 28120 17759
rect 29104 17740 29132 17768
rect 25823 17700 28120 17728
rect 25823 17697 25835 17700
rect 25777 17691 25835 17697
rect 28994 17688 29000 17740
rect 29052 17688 29058 17740
rect 29086 17688 29092 17740
rect 29144 17688 29150 17740
rect 29181 17731 29239 17737
rect 29181 17697 29193 17731
rect 29227 17697 29239 17731
rect 29181 17691 29239 17697
rect 20732 17660 20760 17688
rect 24556 17663 24614 17669
rect 24556 17660 24568 17663
rect 20456 17632 20760 17660
rect 24320 17632 24568 17660
rect 20349 17623 20407 17629
rect 20254 17592 20260 17604
rect 19812 17564 20260 17592
rect 19705 17555 19763 17561
rect 15764 17496 17908 17524
rect 18322 17484 18328 17536
rect 18380 17484 18386 17536
rect 18506 17484 18512 17536
rect 18564 17524 18570 17536
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 18564 17496 19257 17524
rect 18564 17484 18570 17496
rect 19245 17493 19257 17496
rect 19291 17524 19303 17527
rect 19720 17524 19748 17555
rect 20254 17552 20260 17564
rect 20312 17592 20318 17604
rect 20438 17592 20444 17604
rect 20312 17564 20444 17592
rect 20312 17552 20318 17564
rect 20438 17552 20444 17564
rect 20496 17552 20502 17604
rect 24320 17601 24348 17632
rect 24556 17629 24568 17632
rect 24602 17629 24614 17663
rect 24556 17623 24614 17629
rect 24946 17620 24952 17672
rect 25004 17660 25010 17672
rect 25041 17663 25099 17669
rect 25041 17660 25053 17663
rect 25004 17632 25053 17660
rect 25004 17620 25010 17632
rect 25041 17629 25053 17632
rect 25087 17629 25099 17663
rect 25041 17623 25099 17629
rect 26602 17620 26608 17672
rect 26660 17620 26666 17672
rect 27522 17620 27528 17672
rect 27580 17620 27586 17672
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 29196 17660 29224 17691
rect 29270 17688 29276 17740
rect 29328 17688 29334 17740
rect 29380 17737 29408 17768
rect 29908 17759 29920 17768
rect 29914 17756 29920 17759
rect 29972 17756 29978 17808
rect 29365 17731 29423 17737
rect 29365 17697 29377 17731
rect 29411 17697 29423 17731
rect 29365 17691 29423 17697
rect 29546 17688 29552 17740
rect 29604 17688 29610 17740
rect 28868 17632 29224 17660
rect 29288 17660 29316 17688
rect 29641 17663 29699 17669
rect 29641 17660 29653 17663
rect 29288 17632 29653 17660
rect 28868 17620 28874 17632
rect 24305 17595 24363 17601
rect 24305 17561 24317 17595
rect 24351 17561 24363 17595
rect 24305 17555 24363 17561
rect 24854 17552 24860 17604
rect 24912 17592 24918 17604
rect 26421 17595 26479 17601
rect 26421 17592 26433 17595
rect 24912 17564 26433 17592
rect 24912 17552 24918 17564
rect 26421 17561 26433 17564
rect 26467 17561 26479 17595
rect 26421 17555 26479 17561
rect 27157 17595 27215 17601
rect 27157 17561 27169 17595
rect 27203 17592 27215 17595
rect 27982 17592 27988 17604
rect 27203 17564 27988 17592
rect 27203 17561 27215 17564
rect 27157 17555 27215 17561
rect 27982 17552 27988 17564
rect 28040 17592 28046 17604
rect 28077 17595 28135 17601
rect 28077 17592 28089 17595
rect 28040 17564 28089 17592
rect 28040 17552 28046 17564
rect 28077 17561 28089 17564
rect 28123 17561 28135 17595
rect 29196 17592 29224 17632
rect 29641 17629 29653 17632
rect 29687 17629 29699 17663
rect 29641 17623 29699 17629
rect 29454 17592 29460 17604
rect 29196 17564 29460 17592
rect 28077 17555 28135 17561
rect 29454 17552 29460 17564
rect 29512 17552 29518 17604
rect 19291 17496 19748 17524
rect 19291 17493 19303 17496
rect 19245 17487 19303 17493
rect 21082 17484 21088 17536
rect 21140 17484 21146 17536
rect 22646 17484 22652 17536
rect 22704 17524 22710 17536
rect 23566 17524 23572 17536
rect 22704 17496 23572 17524
rect 22704 17484 22710 17496
rect 23566 17484 23572 17496
rect 23624 17484 23630 17536
rect 24394 17484 24400 17536
rect 24452 17484 24458 17536
rect 25685 17527 25743 17533
rect 25685 17493 25697 17527
rect 25731 17524 25743 17527
rect 26142 17524 26148 17536
rect 25731 17496 26148 17524
rect 25731 17493 25743 17496
rect 25685 17487 25743 17493
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 26326 17484 26332 17536
rect 26384 17524 26390 17536
rect 28166 17524 28172 17536
rect 26384 17496 28172 17524
rect 26384 17484 26390 17496
rect 28166 17484 28172 17496
rect 28224 17484 28230 17536
rect 31018 17484 31024 17536
rect 31076 17484 31082 17536
rect 552 17434 31648 17456
rect 552 17382 4285 17434
rect 4337 17382 4349 17434
rect 4401 17382 4413 17434
rect 4465 17382 4477 17434
rect 4529 17382 4541 17434
rect 4593 17382 12059 17434
rect 12111 17382 12123 17434
rect 12175 17382 12187 17434
rect 12239 17382 12251 17434
rect 12303 17382 12315 17434
rect 12367 17382 19833 17434
rect 19885 17382 19897 17434
rect 19949 17382 19961 17434
rect 20013 17382 20025 17434
rect 20077 17382 20089 17434
rect 20141 17382 27607 17434
rect 27659 17382 27671 17434
rect 27723 17382 27735 17434
rect 27787 17382 27799 17434
rect 27851 17382 27863 17434
rect 27915 17382 31648 17434
rect 552 17360 31648 17382
rect 5092 17292 6592 17320
rect 4617 17255 4675 17261
rect 4617 17221 4629 17255
rect 4663 17252 4675 17255
rect 5092 17252 5120 17292
rect 4663 17224 5120 17252
rect 6564 17252 6592 17292
rect 6730 17280 6736 17332
rect 6788 17320 6794 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6788 17292 6837 17320
rect 6788 17280 6794 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 9582 17320 9588 17332
rect 6825 17283 6883 17289
rect 8404 17292 9588 17320
rect 8404 17252 8432 17292
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10137 17323 10195 17329
rect 10137 17320 10149 17323
rect 9824 17292 10149 17320
rect 9824 17280 9830 17292
rect 10137 17289 10149 17292
rect 10183 17320 10195 17323
rect 10183 17292 10456 17320
rect 10183 17289 10195 17292
rect 10137 17283 10195 17289
rect 10428 17264 10456 17292
rect 10502 17280 10508 17332
rect 10560 17280 10566 17332
rect 10686 17280 10692 17332
rect 10744 17280 10750 17332
rect 13265 17323 13323 17329
rect 13265 17289 13277 17323
rect 13311 17320 13323 17323
rect 13446 17320 13452 17332
rect 13311 17292 13452 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13814 17280 13820 17332
rect 13872 17280 13878 17332
rect 14366 17280 14372 17332
rect 14424 17280 14430 17332
rect 14734 17280 14740 17332
rect 14792 17280 14798 17332
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14884 17292 15117 17320
rect 14884 17280 14890 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 15105 17283 15163 17289
rect 18138 17280 18144 17332
rect 18196 17280 18202 17332
rect 19518 17320 19524 17332
rect 19306 17292 19524 17320
rect 6564 17224 8432 17252
rect 4663 17221 4675 17224
rect 4617 17215 4675 17221
rect 9950 17212 9956 17264
rect 10008 17252 10014 17264
rect 10045 17255 10103 17261
rect 10045 17252 10057 17255
rect 10008 17224 10057 17252
rect 10008 17212 10014 17224
rect 10045 17221 10057 17224
rect 10091 17252 10103 17255
rect 10321 17255 10379 17261
rect 10321 17252 10333 17255
rect 10091 17224 10333 17252
rect 10091 17221 10103 17224
rect 10045 17215 10103 17221
rect 10321 17221 10333 17224
rect 10367 17221 10379 17255
rect 10321 17215 10379 17221
rect 10410 17212 10416 17264
rect 10468 17212 10474 17264
rect 10520 17252 10548 17280
rect 10520 17224 10640 17252
rect 5074 17184 5080 17196
rect 4724 17156 5080 17184
rect 1210 17076 1216 17128
rect 1268 17076 1274 17128
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17116 3295 17119
rect 3326 17116 3332 17128
rect 3283 17088 3332 17116
rect 3283 17085 3295 17088
rect 3237 17079 3295 17085
rect 3326 17076 3332 17088
rect 3384 17116 3390 17128
rect 4724 17116 4752 17156
rect 5074 17144 5080 17156
rect 5132 17144 5138 17196
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6696 17156 6868 17184
rect 6696 17144 6702 17156
rect 3384 17088 4752 17116
rect 4801 17119 4859 17125
rect 3384 17076 3390 17088
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 4982 17116 4988 17128
rect 4847 17088 4988 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 6840 17125 6868 17156
rect 7024 17156 7604 17184
rect 7024 17128 7052 17156
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7006 17076 7012 17128
rect 7064 17076 7070 17128
rect 7098 17076 7104 17128
rect 7156 17116 7162 17128
rect 7576 17125 7604 17156
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 10502 17184 10508 17196
rect 7708 17156 8524 17184
rect 7708 17144 7714 17156
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 7156 17088 7297 17116
rect 7156 17076 7162 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 7561 17119 7619 17125
rect 7561 17085 7573 17119
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 7742 17076 7748 17128
rect 7800 17116 7806 17128
rect 8389 17119 8447 17125
rect 8389 17116 8401 17119
rect 7800 17088 8401 17116
rect 7800 17076 7806 17088
rect 8389 17085 8401 17088
rect 8435 17085 8447 17119
rect 8496 17116 8524 17156
rect 9876 17156 10508 17184
rect 9876 17116 9904 17156
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 10612 17193 10640 17224
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 8496 17088 9904 17116
rect 9953 17119 10011 17125
rect 8389 17079 8447 17085
rect 9953 17085 9965 17119
rect 9999 17116 10011 17119
rect 10042 17116 10048 17128
rect 9999 17088 10048 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 10042 17076 10048 17088
rect 10100 17116 10106 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 10100 17088 10333 17116
rect 10100 17076 10106 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10321 17079 10379 17085
rect 10410 17076 10416 17128
rect 10468 17076 10474 17128
rect 10704 17125 10732 17280
rect 12345 17255 12403 17261
rect 12345 17221 12357 17255
rect 12391 17252 12403 17255
rect 13722 17252 13728 17264
rect 12391 17224 13728 17252
rect 12391 17221 12403 17224
rect 12345 17215 12403 17221
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 10796 17156 11100 17184
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 1486 17008 1492 17060
rect 1544 17008 1550 17060
rect 2222 17008 2228 17060
rect 2280 17008 2286 17060
rect 3482 17051 3540 17057
rect 3482 17048 3494 17051
rect 2976 17020 3494 17048
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 2976 16989 3004 17020
rect 3482 17017 3494 17020
rect 3528 17017 3540 17051
rect 5322 17051 5380 17057
rect 5322 17048 5334 17051
rect 3482 17011 3540 17017
rect 5000 17020 5334 17048
rect 5000 16989 5028 17020
rect 5322 17017 5334 17020
rect 5368 17017 5380 17051
rect 7650 17048 7656 17060
rect 5322 17011 5380 17017
rect 6472 17020 7656 17048
rect 6472 16989 6500 17020
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 8634 17051 8692 17057
rect 8634 17048 8646 17051
rect 7760 17020 8646 17048
rect 2961 16983 3019 16989
rect 2961 16980 2973 16983
rect 1452 16952 2973 16980
rect 1452 16940 1458 16952
rect 2961 16949 2973 16952
rect 3007 16949 3019 16983
rect 2961 16943 3019 16949
rect 4985 16983 5043 16989
rect 4985 16949 4997 16983
rect 5031 16949 5043 16983
rect 4985 16943 5043 16949
rect 6457 16983 6515 16989
rect 6457 16949 6469 16983
rect 6503 16949 6515 16983
rect 6457 16943 6515 16949
rect 7098 16940 7104 16992
rect 7156 16940 7162 16992
rect 7760 16989 7788 17020
rect 8634 17017 8646 17020
rect 8680 17017 8692 17051
rect 10229 17051 10287 17057
rect 8634 17011 8692 17017
rect 9784 17020 10180 17048
rect 9784 16989 9812 17020
rect 7745 16983 7803 16989
rect 7745 16949 7757 16983
rect 7791 16949 7803 16983
rect 7745 16943 7803 16949
rect 9769 16983 9827 16989
rect 9769 16949 9781 16983
rect 9815 16949 9827 16983
rect 10152 16980 10180 17020
rect 10229 17017 10241 17051
rect 10275 17048 10287 17051
rect 10594 17048 10600 17060
rect 10275 17020 10600 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 10594 17008 10600 17020
rect 10652 17008 10658 17060
rect 10796 16980 10824 17156
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10928 17088 10977 17116
rect 10928 17076 10934 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 11072 17116 11100 17156
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 12032 17156 13032 17184
rect 12032 17144 12038 17156
rect 13004 17125 13032 17156
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 11072 17088 12725 17116
rect 10965 17079 11023 17085
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17085 13047 17119
rect 12989 17079 13047 17085
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13170 17116 13176 17128
rect 13127 17088 13176 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 13170 17076 13176 17088
rect 13228 17116 13234 17128
rect 13832 17125 13860 17280
rect 14384 17125 14412 17280
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 16540 17224 17632 17252
rect 16540 17212 16546 17224
rect 14550 17144 14556 17196
rect 14608 17144 14614 17196
rect 16574 17144 16580 17196
rect 16632 17144 16638 17196
rect 17310 17144 17316 17196
rect 17368 17144 17374 17196
rect 13817 17119 13875 17125
rect 13228 17088 13771 17116
rect 13228 17076 13234 17088
rect 11210 17051 11268 17057
rect 11210 17048 11222 17051
rect 10888 17020 11222 17048
rect 10888 16989 10916 17020
rect 11210 17017 11222 17020
rect 11256 17017 11268 17051
rect 11210 17011 11268 17017
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 12897 17051 12955 17057
rect 12897 17048 12909 17051
rect 12584 17020 12909 17048
rect 12584 17008 12590 17020
rect 12897 17017 12909 17020
rect 12943 17048 12955 17051
rect 12943 17020 13676 17048
rect 12943 17017 12955 17020
rect 12897 17011 12955 17017
rect 13648 16992 13676 17020
rect 10152 16952 10824 16980
rect 10873 16983 10931 16989
rect 9769 16943 9827 16949
rect 10873 16949 10885 16983
rect 10919 16949 10931 16983
rect 10873 16943 10931 16949
rect 13630 16940 13636 16992
rect 13688 16940 13694 16992
rect 13743 16980 13771 17088
rect 13817 17085 13829 17119
rect 13863 17085 13875 17119
rect 13817 17079 13875 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17085 14427 17119
rect 14369 17079 14427 17085
rect 14016 17048 14044 17079
rect 15654 17076 15660 17128
rect 15712 17116 15718 17128
rect 16218 17119 16276 17125
rect 16218 17116 16230 17119
rect 15712 17088 16230 17116
rect 15712 17076 15718 17088
rect 16218 17085 16230 17088
rect 16264 17085 16276 17119
rect 16218 17079 16276 17085
rect 16390 17076 16396 17128
rect 16448 17116 16454 17128
rect 16485 17119 16543 17125
rect 16485 17116 16497 17119
rect 16448 17088 16497 17116
rect 16448 17076 16454 17088
rect 16485 17085 16497 17088
rect 16531 17085 16543 17119
rect 16485 17079 16543 17085
rect 17126 17076 17132 17128
rect 17184 17116 17190 17128
rect 17604 17125 17632 17224
rect 18230 17212 18236 17264
rect 18288 17252 18294 17264
rect 19306 17252 19334 17292
rect 19518 17280 19524 17292
rect 19576 17280 19582 17332
rect 23198 17320 23204 17332
rect 19904 17292 23204 17320
rect 18288 17224 19334 17252
rect 18288 17212 18294 17224
rect 17678 17144 17684 17196
rect 17736 17184 17742 17196
rect 17736 17156 18276 17184
rect 17736 17144 17742 17156
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 17184 17088 17233 17116
rect 17184 17076 17190 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17085 17647 17119
rect 17589 17079 17647 17085
rect 17773 17119 17831 17125
rect 17773 17085 17785 17119
rect 17819 17116 17831 17119
rect 17819 17088 18000 17116
rect 17819 17085 17831 17088
rect 17773 17079 17831 17085
rect 17972 17048 18000 17088
rect 18046 17076 18052 17128
rect 18104 17076 18110 17128
rect 18248 17125 18276 17156
rect 18233 17119 18291 17125
rect 18233 17085 18245 17119
rect 18279 17085 18291 17119
rect 18233 17079 18291 17085
rect 18506 17076 18512 17128
rect 18564 17076 18570 17128
rect 18874 17076 18880 17128
rect 18932 17076 18938 17128
rect 18984 17116 19012 17224
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 18984 17088 19073 17116
rect 19061 17085 19073 17088
rect 19107 17085 19119 17119
rect 19061 17079 19119 17085
rect 19242 17076 19248 17128
rect 19300 17076 19306 17128
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 19521 17119 19579 17125
rect 19521 17116 19533 17119
rect 19484 17088 19533 17116
rect 19484 17076 19490 17088
rect 19521 17085 19533 17088
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 14016 17020 17908 17048
rect 17972 17020 18920 17048
rect 16298 16980 16304 16992
rect 13743 16952 16304 16980
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 17880 16989 17908 17020
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16949 17923 16983
rect 17865 16943 17923 16949
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18325 16983 18383 16989
rect 18325 16980 18337 16983
rect 18012 16952 18337 16980
rect 18012 16940 18018 16952
rect 18325 16949 18337 16952
rect 18371 16949 18383 16983
rect 18325 16943 18383 16949
rect 18690 16940 18696 16992
rect 18748 16940 18754 16992
rect 18892 16980 18920 17020
rect 18966 17008 18972 17060
rect 19024 17008 19030 17060
rect 19904 17048 19932 17292
rect 23198 17280 23204 17292
rect 23256 17280 23262 17332
rect 24486 17280 24492 17332
rect 24544 17280 24550 17332
rect 26602 17280 26608 17332
rect 26660 17320 26666 17332
rect 27433 17323 27491 17329
rect 27433 17320 27445 17323
rect 26660 17292 27445 17320
rect 26660 17280 26666 17292
rect 27433 17289 27445 17292
rect 27479 17289 27491 17323
rect 27433 17283 27491 17289
rect 29457 17323 29515 17329
rect 29457 17289 29469 17323
rect 29503 17320 29515 17323
rect 29546 17320 29552 17332
rect 29503 17292 29552 17320
rect 29503 17289 29515 17292
rect 29457 17283 29515 17289
rect 29546 17280 29552 17292
rect 29604 17280 29610 17332
rect 20254 17212 20260 17264
rect 20312 17212 20318 17264
rect 24305 17255 24363 17261
rect 24305 17221 24317 17255
rect 24351 17252 24363 17255
rect 24670 17252 24676 17264
rect 24351 17224 24676 17252
rect 24351 17221 24363 17224
rect 24305 17215 24363 17221
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 26694 17252 26700 17264
rect 25884 17224 26700 17252
rect 20272 17184 20300 17212
rect 25884 17184 25912 17224
rect 26694 17212 26700 17224
rect 26752 17212 26758 17264
rect 19996 17156 20300 17184
rect 24228 17156 25912 17184
rect 26053 17187 26111 17193
rect 19996 17125 20024 17156
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 20257 17119 20315 17125
rect 20257 17085 20269 17119
rect 20303 17116 20315 17119
rect 20346 17116 20352 17128
rect 20303 17088 20352 17116
rect 20303 17085 20315 17088
rect 20257 17079 20315 17085
rect 20346 17076 20352 17088
rect 20404 17116 20410 17128
rect 20990 17116 20996 17128
rect 20404 17088 20996 17116
rect 20404 17076 20410 17088
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 21082 17076 21088 17128
rect 21140 17076 21146 17128
rect 21729 17119 21787 17125
rect 21729 17085 21741 17119
rect 21775 17116 21787 17119
rect 22278 17116 22284 17128
rect 21775 17088 22284 17116
rect 21775 17085 21787 17088
rect 21729 17079 21787 17085
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 24228 17116 24256 17156
rect 26053 17153 26065 17187
rect 26099 17184 26111 17187
rect 27065 17187 27123 17193
rect 26099 17156 27016 17184
rect 26099 17153 26111 17156
rect 26053 17147 26111 17153
rect 26068 17116 26096 17147
rect 22612 17088 24256 17116
rect 24320 17088 26096 17116
rect 22612 17076 22618 17088
rect 20502 17051 20560 17057
rect 20502 17048 20514 17051
rect 19067 17020 19932 17048
rect 20180 17020 20514 17048
rect 19067 16980 19095 17020
rect 18892 16952 19095 16980
rect 19334 16940 19340 16992
rect 19392 16940 19398 16992
rect 20180 16989 20208 17020
rect 20502 17017 20514 17020
rect 20548 17017 20560 17051
rect 21100 17048 21128 17076
rect 21974 17051 22032 17057
rect 21974 17048 21986 17051
rect 21100 17020 21986 17048
rect 20502 17011 20560 17017
rect 21974 17017 21986 17020
rect 22020 17017 22032 17051
rect 21974 17011 22032 17017
rect 22094 17008 22100 17060
rect 22152 17048 22158 17060
rect 24320 17048 24348 17088
rect 26326 17076 26332 17128
rect 26384 17076 26390 17128
rect 26418 17076 26424 17128
rect 26476 17116 26482 17128
rect 26988 17125 27016 17156
rect 27065 17153 27077 17187
rect 27111 17184 27123 17187
rect 27798 17184 27804 17196
rect 27111 17156 27804 17184
rect 27111 17153 27123 17156
rect 27065 17147 27123 17153
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 30374 17184 30380 17196
rect 28736 17156 30380 17184
rect 26789 17119 26847 17125
rect 26789 17116 26801 17119
rect 26476 17088 26801 17116
rect 26476 17076 26482 17088
rect 26789 17085 26801 17088
rect 26835 17085 26847 17119
rect 26789 17079 26847 17085
rect 26973 17119 27031 17125
rect 26973 17085 26985 17119
rect 27019 17085 27031 17119
rect 28736 17116 28764 17156
rect 30374 17144 30380 17156
rect 30432 17144 30438 17196
rect 26973 17079 27031 17085
rect 27172 17088 28764 17116
rect 28813 17119 28871 17125
rect 22152 17020 24348 17048
rect 22152 17008 22158 17020
rect 24762 17008 24768 17060
rect 24820 17048 24826 17060
rect 24857 17051 24915 17057
rect 24857 17048 24869 17051
rect 24820 17020 24869 17048
rect 24820 17008 24826 17020
rect 24857 17017 24869 17020
rect 24903 17017 24915 17051
rect 27172 17048 27200 17088
rect 28813 17085 28825 17119
rect 28859 17085 28871 17119
rect 28813 17079 28871 17085
rect 24857 17011 24915 17017
rect 26804 17020 27200 17048
rect 27249 17051 27307 17057
rect 20165 16983 20223 16989
rect 20165 16949 20177 16983
rect 20211 16949 20223 16983
rect 20165 16943 20223 16949
rect 21634 16940 21640 16992
rect 21692 16940 21698 16992
rect 22462 16940 22468 16992
rect 22520 16980 22526 16992
rect 22922 16980 22928 16992
rect 22520 16952 22928 16980
rect 22520 16940 22526 16952
rect 22922 16940 22928 16952
rect 22980 16940 22986 16992
rect 23106 16940 23112 16992
rect 23164 16940 23170 16992
rect 24480 16983 24538 16989
rect 24480 16949 24492 16983
rect 24526 16980 24538 16983
rect 24946 16980 24952 16992
rect 24526 16952 24952 16980
rect 24526 16949 24538 16952
rect 24480 16943 24538 16949
rect 24946 16940 24952 16952
rect 25004 16940 25010 16992
rect 25314 16940 25320 16992
rect 25372 16980 25378 16992
rect 26804 16980 26832 17020
rect 27249 17017 27261 17051
rect 27295 17048 27307 17051
rect 27982 17048 27988 17060
rect 27295 17020 27988 17048
rect 27295 17017 27307 17020
rect 27249 17011 27307 17017
rect 27982 17008 27988 17020
rect 28040 17008 28046 17060
rect 28074 17008 28080 17060
rect 28132 17048 28138 17060
rect 28546 17051 28604 17057
rect 28546 17048 28558 17051
rect 28132 17020 28558 17048
rect 28132 17008 28138 17020
rect 28546 17017 28558 17020
rect 28592 17017 28604 17051
rect 28828 17048 28856 17079
rect 28902 17076 28908 17128
rect 28960 17116 28966 17128
rect 28997 17119 29055 17125
rect 28997 17116 29009 17119
rect 28960 17088 29009 17116
rect 28960 17076 28966 17088
rect 28997 17085 29009 17088
rect 29043 17085 29055 17119
rect 28997 17079 29055 17085
rect 29086 17076 29092 17128
rect 29144 17116 29150 17128
rect 29733 17119 29791 17125
rect 29733 17116 29745 17119
rect 29144 17088 29745 17116
rect 29144 17076 29150 17088
rect 29733 17085 29745 17088
rect 29779 17085 29791 17119
rect 29733 17079 29791 17085
rect 29178 17048 29184 17060
rect 28828 17020 29184 17048
rect 28546 17011 28604 17017
rect 29178 17008 29184 17020
rect 29236 17008 29242 17060
rect 29270 17008 29276 17060
rect 29328 17008 29334 17060
rect 25372 16952 26832 16980
rect 25372 16940 25378 16952
rect 26878 16940 26884 16992
rect 26936 16940 26942 16992
rect 28994 16940 29000 16992
rect 29052 16940 29058 16992
rect 29196 16980 29224 17008
rect 29822 16980 29828 16992
rect 29196 16952 29828 16980
rect 29822 16940 29828 16952
rect 29880 16940 29886 16992
rect 29914 16940 29920 16992
rect 29972 16940 29978 16992
rect 552 16890 31808 16912
rect 552 16838 8172 16890
rect 8224 16838 8236 16890
rect 8288 16838 8300 16890
rect 8352 16838 8364 16890
rect 8416 16838 8428 16890
rect 8480 16838 15946 16890
rect 15998 16838 16010 16890
rect 16062 16838 16074 16890
rect 16126 16838 16138 16890
rect 16190 16838 16202 16890
rect 16254 16838 23720 16890
rect 23772 16838 23784 16890
rect 23836 16838 23848 16890
rect 23900 16838 23912 16890
rect 23964 16838 23976 16890
rect 24028 16838 31494 16890
rect 31546 16838 31558 16890
rect 31610 16838 31622 16890
rect 31674 16838 31686 16890
rect 31738 16838 31750 16890
rect 31802 16838 31808 16890
rect 552 16816 31808 16838
rect 1486 16736 1492 16788
rect 1544 16736 1550 16788
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 2317 16779 2375 16785
rect 2317 16776 2329 16779
rect 2280 16748 2329 16776
rect 2280 16736 2286 16748
rect 2317 16745 2329 16748
rect 2363 16745 2375 16779
rect 2317 16739 2375 16745
rect 4893 16779 4951 16785
rect 4893 16745 4905 16779
rect 4939 16745 4951 16779
rect 4893 16739 4951 16745
rect 1504 16708 1532 16736
rect 4798 16708 4804 16720
rect 1504 16680 1624 16708
rect 1213 16643 1271 16649
rect 1213 16609 1225 16643
rect 1259 16640 1271 16643
rect 1394 16640 1400 16652
rect 1259 16612 1400 16640
rect 1259 16609 1271 16612
rect 1213 16603 1271 16609
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1302 16532 1308 16584
rect 1360 16532 1366 16584
rect 1596 16581 1624 16680
rect 2700 16680 4804 16708
rect 2406 16600 2412 16652
rect 2464 16600 2470 16652
rect 2700 16649 2728 16680
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 4908 16708 4936 16739
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7193 16779 7251 16785
rect 7193 16776 7205 16779
rect 7064 16748 7205 16776
rect 7064 16736 7070 16748
rect 7193 16745 7205 16748
rect 7239 16776 7251 16779
rect 7650 16776 7656 16788
rect 7239 16748 7656 16776
rect 7239 16745 7251 16748
rect 7193 16739 7251 16745
rect 7650 16736 7656 16748
rect 7708 16736 7714 16788
rect 9950 16736 9956 16788
rect 10008 16736 10014 16788
rect 10321 16779 10379 16785
rect 10321 16745 10333 16779
rect 10367 16745 10379 16779
rect 10321 16739 10379 16745
rect 10505 16779 10563 16785
rect 10505 16745 10517 16779
rect 10551 16776 10563 16779
rect 10594 16776 10600 16788
rect 10551 16748 10600 16776
rect 10551 16745 10563 16748
rect 10505 16739 10563 16745
rect 4908 16680 9720 16708
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 3326 16600 3332 16652
rect 3384 16640 3390 16652
rect 3786 16649 3792 16652
rect 3513 16643 3571 16649
rect 3513 16640 3525 16643
rect 3384 16612 3525 16640
rect 3384 16600 3390 16612
rect 3513 16609 3525 16612
rect 3559 16609 3571 16643
rect 3780 16640 3792 16649
rect 3747 16612 3792 16640
rect 3513 16603 3571 16609
rect 3780 16603 3792 16612
rect 3786 16600 3792 16603
rect 3844 16600 3850 16652
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 7374 16640 7380 16652
rect 7239 16612 7380 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 7374 16600 7380 16612
rect 7432 16640 7438 16652
rect 7561 16643 7619 16649
rect 7561 16640 7573 16643
rect 7432 16612 7573 16640
rect 7432 16600 7438 16612
rect 7561 16609 7573 16612
rect 7607 16609 7619 16643
rect 7561 16603 7619 16609
rect 7650 16600 7656 16652
rect 7708 16600 7714 16652
rect 9692 16640 9720 16680
rect 9968 16640 9996 16736
rect 10336 16652 10364 16739
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 10686 16736 10692 16788
rect 10744 16736 10750 16788
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 13909 16779 13967 16785
rect 13909 16776 13921 16779
rect 13596 16748 13921 16776
rect 13596 16736 13602 16748
rect 13909 16745 13921 16748
rect 13955 16745 13967 16779
rect 13909 16739 13967 16745
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 14829 16779 14887 16785
rect 14829 16776 14841 16779
rect 14056 16748 14841 16776
rect 14056 16736 14062 16748
rect 14829 16745 14841 16748
rect 14875 16776 14887 16779
rect 15933 16779 15991 16785
rect 14875 16748 15332 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 10704 16708 10732 16736
rect 10428 16680 10732 16708
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9692 16612 9904 16640
rect 9968 16612 10149 16640
rect 1581 16575 1639 16581
rect 1581 16541 1593 16575
rect 1627 16541 1639 16575
rect 1581 16535 1639 16541
rect 7466 16532 7472 16584
rect 7524 16532 7530 16584
rect 7834 16532 7840 16584
rect 7892 16532 7898 16584
rect 7285 16507 7343 16513
rect 7285 16473 7297 16507
rect 7331 16504 7343 16507
rect 7558 16504 7564 16516
rect 7331 16476 7564 16504
rect 7331 16473 7343 16476
rect 7285 16467 7343 16473
rect 7558 16464 7564 16476
rect 7616 16464 7622 16516
rect 9876 16504 9904 16612
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 10318 16600 10324 16652
rect 10376 16600 10382 16652
rect 10428 16649 10456 16680
rect 10778 16668 10784 16720
rect 10836 16708 10842 16720
rect 10836 16680 13584 16708
rect 10836 16668 10842 16680
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 10413 16603 10471 16609
rect 10502 16600 10508 16652
rect 10560 16600 10566 16652
rect 10597 16643 10655 16649
rect 10597 16609 10609 16643
rect 10643 16640 10655 16643
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 10643 16612 10977 16640
rect 10643 16609 10655 16612
rect 10597 16603 10655 16609
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 10965 16603 11023 16609
rect 11236 16612 12909 16640
rect 10520 16572 10548 16600
rect 11236 16572 11264 16612
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 13078 16600 13084 16652
rect 13136 16600 13142 16652
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 10520 16544 11264 16572
rect 12986 16532 12992 16584
rect 13044 16572 13050 16584
rect 13188 16572 13216 16603
rect 13262 16600 13268 16652
rect 13320 16600 13326 16652
rect 13556 16649 13584 16680
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 14016 16708 14044 16736
rect 13688 16680 14044 16708
rect 13688 16668 13694 16680
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 14921 16643 14979 16649
rect 13771 16612 14780 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 13044 16544 13216 16572
rect 13280 16572 13308 16600
rect 13740 16572 13768 16603
rect 14752 16584 14780 16612
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15102 16640 15108 16652
rect 14967 16612 15108 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 15102 16600 15108 16612
rect 15160 16600 15166 16652
rect 13280 16544 13768 16572
rect 13044 16532 13050 16544
rect 10778 16504 10784 16516
rect 9876 16476 10784 16504
rect 10778 16464 10784 16476
rect 10836 16464 10842 16516
rect 13170 16464 13176 16516
rect 13228 16504 13234 16516
rect 13280 16504 13308 16544
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 14274 16572 14280 16584
rect 13872 16544 14280 16572
rect 13872 16532 13878 16544
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 14734 16532 14740 16584
rect 14792 16532 14798 16584
rect 15304 16572 15332 16748
rect 15933 16745 15945 16779
rect 15979 16776 15991 16779
rect 17678 16776 17684 16788
rect 15979 16748 17684 16776
rect 15979 16745 15991 16748
rect 15933 16739 15991 16745
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 17773 16779 17831 16785
rect 17773 16745 17785 16779
rect 17819 16745 17831 16779
rect 18874 16776 18880 16788
rect 17773 16739 17831 16745
rect 18524 16748 18880 16776
rect 16758 16708 16764 16720
rect 15580 16680 16764 16708
rect 15580 16649 15608 16680
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 17788 16708 17816 16739
rect 17788 16680 18460 16708
rect 15565 16643 15623 16649
rect 15565 16609 15577 16643
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15746 16600 15752 16652
rect 15804 16600 15810 16652
rect 16660 16643 16718 16649
rect 16660 16609 16672 16643
rect 16706 16640 16718 16643
rect 17954 16640 17960 16652
rect 16706 16612 17960 16640
rect 16706 16609 16718 16612
rect 16660 16603 16718 16609
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16609 18107 16643
rect 18049 16603 18107 16609
rect 15304 16544 15792 16572
rect 13228 16476 13308 16504
rect 13449 16507 13507 16513
rect 13228 16464 13234 16476
rect 13449 16473 13461 16507
rect 13495 16504 13507 16507
rect 13495 16476 15700 16504
rect 13495 16473 13507 16476
rect 13449 16467 13507 16473
rect 2590 16396 2596 16448
rect 2648 16396 2654 16448
rect 7742 16396 7748 16448
rect 7800 16436 7806 16448
rect 13262 16436 13268 16448
rect 7800 16408 13268 16436
rect 7800 16396 7806 16408
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 15672 16445 15700 16476
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16405 15715 16439
rect 15764 16436 15792 16544
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16390 16572 16396 16584
rect 15896 16544 16396 16572
rect 15896 16532 15902 16544
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 17586 16532 17592 16584
rect 17644 16532 17650 16584
rect 18064 16572 18092 16603
rect 18138 16600 18144 16652
rect 18196 16600 18202 16652
rect 18230 16600 18236 16652
rect 18288 16600 18294 16652
rect 18432 16649 18460 16680
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16609 18475 16643
rect 18417 16603 18475 16609
rect 18524 16572 18552 16748
rect 18874 16736 18880 16748
rect 18932 16776 18938 16788
rect 18932 16748 19472 16776
rect 18932 16736 18938 16748
rect 18782 16668 18788 16720
rect 18840 16668 18846 16720
rect 19052 16711 19110 16717
rect 19052 16677 19064 16711
rect 19098 16708 19110 16711
rect 19334 16708 19340 16720
rect 19098 16680 19340 16708
rect 19098 16677 19110 16680
rect 19052 16671 19110 16677
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 19444 16708 19472 16748
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 22462 16776 22468 16788
rect 19576 16748 22468 16776
rect 19576 16736 19582 16748
rect 20990 16708 20996 16720
rect 19444 16680 20996 16708
rect 20990 16668 20996 16680
rect 21048 16668 21054 16720
rect 21836 16717 21864 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 23106 16776 23112 16788
rect 22940 16748 23112 16776
rect 21821 16711 21879 16717
rect 21821 16677 21833 16711
rect 21867 16677 21879 16711
rect 21821 16671 21879 16677
rect 21913 16711 21971 16717
rect 21913 16677 21925 16711
rect 21959 16708 21971 16711
rect 22554 16708 22560 16720
rect 21959 16680 22560 16708
rect 21959 16677 21971 16680
rect 21913 16671 21971 16677
rect 22554 16668 22560 16680
rect 22612 16668 22618 16720
rect 22830 16708 22836 16720
rect 22664 16680 22836 16708
rect 18800 16640 18828 16668
rect 21542 16640 21548 16652
rect 18800 16612 21548 16640
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 21634 16600 21640 16652
rect 21692 16600 21698 16652
rect 22005 16643 22063 16649
rect 22005 16640 22017 16643
rect 21744 16612 22017 16640
rect 18064 16544 18552 16572
rect 17604 16504 17632 16532
rect 17865 16507 17923 16513
rect 17865 16504 17877 16507
rect 17604 16476 17877 16504
rect 17865 16473 17877 16476
rect 17911 16473 17923 16507
rect 17865 16467 17923 16473
rect 16574 16436 16580 16448
rect 15764 16408 16580 16436
rect 15657 16399 15715 16405
rect 16574 16396 16580 16408
rect 16632 16436 16638 16448
rect 18064 16436 18092 16544
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 18785 16575 18843 16581
rect 18785 16572 18797 16575
rect 18656 16544 18797 16572
rect 18656 16532 18662 16544
rect 18785 16541 18797 16544
rect 18831 16541 18843 16575
rect 18785 16535 18843 16541
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 21744 16572 21772 16612
rect 22005 16609 22017 16612
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 22462 16600 22468 16652
rect 22520 16640 22526 16652
rect 22664 16640 22692 16680
rect 22830 16668 22836 16680
rect 22888 16668 22894 16720
rect 22940 16717 22968 16748
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 23198 16736 23204 16788
rect 23256 16776 23262 16788
rect 23937 16779 23995 16785
rect 23937 16776 23949 16779
rect 23256 16748 23949 16776
rect 23256 16736 23262 16748
rect 23937 16745 23949 16748
rect 23983 16745 23995 16779
rect 24854 16776 24860 16788
rect 23937 16739 23995 16745
rect 24044 16748 24860 16776
rect 22925 16711 22983 16717
rect 22925 16677 22937 16711
rect 22971 16677 22983 16711
rect 24044 16708 24072 16748
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25041 16779 25099 16785
rect 25041 16745 25053 16779
rect 25087 16745 25099 16779
rect 25041 16739 25099 16745
rect 24397 16711 24455 16717
rect 24397 16708 24409 16711
rect 22925 16671 22983 16677
rect 23124 16680 24072 16708
rect 24228 16680 24409 16708
rect 23124 16649 23152 16680
rect 22520 16612 22692 16640
rect 22741 16643 22799 16649
rect 22520 16600 22526 16612
rect 22741 16609 22753 16643
rect 22787 16609 22799 16643
rect 22741 16603 22799 16609
rect 23109 16643 23167 16649
rect 23109 16609 23121 16643
rect 23155 16609 23167 16643
rect 23109 16603 23167 16609
rect 21048 16544 21772 16572
rect 21048 16532 21054 16544
rect 22094 16532 22100 16584
rect 22152 16572 22158 16584
rect 22756 16572 22784 16603
rect 23198 16600 23204 16652
rect 23256 16600 23262 16652
rect 23290 16600 23296 16652
rect 23348 16600 23354 16652
rect 23566 16600 23572 16652
rect 23624 16640 23630 16652
rect 24228 16649 24256 16680
rect 24397 16677 24409 16680
rect 24443 16677 24455 16711
rect 25056 16708 25084 16739
rect 26878 16736 26884 16788
rect 26936 16776 26942 16788
rect 26936 16748 27384 16776
rect 26936 16736 26942 16748
rect 27356 16717 27384 16748
rect 27430 16736 27436 16788
rect 27488 16776 27494 16788
rect 27617 16779 27675 16785
rect 27617 16776 27629 16779
rect 27488 16748 27629 16776
rect 27488 16736 27494 16748
rect 27617 16745 27629 16748
rect 27663 16776 27675 16779
rect 27663 16748 28028 16776
rect 27663 16745 27675 16748
rect 27617 16739 27675 16745
rect 25961 16711 26019 16717
rect 25961 16708 25973 16711
rect 24397 16671 24455 16677
rect 24504 16680 25084 16708
rect 25240 16680 25973 16708
rect 23661 16643 23719 16649
rect 23661 16640 23673 16643
rect 23624 16612 23673 16640
rect 23624 16600 23630 16612
rect 23661 16609 23673 16612
rect 23707 16609 23719 16643
rect 23661 16603 23719 16609
rect 24213 16643 24271 16649
rect 24213 16609 24225 16643
rect 24259 16609 24271 16643
rect 24213 16603 24271 16609
rect 24305 16643 24363 16649
rect 24305 16609 24317 16643
rect 24351 16640 24363 16643
rect 24504 16640 24532 16680
rect 25240 16652 25268 16680
rect 25961 16677 25973 16680
rect 26007 16677 26019 16711
rect 27341 16711 27399 16717
rect 25961 16671 26019 16677
rect 26620 16680 26924 16708
rect 24351 16612 24532 16640
rect 24581 16643 24639 16649
rect 24351 16609 24363 16612
rect 24305 16603 24363 16609
rect 24581 16609 24593 16643
rect 24627 16640 24639 16643
rect 24670 16640 24676 16652
rect 24627 16612 24676 16640
rect 24627 16609 24639 16612
rect 24581 16603 24639 16609
rect 23308 16572 23336 16600
rect 22152 16544 23336 16572
rect 23676 16572 23704 16603
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 24762 16600 24768 16652
rect 24820 16600 24826 16652
rect 25222 16649 25228 16652
rect 25220 16640 25228 16649
rect 25183 16612 25228 16640
rect 25220 16603 25228 16612
rect 25222 16600 25228 16603
rect 25280 16600 25286 16652
rect 25314 16600 25320 16652
rect 25372 16600 25378 16652
rect 25406 16600 25412 16652
rect 25464 16600 25470 16652
rect 25498 16600 25504 16652
rect 25556 16649 25562 16652
rect 25556 16643 25595 16649
rect 25583 16609 25595 16643
rect 25556 16603 25595 16609
rect 25556 16600 25562 16603
rect 25682 16600 25688 16652
rect 25740 16600 25746 16652
rect 26620 16649 26648 16680
rect 26896 16649 26924 16680
rect 27341 16677 27353 16711
rect 27387 16677 27399 16711
rect 28000 16708 28028 16748
rect 28074 16736 28080 16788
rect 28132 16736 28138 16788
rect 28905 16779 28963 16785
rect 28905 16745 28917 16779
rect 28951 16776 28963 16779
rect 29086 16776 29092 16788
rect 28951 16748 29092 16776
rect 28951 16745 28963 16748
rect 28905 16739 28963 16745
rect 29086 16736 29092 16748
rect 29144 16736 29150 16788
rect 29270 16736 29276 16788
rect 29328 16776 29334 16788
rect 29641 16779 29699 16785
rect 29641 16776 29653 16779
rect 29328 16748 29653 16776
rect 29328 16736 29334 16748
rect 29641 16745 29653 16748
rect 29687 16745 29699 16779
rect 29641 16739 29699 16745
rect 29914 16736 29920 16788
rect 29972 16736 29978 16788
rect 31294 16736 31300 16788
rect 31352 16736 31358 16788
rect 29932 16708 29960 16736
rect 30162 16711 30220 16717
rect 30162 16708 30174 16711
rect 28000 16680 29776 16708
rect 29932 16680 30174 16708
rect 27341 16671 27399 16677
rect 27617 16649 27675 16655
rect 26605 16643 26663 16649
rect 26605 16609 26617 16643
rect 26651 16609 26663 16643
rect 26605 16603 26663 16609
rect 26697 16643 26755 16649
rect 26697 16609 26709 16643
rect 26743 16609 26755 16643
rect 26697 16603 26755 16609
rect 26881 16643 26939 16649
rect 26881 16609 26893 16643
rect 26927 16609 26939 16643
rect 26881 16603 26939 16609
rect 27249 16643 27307 16649
rect 27617 16646 27629 16649
rect 27249 16609 27261 16643
rect 27295 16640 27307 16643
rect 27448 16640 27629 16646
rect 27295 16618 27629 16640
rect 27295 16612 27476 16618
rect 27617 16615 27629 16618
rect 27663 16615 27675 16649
rect 27295 16609 27307 16612
rect 27617 16609 27675 16615
rect 27249 16603 27307 16609
rect 26712 16572 26740 16603
rect 23676 16544 26740 16572
rect 26789 16575 26847 16581
rect 22152 16532 22158 16544
rect 26789 16541 26801 16575
rect 26835 16572 26847 16575
rect 26973 16575 27031 16581
rect 26973 16572 26985 16575
rect 26835 16544 26985 16572
rect 26835 16541 26847 16544
rect 26789 16535 26847 16541
rect 26973 16541 26985 16544
rect 27019 16541 27031 16575
rect 26973 16535 27031 16541
rect 27157 16575 27215 16581
rect 27157 16541 27169 16575
rect 27203 16572 27215 16575
rect 27430 16572 27436 16584
rect 27203 16544 27436 16572
rect 27203 16541 27215 16544
rect 27157 16535 27215 16541
rect 27430 16532 27436 16544
rect 27488 16532 27494 16584
rect 27632 16572 27660 16609
rect 27798 16600 27804 16652
rect 27856 16640 27862 16652
rect 28276 16649 28304 16680
rect 27985 16643 28043 16649
rect 27985 16640 27997 16643
rect 27856 16612 27997 16640
rect 27856 16600 27862 16612
rect 27985 16609 27997 16612
rect 28031 16609 28043 16643
rect 27985 16603 28043 16609
rect 28261 16643 28319 16649
rect 28261 16609 28273 16643
rect 28307 16609 28319 16643
rect 28902 16640 28908 16652
rect 28261 16603 28319 16609
rect 28368 16612 28908 16640
rect 27632 16544 27844 16572
rect 25774 16504 25780 16516
rect 19720 16476 25780 16504
rect 16632 16408 18092 16436
rect 16632 16396 16638 16408
rect 18230 16396 18236 16448
rect 18288 16436 18294 16448
rect 19720 16436 19748 16476
rect 25774 16464 25780 16476
rect 25832 16464 25838 16516
rect 27246 16464 27252 16516
rect 27304 16504 27310 16516
rect 27816 16513 27844 16544
rect 27525 16507 27583 16513
rect 27525 16504 27537 16507
rect 27304 16476 27537 16504
rect 27304 16464 27310 16476
rect 27525 16473 27537 16476
rect 27571 16473 27583 16507
rect 27525 16467 27583 16473
rect 27801 16507 27859 16513
rect 27801 16473 27813 16507
rect 27847 16504 27859 16507
rect 28368 16504 28396 16612
rect 28902 16600 28908 16612
rect 28960 16600 28966 16652
rect 29273 16643 29331 16649
rect 29273 16640 29285 16643
rect 29012 16612 29285 16640
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16572 28871 16575
rect 29012 16572 29040 16612
rect 29273 16609 29285 16612
rect 29319 16609 29331 16643
rect 29273 16603 29331 16609
rect 29457 16643 29515 16649
rect 29457 16609 29469 16643
rect 29503 16609 29515 16643
rect 29457 16603 29515 16609
rect 28859 16544 29040 16572
rect 29181 16575 29239 16581
rect 28859 16541 28871 16544
rect 28813 16535 28871 16541
rect 29181 16541 29193 16575
rect 29227 16572 29239 16575
rect 29365 16575 29423 16581
rect 29365 16572 29377 16575
rect 29227 16544 29377 16572
rect 29227 16541 29239 16544
rect 29181 16535 29239 16541
rect 29365 16541 29377 16544
rect 29411 16541 29423 16575
rect 29365 16535 29423 16541
rect 27847 16476 28396 16504
rect 27847 16473 27859 16476
rect 27801 16467 27859 16473
rect 18288 16408 19748 16436
rect 20165 16439 20223 16445
rect 18288 16396 18294 16408
rect 20165 16405 20177 16439
rect 20211 16436 20223 16439
rect 20438 16436 20444 16448
rect 20211 16408 20444 16436
rect 20211 16405 20223 16408
rect 20165 16399 20223 16405
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 22186 16396 22192 16448
rect 22244 16396 22250 16448
rect 22554 16396 22560 16448
rect 22612 16396 22618 16448
rect 23842 16396 23848 16448
rect 23900 16396 23906 16448
rect 24210 16396 24216 16448
rect 24268 16396 24274 16448
rect 27540 16436 27568 16467
rect 28994 16464 29000 16516
rect 29052 16464 29058 16516
rect 29472 16504 29500 16603
rect 29546 16600 29552 16652
rect 29604 16600 29610 16652
rect 29748 16649 29776 16680
rect 30162 16677 30174 16680
rect 30208 16677 30220 16711
rect 30162 16671 30220 16677
rect 29733 16643 29791 16649
rect 29733 16609 29745 16643
rect 29779 16609 29791 16643
rect 29733 16603 29791 16609
rect 29822 16600 29828 16652
rect 29880 16640 29886 16652
rect 29917 16643 29975 16649
rect 29917 16640 29929 16643
rect 29880 16612 29929 16640
rect 29880 16600 29886 16612
rect 29917 16609 29929 16612
rect 29963 16609 29975 16643
rect 29917 16603 29975 16609
rect 29104 16476 29500 16504
rect 29104 16436 29132 16476
rect 27540 16408 29132 16436
rect 552 16346 31648 16368
rect 552 16294 4285 16346
rect 4337 16294 4349 16346
rect 4401 16294 4413 16346
rect 4465 16294 4477 16346
rect 4529 16294 4541 16346
rect 4593 16294 12059 16346
rect 12111 16294 12123 16346
rect 12175 16294 12187 16346
rect 12239 16294 12251 16346
rect 12303 16294 12315 16346
rect 12367 16294 19833 16346
rect 19885 16294 19897 16346
rect 19949 16294 19961 16346
rect 20013 16294 20025 16346
rect 20077 16294 20089 16346
rect 20141 16294 27607 16346
rect 27659 16294 27671 16346
rect 27723 16294 27735 16346
rect 27787 16294 27799 16346
rect 27851 16294 27863 16346
rect 27915 16294 31648 16346
rect 552 16272 31648 16294
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 7742 16232 7748 16244
rect 4755 16204 7748 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 7834 16192 7840 16244
rect 7892 16232 7898 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7892 16204 8033 16232
rect 7892 16192 7898 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 9674 16232 9680 16244
rect 8021 16195 8079 16201
rect 8772 16204 9680 16232
rect 7929 16167 7987 16173
rect 7929 16133 7941 16167
rect 7975 16133 7987 16167
rect 8772 16164 8800 16204
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16232 10195 16235
rect 13357 16235 13415 16241
rect 10183 16204 12848 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 7929 16127 7987 16133
rect 8036 16136 8800 16164
rect 12621 16167 12679 16173
rect 1118 16056 1124 16108
rect 1176 16096 1182 16108
rect 1305 16099 1363 16105
rect 1305 16096 1317 16099
rect 1176 16068 1317 16096
rect 1176 16056 1182 16068
rect 1305 16065 1317 16068
rect 1351 16065 1363 16099
rect 1305 16059 1363 16065
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 1029 16031 1087 16037
rect 1029 15997 1041 16031
rect 1075 15997 1087 16031
rect 1029 15991 1087 15997
rect 1044 15892 1072 15991
rect 1210 15988 1216 16040
rect 1268 15988 1274 16040
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 16028 3387 16031
rect 4982 16028 4988 16040
rect 3375 16000 4988 16028
rect 3375 15997 3387 16000
rect 3329 15991 3387 15997
rect 4982 15988 4988 16000
rect 5040 15988 5046 16040
rect 6816 16031 6874 16037
rect 6816 15997 6828 16031
rect 6862 16028 6874 16031
rect 7098 16028 7104 16040
rect 6862 16000 7104 16028
rect 6862 15997 6874 16000
rect 6816 15991 6874 15997
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 1121 15963 1179 15969
rect 1121 15929 1133 15963
rect 1167 15960 1179 15963
rect 1581 15963 1639 15969
rect 1581 15960 1593 15963
rect 1167 15932 1593 15960
rect 1167 15929 1179 15932
rect 1121 15923 1179 15929
rect 1581 15929 1593 15932
rect 1627 15929 1639 15963
rect 1581 15923 1639 15929
rect 2590 15920 2596 15972
rect 2648 15920 2654 15972
rect 3574 15963 3632 15969
rect 3574 15960 3586 15963
rect 3068 15932 3586 15960
rect 1302 15892 1308 15904
rect 1044 15864 1308 15892
rect 1302 15852 1308 15864
rect 1360 15852 1366 15904
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 3068 15901 3096 15932
rect 3574 15929 3586 15932
rect 3620 15929 3632 15963
rect 3574 15923 3632 15929
rect 5074 15920 5080 15972
rect 5132 15960 5138 15972
rect 5230 15963 5288 15969
rect 5230 15960 5242 15963
rect 5132 15932 5242 15960
rect 5132 15920 5138 15932
rect 5230 15929 5242 15932
rect 5276 15929 5288 15963
rect 7944 15960 7972 16127
rect 8036 16037 8064 16136
rect 12621 16133 12633 16167
rect 12667 16133 12679 16167
rect 12621 16127 12679 16133
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 8680 16068 8769 16096
rect 8680 16040 8708 16068
rect 8757 16065 8769 16068
rect 8803 16065 8815 16099
rect 12526 16096 12532 16108
rect 8757 16059 8815 16065
rect 12452 16068 12532 16096
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8110 15988 8116 16040
rect 8168 16028 8174 16040
rect 8205 16031 8263 16037
rect 8205 16028 8217 16031
rect 8168 16000 8217 16028
rect 8168 15988 8174 16000
rect 8205 15997 8217 16000
rect 8251 15997 8263 16031
rect 8205 15991 8263 15997
rect 8662 15988 8668 16040
rect 8720 15988 8726 16040
rect 9030 16037 9036 16040
rect 9024 16028 9036 16037
rect 8991 16000 9036 16028
rect 9024 15991 9036 16000
rect 9030 15988 9036 15991
rect 9088 15988 9094 16040
rect 10226 15988 10232 16040
rect 10284 15988 10290 16040
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 12452 16037 12480 16068
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 10485 16031 10543 16037
rect 10485 16028 10497 16031
rect 10376 16000 10497 16028
rect 10376 15988 10382 16000
rect 10485 15997 10497 16000
rect 10531 15997 10543 16031
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 10485 15991 10543 15997
rect 10888 16000 12081 16028
rect 10778 15960 10784 15972
rect 7944 15932 10784 15960
rect 5230 15923 5288 15929
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 3053 15895 3111 15901
rect 3053 15892 3065 15895
rect 2464 15864 3065 15892
rect 2464 15852 2470 15864
rect 3053 15861 3065 15864
rect 3099 15861 3111 15895
rect 3053 15855 3111 15861
rect 6365 15895 6423 15901
rect 6365 15861 6377 15895
rect 6411 15892 6423 15895
rect 10888 15892 10916 16000
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12345 16031 12403 16037
rect 12345 16028 12357 16031
rect 12069 15991 12127 15997
rect 12176 16000 12357 16028
rect 10962 15920 10968 15972
rect 11020 15960 11026 15972
rect 12176 15960 12204 16000
rect 12345 15997 12357 16000
rect 12391 15997 12403 16031
rect 12345 15991 12403 15997
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12636 16028 12664 16127
rect 12820 16037 12848 16204
rect 13357 16201 13369 16235
rect 13403 16232 13415 16235
rect 14182 16232 14188 16244
rect 13403 16204 14188 16232
rect 13403 16201 13415 16204
rect 13357 16195 13415 16201
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 15746 16192 15752 16244
rect 15804 16232 15810 16244
rect 16117 16235 16175 16241
rect 16117 16232 16129 16235
rect 15804 16204 16129 16232
rect 15804 16192 15810 16204
rect 16117 16201 16129 16204
rect 16163 16201 16175 16235
rect 16117 16195 16175 16201
rect 16758 16192 16764 16244
rect 16816 16192 16822 16244
rect 17957 16235 18015 16241
rect 17957 16201 17969 16235
rect 18003 16232 18015 16235
rect 18046 16232 18052 16244
rect 18003 16204 18052 16232
rect 18003 16201 18015 16204
rect 17957 16195 18015 16201
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 20530 16232 20536 16244
rect 18380 16204 20536 16232
rect 18380 16192 18386 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 20806 16192 20812 16244
rect 20864 16192 20870 16244
rect 21085 16235 21143 16241
rect 21085 16201 21097 16235
rect 21131 16201 21143 16235
rect 21085 16195 21143 16201
rect 22281 16235 22339 16241
rect 22281 16201 22293 16235
rect 22327 16232 22339 16235
rect 22370 16232 22376 16244
rect 22327 16204 22376 16232
rect 22327 16201 22339 16204
rect 22281 16195 22339 16201
rect 14458 16164 14464 16176
rect 13740 16136 14464 16164
rect 13740 16096 13768 16136
rect 14458 16124 14464 16136
rect 14516 16124 14522 16176
rect 14734 16124 14740 16176
rect 14792 16164 14798 16176
rect 21100 16164 21128 16195
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 22462 16192 22468 16244
rect 22520 16192 22526 16244
rect 22646 16192 22652 16244
rect 22704 16192 22710 16244
rect 24394 16232 24400 16244
rect 22940 16204 24400 16232
rect 21358 16164 21364 16176
rect 14792 16136 19334 16164
rect 14792 16124 14798 16136
rect 14090 16096 14096 16108
rect 13004 16068 13768 16096
rect 13004 16037 13032 16068
rect 13740 16040 13768 16068
rect 13832 16068 14096 16096
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 12636 16000 12725 16028
rect 12437 15991 12495 15997
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 12806 16031 12864 16037
rect 12806 15997 12818 16031
rect 12852 15997 12864 16031
rect 12806 15991 12864 15997
rect 12989 16031 13047 16037
rect 12989 15997 13001 16031
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 13219 16031 13277 16037
rect 13219 15997 13231 16031
rect 13265 16028 13277 16031
rect 13630 16028 13636 16040
rect 13265 16000 13636 16028
rect 13265 15997 13277 16000
rect 13219 15991 13277 15997
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 13722 15988 13728 16040
rect 13780 15988 13786 16040
rect 13832 16037 13860 16068
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 14642 16096 14648 16108
rect 14477 16068 14648 16096
rect 13817 16031 13875 16037
rect 13817 15997 13829 16031
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 13910 16031 13968 16037
rect 13910 15997 13922 16031
rect 13956 15997 13968 16031
rect 14323 16031 14381 16037
rect 14323 16028 14335 16031
rect 13910 15991 13968 15997
rect 14016 16000 14335 16028
rect 11020 15932 12204 15960
rect 12253 15963 12311 15969
rect 11020 15920 11026 15932
rect 12253 15929 12265 15963
rect 12299 15960 12311 15963
rect 12526 15960 12532 15972
rect 12299 15932 12532 15960
rect 12299 15929 12311 15932
rect 12253 15923 12311 15929
rect 12526 15920 12532 15932
rect 12584 15920 12590 15972
rect 13078 15920 13084 15972
rect 13136 15920 13142 15972
rect 13924 15960 13952 15991
rect 13280 15932 13952 15960
rect 6411 15864 10916 15892
rect 11609 15895 11667 15901
rect 6411 15861 6423 15864
rect 6365 15855 6423 15861
rect 11609 15861 11621 15895
rect 11655 15892 11667 15895
rect 13280 15892 13308 15932
rect 11655 15864 13308 15892
rect 11655 15861 11667 15864
rect 11609 15855 11667 15861
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 14016 15892 14044 16000
rect 14323 15997 14335 16000
rect 14369 16028 14381 16031
rect 14477 16028 14505 16068
rect 14642 16056 14648 16068
rect 14700 16096 14706 16108
rect 14700 16068 15148 16096
rect 14700 16056 14706 16068
rect 15120 16040 15148 16068
rect 15562 16056 15568 16108
rect 15620 16096 15626 16108
rect 16025 16099 16083 16105
rect 16025 16096 16037 16099
rect 15620 16068 16037 16096
rect 15620 16056 15626 16068
rect 16025 16065 16037 16068
rect 16071 16065 16083 16099
rect 18230 16096 18236 16108
rect 16025 16059 16083 16065
rect 16316 16068 18236 16096
rect 16316 16040 16344 16068
rect 14369 16000 14505 16028
rect 14369 15997 14381 16000
rect 14323 15991 14381 15997
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 15102 15988 15108 16040
rect 15160 15988 15166 16040
rect 15197 16031 15255 16037
rect 15197 15997 15209 16031
rect 15243 15997 15255 16031
rect 15197 15991 15255 15997
rect 14093 15963 14151 15969
rect 14093 15929 14105 15963
rect 14139 15929 14151 15963
rect 14093 15923 14151 15929
rect 13872 15864 14044 15892
rect 14108 15892 14136 15923
rect 14182 15920 14188 15972
rect 14240 15920 14246 15972
rect 14568 15960 14596 15988
rect 14292 15932 14596 15960
rect 14292 15892 14320 15932
rect 14108 15864 14320 15892
rect 14461 15895 14519 15901
rect 13872 15852 13878 15864
rect 14461 15861 14473 15895
rect 14507 15892 14519 15895
rect 15212 15892 15240 15991
rect 15286 15988 15292 16040
rect 15344 16037 15350 16040
rect 15344 16031 15393 16037
rect 15344 15997 15347 16031
rect 15381 15997 15393 16031
rect 15344 15991 15393 15997
rect 15344 15988 15350 15991
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 16298 15988 16304 16040
rect 16356 15988 16362 16040
rect 16390 15988 16396 16040
rect 16448 15988 16454 16040
rect 16485 16031 16543 16037
rect 16485 15997 16497 16031
rect 16531 16028 16543 16031
rect 16574 16028 16580 16040
rect 16531 16000 16580 16028
rect 16531 15997 16543 16000
rect 16485 15991 16543 15997
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 16669 16031 16727 16037
rect 16669 15997 16681 16031
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17034 16028 17040 16040
rect 16991 16000 17040 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 16684 15960 16712 15991
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 16028 17279 16031
rect 17494 16028 17500 16040
rect 17267 16000 17500 16028
rect 17267 15997 17279 16000
rect 17221 15991 17279 15997
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 17696 16037 17724 16068
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 17681 16031 17739 16037
rect 17681 15997 17693 16031
rect 17727 15997 17739 16031
rect 17681 15991 17739 15997
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 18322 16028 18328 16040
rect 18196 16000 18328 16028
rect 18196 15988 18202 16000
rect 18322 15988 18328 16000
rect 18380 15988 18386 16040
rect 18417 16031 18475 16037
rect 18417 15997 18429 16031
rect 18463 15997 18475 16031
rect 19306 16028 19334 16136
rect 21100 16136 21364 16164
rect 20254 16096 20260 16108
rect 20180 16068 20260 16096
rect 20070 16028 20076 16040
rect 19306 16000 20076 16028
rect 18417 15991 18475 15997
rect 15580 15932 16712 15960
rect 15580 15904 15608 15932
rect 18432 15904 18460 15991
rect 20070 15988 20076 16000
rect 20128 15988 20134 16040
rect 20180 16037 20208 16068
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 21100 16096 21128 16136
rect 21358 16124 21364 16136
rect 21416 16164 21422 16176
rect 22480 16164 22508 16192
rect 21416 16136 22508 16164
rect 21416 16124 21422 16136
rect 20548 16068 21128 16096
rect 21729 16099 21787 16105
rect 20548 16037 20576 16068
rect 21729 16065 21741 16099
rect 21775 16096 21787 16099
rect 21818 16096 21824 16108
rect 21775 16068 21824 16096
rect 21775 16065 21787 16068
rect 21729 16059 21787 16065
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 20165 16031 20223 16037
rect 20165 15997 20177 16031
rect 20211 15997 20223 16031
rect 20165 15991 20223 15997
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 16028 20683 16031
rect 20671 16000 21128 16028
rect 20671 15997 20683 16000
rect 20625 15991 20683 15997
rect 20303 15963 20361 15969
rect 20303 15929 20315 15963
rect 20349 15929 20361 15963
rect 20303 15923 20361 15929
rect 14507 15864 15240 15892
rect 14507 15861 14519 15864
rect 14461 15855 14519 15861
rect 15562 15852 15568 15904
rect 15620 15852 15626 15904
rect 17126 15852 17132 15904
rect 17184 15852 17190 15904
rect 17497 15895 17555 15901
rect 17497 15861 17509 15895
rect 17543 15892 17555 15895
rect 17586 15892 17592 15904
rect 17543 15864 17592 15892
rect 17543 15861 17555 15864
rect 17497 15855 17555 15861
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 18322 15852 18328 15904
rect 18380 15852 18386 15904
rect 18414 15852 18420 15904
rect 18472 15892 18478 15904
rect 19889 15895 19947 15901
rect 19889 15892 19901 15895
rect 18472 15864 19901 15892
rect 18472 15852 18478 15864
rect 19889 15861 19901 15864
rect 19935 15892 19947 15895
rect 20318 15892 20346 15923
rect 20438 15920 20444 15972
rect 20496 15920 20502 15972
rect 20898 15920 20904 15972
rect 20956 15920 20962 15972
rect 21100 15969 21128 16000
rect 21450 15988 21456 16040
rect 21508 15988 21514 16040
rect 22462 16037 22468 16040
rect 22460 16028 22468 16037
rect 21560 16000 22048 16028
rect 22423 16000 22468 16028
rect 21100 15963 21175 15969
rect 21100 15932 21129 15963
rect 21117 15929 21129 15932
rect 21163 15960 21175 15963
rect 21560 15960 21588 16000
rect 22020 15972 22048 16000
rect 22460 15991 22468 16000
rect 22462 15988 22468 15991
rect 22520 15988 22526 16040
rect 22664 16037 22692 16192
rect 22649 16031 22707 16037
rect 22649 15997 22661 16031
rect 22695 15997 22707 16031
rect 22649 15991 22707 15997
rect 22830 15988 22836 16040
rect 22888 15988 22894 16040
rect 22940 16037 22968 16204
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 25498 16192 25504 16244
rect 25556 16192 25562 16244
rect 26326 16192 26332 16244
rect 26384 16232 26390 16244
rect 28997 16235 29055 16241
rect 28997 16232 29009 16235
rect 26384 16204 29009 16232
rect 26384 16192 26390 16204
rect 28997 16201 29009 16204
rect 29043 16201 29055 16235
rect 28997 16195 29055 16201
rect 29472 16204 30420 16232
rect 23842 16124 23848 16176
rect 23900 16124 23906 16176
rect 26694 16124 26700 16176
rect 26752 16124 26758 16176
rect 28537 16167 28595 16173
rect 28537 16164 28549 16167
rect 28092 16136 28549 16164
rect 23860 16096 23888 16124
rect 23860 16068 24256 16096
rect 22925 16031 22983 16037
rect 22925 15997 22937 16031
rect 22971 15997 22983 16031
rect 22925 15991 22983 15997
rect 23014 15988 23020 16040
rect 23072 16028 23078 16040
rect 23201 16031 23259 16037
rect 23201 16028 23213 16031
rect 23072 16000 23213 16028
rect 23072 15988 23078 16000
rect 23201 15997 23213 16000
rect 23247 15997 23259 16031
rect 23201 15991 23259 15997
rect 23569 16031 23627 16037
rect 23569 15997 23581 16031
rect 23615 16028 23627 16031
rect 24026 16028 24032 16040
rect 23615 16000 24032 16028
rect 23615 15997 23627 16000
rect 23569 15991 23627 15997
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24121 16031 24179 16037
rect 24121 15997 24133 16031
rect 24167 15997 24179 16031
rect 24228 16028 24256 16068
rect 28092 16037 28120 16136
rect 28537 16133 28549 16136
rect 28583 16164 28595 16167
rect 28626 16164 28632 16176
rect 28583 16136 28632 16164
rect 28583 16133 28595 16136
rect 28537 16127 28595 16133
rect 28626 16124 28632 16136
rect 28684 16164 28690 16176
rect 29472 16164 29500 16204
rect 28684 16136 29500 16164
rect 28684 16124 28690 16136
rect 28994 16096 29000 16108
rect 28276 16068 29000 16096
rect 28276 16037 28304 16068
rect 28994 16056 29000 16068
rect 29052 16056 29058 16108
rect 30392 16105 30420 16204
rect 30377 16099 30435 16105
rect 30377 16065 30389 16099
rect 30423 16065 30435 16099
rect 30377 16059 30435 16065
rect 28077 16031 28135 16037
rect 28077 16028 28089 16031
rect 24228 16000 24348 16028
rect 24121 15991 24179 15997
rect 21163 15932 21588 15960
rect 21163 15929 21175 15932
rect 21117 15923 21175 15929
rect 22002 15920 22008 15972
rect 22060 15920 22066 15972
rect 22278 15920 22284 15972
rect 22336 15960 22342 15972
rect 22557 15963 22615 15969
rect 22557 15960 22569 15963
rect 22336 15932 22569 15960
rect 22336 15920 22342 15932
rect 22557 15929 22569 15932
rect 22603 15929 22615 15963
rect 22557 15923 22615 15929
rect 23293 15963 23351 15969
rect 23293 15929 23305 15963
rect 23339 15929 23351 15963
rect 23293 15923 23351 15929
rect 19935 15864 20346 15892
rect 19935 15861 19947 15864
rect 19889 15855 19947 15861
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 21542 15852 21548 15904
rect 21600 15892 21606 15904
rect 23017 15895 23075 15901
rect 23017 15892 23029 15895
rect 21600 15864 23029 15892
rect 21600 15852 21606 15864
rect 23017 15861 23029 15864
rect 23063 15861 23075 15895
rect 23308 15892 23336 15923
rect 23382 15920 23388 15972
rect 23440 15920 23446 15972
rect 24136 15960 24164 15991
rect 24320 15960 24348 16000
rect 27908 16000 28089 16028
rect 24377 15963 24435 15969
rect 24377 15960 24389 15963
rect 24136 15932 24256 15960
rect 24320 15932 24389 15960
rect 24118 15892 24124 15904
rect 23308 15864 24124 15892
rect 23017 15855 23075 15861
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 24228 15892 24256 15932
rect 24377 15929 24389 15932
rect 24423 15929 24435 15963
rect 24377 15923 24435 15929
rect 27154 15920 27160 15972
rect 27212 15960 27218 15972
rect 27810 15963 27868 15969
rect 27810 15960 27822 15963
rect 27212 15932 27822 15960
rect 27212 15920 27218 15932
rect 27810 15929 27822 15932
rect 27856 15929 27868 15963
rect 27810 15923 27868 15929
rect 25866 15892 25872 15904
rect 24228 15864 25872 15892
rect 25866 15852 25872 15864
rect 25924 15892 25930 15904
rect 27908 15892 27936 16000
rect 28077 15997 28089 16000
rect 28123 15997 28135 16031
rect 28077 15991 28135 15997
rect 28261 16031 28319 16037
rect 28261 15997 28273 16031
rect 28307 15997 28319 16031
rect 30110 16031 30168 16037
rect 30110 16028 30122 16031
rect 28261 15991 28319 15997
rect 28460 16000 30122 16028
rect 28460 15901 28488 16000
rect 30110 15997 30122 16000
rect 30156 15997 30168 16031
rect 30110 15991 30168 15997
rect 28721 15963 28779 15969
rect 28721 15929 28733 15963
rect 28767 15960 28779 15963
rect 29638 15960 29644 15972
rect 28767 15932 29644 15960
rect 28767 15929 28779 15932
rect 28721 15923 28779 15929
rect 29638 15920 29644 15932
rect 29696 15920 29702 15972
rect 25924 15864 27936 15892
rect 28445 15895 28503 15901
rect 25924 15852 25930 15864
rect 28445 15861 28457 15895
rect 28491 15861 28503 15895
rect 28445 15855 28503 15861
rect 552 15802 31808 15824
rect 552 15750 8172 15802
rect 8224 15750 8236 15802
rect 8288 15750 8300 15802
rect 8352 15750 8364 15802
rect 8416 15750 8428 15802
rect 8480 15750 15946 15802
rect 15998 15750 16010 15802
rect 16062 15750 16074 15802
rect 16126 15750 16138 15802
rect 16190 15750 16202 15802
rect 16254 15750 23720 15802
rect 23772 15750 23784 15802
rect 23836 15750 23848 15802
rect 23900 15750 23912 15802
rect 23964 15750 23976 15802
rect 24028 15750 31494 15802
rect 31546 15750 31558 15802
rect 31610 15750 31622 15802
rect 31674 15750 31686 15802
rect 31738 15750 31750 15802
rect 31802 15750 31808 15802
rect 552 15728 31808 15750
rect 1210 15648 1216 15700
rect 1268 15648 1274 15700
rect 1302 15648 1308 15700
rect 1360 15688 1366 15700
rect 1489 15691 1547 15697
rect 1489 15688 1501 15691
rect 1360 15660 1501 15688
rect 1360 15648 1366 15660
rect 1489 15657 1501 15660
rect 1535 15657 1547 15691
rect 2225 15691 2283 15697
rect 2225 15688 2237 15691
rect 1489 15651 1547 15657
rect 1688 15660 2237 15688
rect 1228 15620 1256 15648
rect 1688 15620 1716 15660
rect 2225 15657 2237 15660
rect 2271 15657 2283 15691
rect 2406 15688 2412 15700
rect 2225 15651 2283 15657
rect 2332 15660 2412 15688
rect 1228 15592 1716 15620
rect 1765 15623 1823 15629
rect 1765 15589 1777 15623
rect 1811 15620 1823 15623
rect 2332 15620 2360 15660
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3694 15688 3700 15700
rect 3108 15660 3700 15688
rect 3108 15648 3114 15660
rect 3694 15648 3700 15660
rect 3752 15688 3758 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 3752 15660 3801 15688
rect 3752 15648 3758 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 7466 15688 7472 15700
rect 7423 15660 7472 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 10689 15691 10747 15697
rect 9539 15660 10640 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 8036 15620 8064 15651
rect 8358 15623 8416 15629
rect 8358 15620 8370 15623
rect 1811 15592 2360 15620
rect 2424 15592 3004 15620
rect 1811 15589 1823 15592
rect 1765 15583 1823 15589
rect 2148 15561 2176 15592
rect 2424 15561 2452 15592
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15521 1731 15555
rect 1673 15515 1731 15521
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15521 2191 15555
rect 2409 15555 2467 15561
rect 2409 15552 2421 15555
rect 2133 15515 2191 15521
rect 2240 15524 2421 15552
rect 1688 15360 1716 15515
rect 1872 15484 1900 15515
rect 2240 15484 2268 15524
rect 2409 15521 2421 15524
rect 2455 15521 2467 15555
rect 2409 15515 2467 15521
rect 2501 15555 2559 15561
rect 2501 15521 2513 15555
rect 2547 15521 2559 15555
rect 2501 15515 2559 15521
rect 1872 15456 2268 15484
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15453 2375 15487
rect 2317 15447 2375 15453
rect 2038 15376 2044 15428
rect 2096 15416 2102 15428
rect 2332 15416 2360 15447
rect 2096 15388 2360 15416
rect 2516 15416 2544 15515
rect 2976 15496 3004 15592
rect 3896 15592 5764 15620
rect 8036 15592 8370 15620
rect 3896 15564 3924 15592
rect 5736 15564 5764 15592
rect 8358 15589 8370 15592
rect 8404 15589 8416 15623
rect 9769 15623 9827 15629
rect 9769 15620 9781 15623
rect 8358 15583 8416 15589
rect 8680 15592 9781 15620
rect 8680 15564 8708 15592
rect 9769 15589 9781 15592
rect 9815 15589 9827 15623
rect 9769 15583 9827 15589
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15521 3663 15555
rect 3605 15515 3663 15521
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3620 15484 3648 15515
rect 3878 15512 3884 15564
rect 3936 15512 3942 15564
rect 4706 15512 4712 15564
rect 4764 15552 4770 15564
rect 5077 15555 5135 15561
rect 5077 15552 5089 15555
rect 4764 15524 5089 15552
rect 4764 15512 4770 15524
rect 5077 15521 5089 15524
rect 5123 15552 5135 15555
rect 5353 15555 5411 15561
rect 5353 15552 5365 15555
rect 5123 15524 5365 15552
rect 5123 15521 5135 15524
rect 5077 15515 5135 15521
rect 5353 15521 5365 15524
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 5718 15512 5724 15564
rect 5776 15512 5782 15564
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 7374 15552 7380 15564
rect 7331 15524 7380 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 7374 15512 7380 15524
rect 7432 15512 7438 15564
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15552 7527 15555
rect 7561 15555 7619 15561
rect 7561 15552 7573 15555
rect 7515 15524 7573 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 7561 15521 7573 15524
rect 7607 15521 7619 15555
rect 7561 15515 7619 15521
rect 7834 15512 7840 15564
rect 7892 15552 7898 15564
rect 8018 15552 8024 15564
rect 7892 15524 8024 15552
rect 7892 15512 7898 15524
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8662 15552 8668 15564
rect 8128 15524 8668 15552
rect 3016 15456 5120 15484
rect 3016 15444 3022 15456
rect 5092 15428 5120 15456
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 7650 15484 7656 15496
rect 6604 15456 7656 15484
rect 6604 15444 6610 15456
rect 7650 15444 7656 15456
rect 7708 15484 7714 15496
rect 8128 15493 8156 15524
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 9364 15524 9597 15552
rect 9364 15512 9370 15524
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 10410 15512 10416 15564
rect 10468 15552 10474 15564
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 10468 15524 10517 15552
rect 10468 15512 10474 15524
rect 10505 15521 10517 15524
rect 10551 15521 10563 15555
rect 10612 15552 10640 15660
rect 10689 15657 10701 15691
rect 10735 15657 10747 15691
rect 14182 15688 14188 15700
rect 10689 15651 10747 15657
rect 12406 15660 14188 15688
rect 10704 15620 10732 15651
rect 11210 15623 11268 15629
rect 11210 15620 11222 15623
rect 10704 15592 11222 15620
rect 11210 15589 11222 15592
rect 11256 15589 11268 15623
rect 11210 15583 11268 15589
rect 12406 15552 12434 15660
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 14274 15648 14280 15700
rect 14332 15648 14338 15700
rect 14458 15648 14464 15700
rect 14516 15648 14522 15700
rect 15470 15648 15476 15700
rect 15528 15648 15534 15700
rect 18506 15648 18512 15700
rect 18564 15648 18570 15700
rect 20257 15691 20315 15697
rect 20257 15657 20269 15691
rect 20303 15688 20315 15691
rect 20898 15688 20904 15700
rect 20303 15660 20904 15688
rect 20303 15657 20315 15660
rect 20257 15651 20315 15657
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 21450 15648 21456 15700
rect 21508 15688 21514 15700
rect 21637 15691 21695 15697
rect 21637 15688 21649 15691
rect 21508 15660 21649 15688
rect 21508 15648 21514 15660
rect 21637 15657 21649 15660
rect 21683 15657 21695 15691
rect 21637 15651 21695 15657
rect 22278 15648 22284 15700
rect 22336 15688 22342 15700
rect 22336 15660 26087 15688
rect 22336 15648 22342 15660
rect 13630 15620 13636 15632
rect 12999 15592 13636 15620
rect 10612 15524 12434 15552
rect 10505 15515 10563 15521
rect 12618 15512 12624 15564
rect 12676 15552 12682 15564
rect 12999 15561 13027 15592
rect 13630 15580 13636 15592
rect 13688 15620 13694 15632
rect 14476 15620 14504 15648
rect 13688 15592 14136 15620
rect 13688 15580 13694 15592
rect 14108 15564 14136 15592
rect 14200 15592 14504 15620
rect 15488 15620 15516 15648
rect 22094 15620 22100 15632
rect 15488 15592 21036 15620
rect 14200 15564 14228 15592
rect 12984 15555 13042 15561
rect 12676 15524 12940 15552
rect 12676 15512 12682 15524
rect 8113 15487 8171 15493
rect 8113 15484 8125 15487
rect 7708 15456 8125 15484
rect 7708 15444 7714 15456
rect 8113 15453 8125 15456
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10962 15484 10968 15496
rect 10284 15456 10968 15484
rect 10284 15444 10290 15456
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 12912 15484 12940 15524
rect 12984 15521 12996 15555
rect 13030 15521 13042 15555
rect 12984 15515 13042 15521
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15521 13139 15555
rect 13081 15515 13139 15521
rect 13096 15484 13124 15515
rect 13170 15512 13176 15564
rect 13228 15512 13234 15564
rect 13262 15512 13268 15564
rect 13320 15561 13326 15564
rect 13320 15555 13359 15561
rect 13347 15521 13359 15555
rect 13320 15515 13359 15521
rect 13320 15512 13326 15515
rect 13446 15512 13452 15564
rect 13504 15512 13510 15564
rect 13541 15555 13599 15561
rect 13541 15521 13553 15555
rect 13587 15521 13599 15555
rect 13541 15515 13599 15521
rect 12912 15456 13124 15484
rect 3878 15416 3884 15428
rect 2516 15388 3884 15416
rect 2096 15376 2102 15388
rect 1670 15308 1676 15360
rect 1728 15348 1734 15360
rect 2516 15348 2544 15388
rect 3878 15376 3884 15388
rect 3936 15376 3942 15428
rect 5074 15376 5080 15428
rect 5132 15376 5138 15428
rect 1728 15320 2544 15348
rect 1728 15308 1734 15320
rect 3418 15308 3424 15360
rect 3476 15308 3482 15360
rect 5261 15351 5319 15357
rect 5261 15317 5273 15351
rect 5307 15348 5319 15351
rect 5534 15348 5540 15360
rect 5307 15320 5540 15348
rect 5307 15317 5319 15320
rect 5261 15311 5319 15317
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15348 12403 15351
rect 12434 15348 12440 15360
rect 12391 15320 12440 15348
rect 12391 15317 12403 15320
rect 12345 15311 12403 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 12820 15357 12848 15444
rect 13170 15376 13176 15428
rect 13228 15416 13234 15428
rect 13556 15416 13584 15515
rect 13722 15512 13728 15564
rect 13780 15512 13786 15564
rect 13814 15512 13820 15564
rect 13872 15512 13878 15564
rect 13906 15512 13912 15564
rect 13964 15512 13970 15564
rect 14090 15512 14096 15564
rect 14148 15512 14154 15564
rect 14182 15512 14188 15564
rect 14240 15512 14246 15564
rect 14461 15555 14519 15561
rect 14461 15521 14473 15555
rect 14507 15552 14519 15555
rect 15010 15552 15016 15564
rect 14507 15524 15016 15552
rect 14507 15521 14519 15524
rect 14461 15515 14519 15521
rect 13998 15444 14004 15496
rect 14056 15484 14062 15496
rect 14476 15484 14504 15515
rect 15010 15512 15016 15524
rect 15068 15552 15074 15564
rect 15068 15524 15332 15552
rect 15068 15512 15074 15524
rect 14056 15456 14504 15484
rect 14056 15444 14062 15456
rect 13228 15388 13584 15416
rect 14093 15419 14151 15425
rect 13228 15376 13234 15388
rect 14093 15385 14105 15419
rect 14139 15416 14151 15419
rect 15194 15416 15200 15428
rect 14139 15388 15200 15416
rect 14139 15385 14151 15388
rect 14093 15379 14151 15385
rect 15194 15376 15200 15388
rect 15252 15376 15258 15428
rect 15304 15416 15332 15524
rect 15470 15512 15476 15564
rect 15528 15552 15534 15564
rect 17589 15555 17647 15561
rect 17589 15552 17601 15555
rect 15528 15524 17601 15552
rect 15528 15512 15534 15524
rect 17589 15521 17601 15524
rect 17635 15521 17647 15555
rect 17589 15515 17647 15521
rect 17770 15512 17776 15564
rect 17828 15512 17834 15564
rect 18138 15512 18144 15564
rect 18196 15512 18202 15564
rect 18966 15512 18972 15564
rect 19024 15552 19030 15564
rect 19133 15555 19191 15561
rect 19133 15552 19145 15555
rect 19024 15524 19145 15552
rect 19024 15512 19030 15524
rect 19133 15521 19145 15524
rect 19179 15521 19191 15555
rect 19133 15515 19191 15521
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15804 15456 16129 15484
rect 15804 15444 15810 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 16298 15444 16304 15496
rect 16356 15484 16362 15496
rect 16393 15487 16451 15493
rect 16393 15484 16405 15487
rect 16356 15456 16405 15484
rect 16356 15444 16362 15456
rect 16393 15453 16405 15456
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 17052 15416 17080 15444
rect 15304 15388 17080 15416
rect 18340 15416 18368 15447
rect 18782 15444 18788 15496
rect 18840 15484 18846 15496
rect 18877 15487 18935 15493
rect 18877 15484 18889 15487
rect 18840 15456 18889 15484
rect 18840 15444 18846 15456
rect 18877 15453 18889 15456
rect 18923 15453 18935 15487
rect 21008 15484 21036 15592
rect 21468 15592 22100 15620
rect 21358 15512 21364 15564
rect 21416 15512 21422 15564
rect 21468 15561 21496 15592
rect 22094 15580 22100 15592
rect 22152 15580 22158 15632
rect 22370 15580 22376 15632
rect 22428 15620 22434 15632
rect 24029 15623 24087 15629
rect 24029 15620 24041 15623
rect 22428 15592 24041 15620
rect 22428 15580 22434 15592
rect 24029 15589 24041 15592
rect 24075 15589 24087 15623
rect 24029 15583 24087 15589
rect 24121 15623 24179 15629
rect 24121 15589 24133 15623
rect 24167 15620 24179 15623
rect 25222 15620 25228 15632
rect 24167 15592 25228 15620
rect 24167 15589 24179 15592
rect 24121 15583 24179 15589
rect 21453 15555 21511 15561
rect 21453 15521 21465 15555
rect 21499 15521 21511 15555
rect 21453 15515 21511 15521
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 22465 15555 22523 15561
rect 22465 15521 22477 15555
rect 22511 15552 22523 15555
rect 22554 15552 22560 15564
rect 22511 15524 22560 15552
rect 22511 15521 22523 15524
rect 22465 15515 22523 15521
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 23566 15512 23572 15564
rect 23624 15552 23630 15564
rect 23845 15555 23903 15561
rect 23845 15552 23857 15555
rect 23624 15524 23857 15552
rect 23624 15512 23630 15524
rect 23845 15521 23857 15524
rect 23891 15521 23903 15555
rect 23845 15515 23903 15521
rect 24044 15484 24072 15583
rect 25222 15580 25228 15592
rect 25280 15580 25286 15632
rect 25774 15580 25780 15632
rect 25832 15580 25838 15632
rect 25866 15580 25872 15632
rect 25924 15580 25930 15632
rect 25958 15580 25964 15632
rect 26016 15629 26022 15632
rect 26016 15583 26028 15629
rect 26059 15620 26087 15660
rect 27154 15648 27160 15700
rect 27212 15648 27218 15700
rect 27985 15691 28043 15697
rect 27985 15657 27997 15691
rect 28031 15657 28043 15691
rect 27985 15651 28043 15657
rect 28000 15620 28028 15651
rect 29086 15648 29092 15700
rect 29144 15688 29150 15700
rect 29144 15660 30205 15688
rect 29144 15648 29150 15660
rect 30177 15629 30205 15660
rect 30374 15648 30380 15700
rect 30432 15688 30438 15700
rect 31297 15691 31355 15697
rect 31297 15688 31309 15691
rect 30432 15660 31309 15688
rect 30432 15648 30438 15660
rect 31297 15657 31309 15660
rect 31343 15657 31355 15691
rect 31297 15651 31355 15657
rect 30162 15623 30220 15629
rect 26059 15592 28028 15620
rect 28736 15592 29500 15620
rect 26016 15580 26022 15583
rect 24213 15555 24271 15561
rect 24213 15521 24225 15555
rect 24259 15552 24271 15555
rect 25792 15552 25820 15580
rect 24259 15524 25820 15552
rect 25884 15552 25912 15580
rect 26237 15555 26295 15561
rect 26237 15552 26249 15555
rect 25884 15524 26249 15552
rect 24259 15521 24271 15524
rect 24213 15515 24271 15521
rect 26237 15521 26249 15524
rect 26283 15521 26295 15555
rect 26237 15515 26295 15521
rect 26973 15555 27031 15561
rect 26973 15521 26985 15555
rect 27019 15552 27031 15555
rect 27246 15552 27252 15564
rect 27019 15524 27252 15552
rect 27019 15521 27031 15524
rect 26973 15515 27031 15521
rect 27246 15512 27252 15524
rect 27304 15512 27310 15564
rect 27982 15512 27988 15564
rect 28040 15552 28046 15564
rect 28350 15552 28356 15564
rect 28040 15524 28356 15552
rect 28040 15512 28046 15524
rect 28350 15512 28356 15524
rect 28408 15552 28414 15564
rect 28736 15552 28764 15592
rect 28408 15524 28764 15552
rect 28408 15512 28414 15524
rect 28810 15512 28816 15564
rect 28868 15552 28874 15564
rect 29472 15561 29500 15592
rect 30162 15589 30174 15623
rect 30208 15589 30220 15623
rect 30162 15583 30220 15589
rect 29098 15555 29156 15561
rect 29098 15552 29110 15555
rect 28868 15524 29110 15552
rect 28868 15512 28874 15524
rect 29098 15521 29110 15524
rect 29144 15521 29156 15555
rect 29098 15515 29156 15521
rect 29457 15555 29515 15561
rect 29457 15521 29469 15555
rect 29503 15521 29515 15555
rect 29457 15515 29515 15521
rect 24670 15484 24676 15496
rect 21008 15456 22692 15484
rect 24044 15456 24676 15484
rect 18877 15447 18935 15453
rect 22664 15425 22692 15456
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 29365 15487 29423 15493
rect 29365 15453 29377 15487
rect 29411 15484 29423 15487
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29411 15456 29929 15484
rect 29411 15453 29423 15456
rect 29365 15447 29423 15453
rect 29917 15453 29929 15456
rect 29963 15453 29975 15487
rect 29917 15447 29975 15453
rect 22649 15419 22707 15425
rect 18340 15388 18920 15416
rect 12805 15351 12863 15357
rect 12805 15317 12817 15351
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 14645 15351 14703 15357
rect 14645 15317 14657 15351
rect 14691 15348 14703 15351
rect 15378 15348 15384 15360
rect 14691 15320 15384 15348
rect 14691 15317 14703 15320
rect 14645 15311 14703 15317
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 18892 15348 18920 15388
rect 22649 15385 22661 15419
rect 22695 15385 22707 15419
rect 22649 15379 22707 15385
rect 24394 15376 24400 15428
rect 24452 15376 24458 15428
rect 20714 15348 20720 15360
rect 18892 15320 20720 15348
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 22186 15308 22192 15360
rect 22244 15348 22250 15360
rect 22281 15351 22339 15357
rect 22281 15348 22293 15351
rect 22244 15320 22293 15348
rect 22244 15308 22250 15320
rect 22281 15317 22293 15320
rect 22327 15317 22339 15351
rect 22281 15311 22339 15317
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 23014 15348 23020 15360
rect 22520 15320 23020 15348
rect 22520 15308 22526 15320
rect 23014 15308 23020 15320
rect 23072 15308 23078 15360
rect 24486 15308 24492 15360
rect 24544 15348 24550 15360
rect 24857 15351 24915 15357
rect 24857 15348 24869 15351
rect 24544 15320 24869 15348
rect 24544 15308 24550 15320
rect 24857 15317 24869 15320
rect 24903 15317 24915 15351
rect 24857 15311 24915 15317
rect 28626 15308 28632 15360
rect 28684 15348 28690 15360
rect 29380 15348 29408 15447
rect 28684 15320 29408 15348
rect 28684 15308 28690 15320
rect 552 15258 31648 15280
rect 552 15206 4285 15258
rect 4337 15206 4349 15258
rect 4401 15206 4413 15258
rect 4465 15206 4477 15258
rect 4529 15206 4541 15258
rect 4593 15206 12059 15258
rect 12111 15206 12123 15258
rect 12175 15206 12187 15258
rect 12239 15206 12251 15258
rect 12303 15206 12315 15258
rect 12367 15206 19833 15258
rect 19885 15206 19897 15258
rect 19949 15206 19961 15258
rect 20013 15206 20025 15258
rect 20077 15206 20089 15258
rect 20141 15206 27607 15258
rect 27659 15206 27671 15258
rect 27723 15206 27735 15258
rect 27787 15206 27799 15258
rect 27851 15206 27863 15258
rect 27915 15206 31648 15258
rect 552 15184 31648 15206
rect 5074 15104 5080 15156
rect 5132 15104 5138 15156
rect 7926 15104 7932 15156
rect 7984 15144 7990 15156
rect 9674 15144 9680 15156
rect 7984 15116 8708 15144
rect 7984 15104 7990 15116
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 8573 15079 8631 15085
rect 8573 15076 8585 15079
rect 7892 15048 8585 15076
rect 7892 15036 7898 15048
rect 8573 15045 8585 15048
rect 8619 15045 8631 15079
rect 8573 15039 8631 15045
rect 4982 14968 4988 15020
rect 5040 15008 5046 15020
rect 5442 15008 5448 15020
rect 5040 14980 5448 15008
rect 5040 14968 5046 14980
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 8113 15011 8171 15017
rect 7432 14980 7972 15008
rect 7432 14968 7438 14980
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 2958 14940 2964 14952
rect 2915 14912 2964 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3050 14900 3056 14952
rect 3108 14900 3114 14952
rect 3326 14900 3332 14952
rect 3384 14900 3390 14952
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 5701 14943 5759 14949
rect 5701 14940 5713 14943
rect 5592 14912 5713 14940
rect 5592 14900 5598 14912
rect 5701 14909 5713 14912
rect 5747 14909 5759 14943
rect 5701 14903 5759 14909
rect 7293 14943 7351 14949
rect 7293 14909 7305 14943
rect 7339 14940 7351 14943
rect 7392 14940 7420 14968
rect 7339 14912 7420 14940
rect 7339 14909 7351 14912
rect 7293 14903 7351 14909
rect 7558 14900 7564 14952
rect 7616 14900 7622 14952
rect 7742 14900 7748 14952
rect 7800 14900 7806 14952
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 7944 14949 7972 14980
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8159 14980 8616 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 7975 14912 8524 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 3068 14872 3096 14900
rect 2884 14844 3096 14872
rect 2884 14816 2912 14844
rect 3602 14832 3608 14884
rect 3660 14832 3666 14884
rect 4338 14832 4344 14884
rect 4396 14832 4402 14884
rect 7653 14875 7711 14881
rect 7653 14841 7665 14875
rect 7699 14872 7711 14875
rect 8389 14875 8447 14881
rect 8389 14872 8401 14875
rect 7699 14844 8401 14872
rect 7699 14841 7711 14844
rect 7653 14835 7711 14841
rect 8389 14841 8401 14844
rect 8435 14841 8447 14875
rect 8389 14835 8447 14841
rect 2866 14764 2872 14816
rect 2924 14764 2930 14816
rect 3050 14764 3056 14816
rect 3108 14764 3114 14816
rect 6822 14764 6828 14816
rect 6880 14764 6886 14816
rect 7466 14764 7472 14816
rect 7524 14764 7530 14816
rect 8496 14804 8524 14912
rect 8588 14872 8616 14980
rect 8680 14952 8708 15116
rect 8772 15116 9680 15144
rect 8662 14900 8668 14952
rect 8720 14900 8726 14952
rect 8772 14949 8800 15116
rect 9674 15104 9680 15116
rect 9732 15144 9738 15156
rect 10502 15144 10508 15156
rect 9732 15116 10508 15144
rect 9732 15104 9738 15116
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 12253 15147 12311 15153
rect 10827 15116 12204 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 12176 15076 12204 15116
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 13814 15144 13820 15156
rect 12299 15116 13820 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 14182 15104 14188 15156
rect 14240 15104 14246 15156
rect 15194 15104 15200 15156
rect 15252 15104 15258 15156
rect 15286 15104 15292 15156
rect 15344 15104 15350 15156
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 16482 15144 16488 15156
rect 15519 15116 16488 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 17681 15147 17739 15153
rect 16684 15116 17080 15144
rect 13170 15076 13176 15088
rect 12176 15048 13176 15076
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 14200 15008 14228 15104
rect 15013 15079 15071 15085
rect 15013 15045 15025 15079
rect 15059 15076 15071 15079
rect 15304 15076 15332 15104
rect 15059 15048 15332 15076
rect 15059 15045 15071 15048
rect 15013 15039 15071 15045
rect 15197 15011 15255 15017
rect 13832 14980 14688 15008
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14909 8815 14943
rect 8757 14903 8815 14909
rect 8953 14943 9011 14949
rect 8953 14909 8965 14943
rect 8999 14940 9011 14943
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8999 14912 9137 14940
rect 8999 14909 9011 14912
rect 8953 14903 9011 14909
rect 9125 14909 9137 14912
rect 9171 14940 9183 14943
rect 9171 14912 9260 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 8849 14875 8907 14881
rect 8849 14872 8861 14875
rect 8588 14844 8861 14872
rect 8849 14841 8861 14844
rect 8895 14841 8907 14875
rect 8849 14835 8907 14841
rect 9232 14816 9260 14912
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 9364 14912 9413 14940
rect 9364 14900 9370 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 10873 14943 10931 14949
rect 10873 14909 10885 14943
rect 10919 14940 10931 14943
rect 10962 14940 10968 14952
rect 10919 14912 10968 14940
rect 10919 14909 10931 14912
rect 10873 14903 10931 14909
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 12434 14900 12440 14952
rect 12492 14900 12498 14952
rect 13538 14900 13544 14952
rect 13596 14900 13602 14952
rect 13630 14900 13636 14952
rect 13688 14900 13694 14952
rect 13832 14949 13860 14980
rect 14090 14949 14096 14952
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 14047 14943 14096 14949
rect 14047 14909 14059 14943
rect 14093 14909 14096 14943
rect 14047 14903 14096 14909
rect 14090 14900 14096 14903
rect 14148 14900 14154 14952
rect 14182 14900 14188 14952
rect 14240 14940 14246 14952
rect 14660 14949 14688 14980
rect 14844 14980 15056 15008
rect 14844 14952 14872 14980
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 14240 14912 14381 14940
rect 14240 14900 14246 14912
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 14462 14943 14520 14949
rect 14462 14909 14474 14943
rect 14508 14909 14520 14943
rect 14462 14903 14520 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 9646 14875 9704 14881
rect 9646 14872 9658 14875
rect 9324 14844 9658 14872
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8496 14776 8677 14804
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 9214 14764 9220 14816
rect 9272 14764 9278 14816
rect 9324 14813 9352 14844
rect 9646 14841 9658 14844
rect 9692 14841 9704 14875
rect 9646 14835 9704 14841
rect 10226 14832 10232 14884
rect 10284 14872 10290 14884
rect 11118 14875 11176 14881
rect 11118 14872 11130 14875
rect 10284 14844 11130 14872
rect 10284 14832 10290 14844
rect 11118 14841 11130 14844
rect 11164 14841 11176 14875
rect 12452 14872 12480 14900
rect 12452 14844 13860 14872
rect 11118 14835 11176 14841
rect 9309 14807 9367 14813
rect 9309 14773 9321 14807
rect 9355 14773 9367 14807
rect 9309 14767 9367 14773
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 13722 14804 13728 14816
rect 9548 14776 13728 14804
rect 9548 14764 9554 14776
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 13832 14804 13860 14844
rect 13906 14832 13912 14884
rect 13964 14832 13970 14884
rect 14477 14872 14505 14903
rect 14826 14900 14832 14952
rect 14884 14949 14890 14952
rect 14884 14903 14892 14949
rect 14884 14900 14890 14903
rect 14108 14844 14505 14872
rect 14108 14804 14136 14844
rect 14734 14832 14740 14884
rect 14792 14832 14798 14884
rect 15028 14872 15056 14980
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15378 15008 15384 15020
rect 15243 14980 15384 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15102 14900 15108 14952
rect 15160 14900 15166 14952
rect 15565 14943 15623 14949
rect 15565 14909 15577 14943
rect 15611 14940 15623 14943
rect 16298 14940 16304 14952
rect 15611 14912 16304 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 16298 14900 16304 14912
rect 16356 14900 16362 14952
rect 15028 14844 15332 14872
rect 13832 14776 14136 14804
rect 14185 14807 14243 14813
rect 14185 14773 14197 14807
rect 14231 14804 14243 14807
rect 15194 14804 15200 14816
rect 14231 14776 15200 14804
rect 14231 14773 14243 14776
rect 14185 14767 14243 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 15304 14804 15332 14844
rect 15654 14832 15660 14884
rect 15712 14872 15718 14884
rect 15810 14875 15868 14881
rect 15810 14872 15822 14875
rect 15712 14844 15822 14872
rect 15712 14832 15718 14844
rect 15810 14841 15822 14844
rect 15856 14841 15868 14875
rect 15810 14835 15868 14841
rect 15930 14832 15936 14884
rect 15988 14872 15994 14884
rect 16684 14872 16712 15116
rect 16945 15079 17003 15085
rect 16945 15045 16957 15079
rect 16991 15045 17003 15079
rect 17052 15076 17080 15116
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 17770 15144 17776 15156
rect 17727 15116 17776 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 22848 15116 24808 15144
rect 19337 15079 19395 15085
rect 19337 15076 19349 15079
rect 17052 15048 19349 15076
rect 16945 15039 17003 15045
rect 19337 15045 19349 15048
rect 19383 15045 19395 15079
rect 19337 15039 19395 15045
rect 16960 15008 16988 15039
rect 16960 14980 17172 15008
rect 17034 14900 17040 14952
rect 17092 14900 17098 14952
rect 17144 14949 17172 14980
rect 17586 14968 17592 15020
rect 17644 15008 17650 15020
rect 17644 14980 20300 15008
rect 17644 14968 17650 14980
rect 17130 14943 17188 14949
rect 17130 14909 17142 14943
rect 17176 14909 17188 14943
rect 17130 14903 17188 14909
rect 17494 14900 17500 14952
rect 17552 14949 17558 14952
rect 17552 14903 17560 14949
rect 17552 14900 17558 14903
rect 15988 14844 16712 14872
rect 15988 14832 15994 14844
rect 17310 14832 17316 14884
rect 17368 14832 17374 14884
rect 17402 14832 17408 14884
rect 17460 14832 17466 14884
rect 17604 14804 17632 14968
rect 18414 14900 18420 14952
rect 18472 14900 18478 14952
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 18874 14949 18880 14952
rect 18841 14943 18880 14949
rect 18841 14909 18853 14943
rect 18841 14903 18880 14909
rect 18874 14900 18880 14903
rect 18932 14900 18938 14952
rect 19199 14943 19257 14949
rect 19199 14909 19211 14943
rect 19245 14940 19257 14943
rect 19306 14940 19334 14980
rect 19245 14912 19334 14940
rect 20073 14943 20131 14949
rect 19245 14909 19257 14912
rect 19199 14903 19257 14909
rect 20073 14909 20085 14943
rect 20119 14940 20131 14943
rect 20162 14940 20168 14952
rect 20119 14912 20168 14940
rect 20119 14909 20131 14912
rect 20073 14903 20131 14909
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 20272 14940 20300 14980
rect 20346 14968 20352 15020
rect 20404 14968 20410 15020
rect 22186 14940 22192 14952
rect 20272 14912 22192 14940
rect 22186 14900 22192 14912
rect 22244 14940 22250 14952
rect 22462 14940 22468 14952
rect 22244 14912 22468 14940
rect 22244 14900 22250 14912
rect 22462 14900 22468 14912
rect 22520 14940 22526 14952
rect 22848 14949 22876 15116
rect 24780 15076 24808 15116
rect 25222 15104 25228 15156
rect 25280 15104 25286 15156
rect 27249 15147 27307 15153
rect 27249 15144 27261 15147
rect 25332 15116 27261 15144
rect 25332 15076 25360 15116
rect 27249 15113 27261 15116
rect 27295 15113 27307 15147
rect 27249 15107 27307 15113
rect 27522 15104 27528 15156
rect 27580 15104 27586 15156
rect 24780 15048 25360 15076
rect 27157 15079 27215 15085
rect 27157 15045 27169 15079
rect 27203 15076 27215 15079
rect 27540 15076 27568 15104
rect 27203 15048 27568 15076
rect 27203 15045 27215 15048
rect 27157 15039 27215 15045
rect 23124 14980 23980 15008
rect 22741 14943 22799 14949
rect 22741 14940 22753 14943
rect 22520 14912 22753 14940
rect 22520 14900 22526 14912
rect 22741 14909 22753 14912
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 22833 14943 22891 14949
rect 22833 14909 22845 14943
rect 22879 14909 22891 14943
rect 22833 14903 22891 14909
rect 22922 14900 22928 14952
rect 22980 14900 22986 14952
rect 23124 14949 23152 14980
rect 23109 14943 23167 14949
rect 23109 14909 23121 14943
rect 23155 14909 23167 14943
rect 23109 14903 23167 14909
rect 23201 14943 23259 14949
rect 23201 14909 23213 14943
rect 23247 14909 23259 14943
rect 23845 14943 23903 14949
rect 23845 14940 23857 14943
rect 23201 14903 23259 14909
rect 23400 14912 23857 14940
rect 18432 14872 18460 14900
rect 18969 14875 19027 14881
rect 18969 14872 18981 14875
rect 18432 14844 18981 14872
rect 18969 14841 18981 14844
rect 19015 14841 19027 14875
rect 18969 14835 19027 14841
rect 19061 14875 19119 14881
rect 19061 14841 19073 14875
rect 19107 14872 19119 14875
rect 19702 14872 19708 14884
rect 19107 14844 19708 14872
rect 19107 14841 19119 14844
rect 19061 14835 19119 14841
rect 19702 14832 19708 14844
rect 19760 14832 19766 14884
rect 20594 14875 20652 14881
rect 20594 14872 20606 14875
rect 20272 14844 20606 14872
rect 20272 14813 20300 14844
rect 20594 14841 20606 14844
rect 20640 14841 20652 14875
rect 22094 14872 22100 14884
rect 20594 14835 20652 14841
rect 21652 14844 22100 14872
rect 15304 14776 17632 14804
rect 20257 14807 20315 14813
rect 20257 14773 20269 14807
rect 20303 14773 20315 14807
rect 20257 14767 20315 14773
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 21652 14804 21680 14844
rect 22094 14832 22100 14844
rect 22152 14872 22158 14884
rect 23216 14872 23244 14903
rect 22152 14844 23244 14872
rect 22152 14832 22158 14844
rect 20404 14776 21680 14804
rect 20404 14764 20410 14776
rect 21726 14764 21732 14816
rect 21784 14764 21790 14816
rect 22002 14764 22008 14816
rect 22060 14804 22066 14816
rect 22557 14807 22615 14813
rect 22557 14804 22569 14807
rect 22060 14776 22569 14804
rect 22060 14764 22066 14776
rect 22557 14773 22569 14776
rect 22603 14773 22615 14807
rect 22557 14767 22615 14773
rect 23290 14764 23296 14816
rect 23348 14804 23354 14816
rect 23400 14813 23428 14912
rect 23845 14909 23857 14912
rect 23891 14909 23903 14943
rect 23952 14940 23980 14980
rect 28626 14968 28632 15020
rect 28684 14968 28690 15020
rect 24486 14940 24492 14952
rect 23952 14912 24492 14940
rect 23845 14903 23903 14909
rect 24486 14900 24492 14912
rect 24544 14900 24550 14952
rect 25777 14943 25835 14949
rect 25777 14909 25789 14943
rect 25823 14940 25835 14943
rect 25866 14940 25872 14952
rect 25823 14912 25872 14940
rect 25823 14909 25835 14912
rect 25777 14903 25835 14909
rect 25866 14900 25872 14912
rect 25924 14900 25930 14952
rect 23474 14832 23480 14884
rect 23532 14872 23538 14884
rect 26050 14881 26056 14884
rect 24090 14875 24148 14881
rect 24090 14872 24102 14875
rect 23532 14844 24102 14872
rect 23532 14832 23538 14844
rect 24090 14841 24102 14844
rect 24136 14841 24148 14875
rect 24090 14835 24148 14841
rect 26044 14835 26056 14881
rect 26050 14832 26056 14835
rect 26108 14832 26114 14884
rect 28384 14875 28442 14881
rect 28384 14841 28396 14875
rect 28430 14872 28442 14875
rect 28718 14872 28724 14884
rect 28430 14844 28724 14872
rect 28430 14841 28442 14844
rect 28384 14835 28442 14841
rect 28718 14832 28724 14844
rect 28776 14832 28782 14884
rect 23385 14807 23443 14813
rect 23385 14804 23397 14807
rect 23348 14776 23397 14804
rect 23348 14764 23354 14776
rect 23385 14773 23397 14776
rect 23431 14773 23443 14807
rect 23385 14767 23443 14773
rect 552 14714 31808 14736
rect 552 14662 8172 14714
rect 8224 14662 8236 14714
rect 8288 14662 8300 14714
rect 8352 14662 8364 14714
rect 8416 14662 8428 14714
rect 8480 14662 15946 14714
rect 15998 14662 16010 14714
rect 16062 14662 16074 14714
rect 16126 14662 16138 14714
rect 16190 14662 16202 14714
rect 16254 14662 23720 14714
rect 23772 14662 23784 14714
rect 23836 14662 23848 14714
rect 23900 14662 23912 14714
rect 23964 14662 23976 14714
rect 24028 14662 31494 14714
rect 31546 14662 31558 14714
rect 31610 14662 31622 14714
rect 31674 14662 31686 14714
rect 31738 14662 31750 14714
rect 31802 14662 31808 14714
rect 552 14640 31808 14662
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3421 14603 3479 14609
rect 3108 14572 3372 14600
rect 3108 14560 3114 14572
rect 1302 14532 1308 14544
rect 1136 14504 1308 14532
rect 1136 14473 1164 14504
rect 1302 14492 1308 14504
rect 1360 14492 1366 14544
rect 3145 14535 3203 14541
rect 3145 14532 3157 14535
rect 2622 14504 3157 14532
rect 3145 14501 3157 14504
rect 3191 14501 3203 14535
rect 3344 14532 3372 14572
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 3602 14600 3608 14612
rect 3467 14572 3608 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4396 14572 4445 14600
rect 4396 14560 4402 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4433 14563 4491 14569
rect 4798 14560 4804 14612
rect 4856 14560 4862 14612
rect 7466 14560 7472 14612
rect 7524 14560 7530 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 8941 14603 8999 14609
rect 7616 14572 8892 14600
rect 7616 14560 7622 14572
rect 3344 14504 3832 14532
rect 3145 14495 3203 14501
rect 1121 14467 1179 14473
rect 1121 14433 1133 14467
rect 1167 14433 1179 14467
rect 1121 14427 1179 14433
rect 3237 14467 3295 14473
rect 3237 14433 3249 14467
rect 3283 14464 3295 14467
rect 3283 14436 3372 14464
rect 3283 14433 3295 14436
rect 3237 14427 3295 14433
rect 1394 14356 1400 14408
rect 1452 14356 1458 14408
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 3344 14328 3372 14436
rect 3418 14424 3424 14476
rect 3476 14464 3482 14476
rect 3804 14473 3832 14504
rect 3605 14467 3663 14473
rect 3605 14464 3617 14467
rect 3476 14436 3617 14464
rect 3476 14424 3482 14436
rect 3605 14433 3617 14436
rect 3651 14433 3663 14467
rect 3605 14427 3663 14433
rect 3789 14467 3847 14473
rect 3789 14433 3801 14467
rect 3835 14433 3847 14467
rect 3789 14427 3847 14433
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14464 4399 14467
rect 4816 14464 4844 14560
rect 7484 14532 7512 14560
rect 7806 14535 7864 14541
rect 7806 14532 7818 14535
rect 7484 14504 7818 14532
rect 7806 14501 7818 14504
rect 7852 14501 7864 14535
rect 7806 14495 7864 14501
rect 8662 14492 8668 14544
rect 8720 14492 8726 14544
rect 4387 14436 4844 14464
rect 4387 14433 4399 14436
rect 4341 14427 4399 14433
rect 3881 14399 3939 14405
rect 3881 14365 3893 14399
rect 3927 14396 3939 14399
rect 4154 14396 4160 14408
rect 3927 14368 4160 14396
rect 3927 14365 3939 14368
rect 3881 14359 3939 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4356 14328 4384 14427
rect 5442 14424 5448 14476
rect 5500 14464 5506 14476
rect 6086 14473 6092 14476
rect 5813 14467 5871 14473
rect 5813 14464 5825 14467
rect 5500 14436 5825 14464
rect 5500 14424 5506 14436
rect 5813 14433 5825 14436
rect 5859 14433 5871 14467
rect 5813 14427 5871 14433
rect 6080 14427 6092 14473
rect 6086 14424 6092 14427
rect 6144 14424 6150 14476
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14464 7619 14467
rect 7650 14464 7656 14476
rect 7607 14436 7656 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 8680 14396 8708 14492
rect 8864 14464 8892 14572
rect 8941 14569 8953 14603
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 9401 14603 9459 14609
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 10226 14600 10232 14612
rect 9447 14572 10232 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 8956 14532 8984 14563
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 12989 14603 13047 14609
rect 12989 14569 13001 14603
rect 13035 14600 13047 14603
rect 13538 14600 13544 14612
rect 13035 14572 13544 14600
rect 13035 14569 13047 14572
rect 12989 14563 13047 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 14182 14600 14188 14612
rect 13679 14572 14188 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 14277 14603 14335 14609
rect 14277 14569 14289 14603
rect 14323 14600 14335 14603
rect 15102 14600 15108 14612
rect 14323 14572 15108 14600
rect 14323 14569 14335 14572
rect 14277 14563 14335 14569
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15657 14603 15715 14609
rect 15657 14569 15669 14603
rect 15703 14600 15715 14603
rect 15703 14572 16160 14600
rect 15703 14569 15715 14572
rect 15657 14563 15715 14569
rect 11330 14532 11336 14544
rect 8956 14504 11336 14532
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 11514 14492 11520 14544
rect 11572 14532 11578 14544
rect 13357 14535 13415 14541
rect 13357 14532 13369 14535
rect 11572 14504 13369 14532
rect 11572 14492 11578 14504
rect 13357 14501 13369 14504
rect 13403 14501 13415 14535
rect 13357 14495 13415 14501
rect 13464 14504 13860 14532
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 8864 14436 9229 14464
rect 9217 14433 9229 14436
rect 9263 14464 9275 14467
rect 9398 14464 9404 14476
rect 9263 14436 9404 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 9398 14424 9404 14436
rect 9456 14424 9462 14476
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14464 9551 14467
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 9539 14436 9873 14464
rect 9539 14433 9551 14436
rect 9493 14427 9551 14433
rect 9861 14433 9873 14436
rect 9907 14433 9919 14467
rect 9861 14427 9919 14433
rect 9508 14396 9536 14427
rect 8680 14368 9536 14396
rect 9766 14356 9772 14408
rect 9824 14356 9830 14408
rect 9876 14396 9904 14427
rect 10502 14424 10508 14476
rect 10560 14424 10566 14476
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10735 14436 10824 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 10137 14399 10195 14405
rect 9876 14368 10088 14396
rect 3292 14300 4384 14328
rect 3292 14288 3298 14300
rect 7190 14288 7196 14340
rect 7248 14288 7254 14340
rect 9214 14288 9220 14340
rect 9272 14328 9278 14340
rect 9585 14331 9643 14337
rect 9585 14328 9597 14331
rect 9272 14300 9597 14328
rect 9272 14288 9278 14300
rect 9585 14297 9597 14300
rect 9631 14328 9643 14331
rect 9861 14331 9919 14337
rect 9861 14328 9873 14331
rect 9631 14300 9873 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 9861 14297 9873 14300
rect 9907 14297 9919 14331
rect 9861 14291 9919 14297
rect 9953 14331 10011 14337
rect 9953 14297 9965 14331
rect 9999 14297 10011 14331
rect 10060 14328 10088 14368
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 10597 14399 10655 14405
rect 10597 14396 10609 14399
rect 10183 14368 10609 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10597 14365 10609 14368
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 10796 14340 10824 14436
rect 10888 14436 11161 14464
rect 10410 14328 10416 14340
rect 10060 14300 10416 14328
rect 9953 14291 10011 14297
rect 1026 14220 1032 14272
rect 1084 14260 1090 14272
rect 2038 14260 2044 14272
rect 1084 14232 2044 14260
rect 1084 14220 1090 14232
rect 2038 14220 2044 14232
rect 2096 14260 2102 14272
rect 2866 14260 2872 14272
rect 2096 14232 2872 14260
rect 2096 14220 2102 14232
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 9398 14220 9404 14272
rect 9456 14260 9462 14272
rect 9493 14263 9551 14269
rect 9493 14260 9505 14263
rect 9456 14232 9505 14260
rect 9456 14220 9462 14232
rect 9493 14229 9505 14232
rect 9539 14260 9551 14263
rect 9968 14260 9996 14291
rect 10410 14288 10416 14300
rect 10468 14288 10474 14340
rect 10778 14288 10784 14340
rect 10836 14288 10842 14340
rect 9539 14232 9996 14260
rect 9539 14229 9551 14232
rect 9493 14223 9551 14229
rect 10226 14220 10232 14272
rect 10284 14220 10290 14272
rect 10318 14220 10324 14272
rect 10376 14260 10382 14272
rect 10888 14260 10916 14436
rect 11149 14433 11161 14436
rect 11195 14464 11207 14467
rect 11238 14464 11244 14476
rect 11195 14436 11244 14464
rect 11195 14433 11207 14436
rect 11149 14427 11207 14433
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 11440 14396 11468 14427
rect 11606 14424 11612 14476
rect 11664 14424 11670 14476
rect 12434 14424 12440 14476
rect 12492 14424 12498 14476
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 12621 14467 12679 14473
rect 12621 14464 12633 14467
rect 12584 14436 12633 14464
rect 12584 14424 12590 14436
rect 12621 14433 12633 14436
rect 12667 14433 12679 14467
rect 12621 14427 12679 14433
rect 12710 14424 12716 14476
rect 12768 14424 12774 14476
rect 12802 14424 12808 14476
rect 12860 14424 12866 14476
rect 13464 14473 13492 14504
rect 13832 14476 13860 14504
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 15838 14532 15844 14544
rect 14424 14504 15844 14532
rect 14424 14492 14430 14504
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 16132 14532 16160 14572
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 17497 14603 17555 14609
rect 17497 14600 17509 14603
rect 17460 14572 17509 14600
rect 17460 14560 17466 14572
rect 17497 14569 17509 14572
rect 17543 14569 17555 14603
rect 17497 14563 17555 14569
rect 19153 14603 19211 14609
rect 19153 14569 19165 14603
rect 19199 14569 19211 14603
rect 19153 14563 19211 14569
rect 16362 14535 16420 14541
rect 16362 14532 16374 14535
rect 16132 14504 16374 14532
rect 16362 14501 16374 14504
rect 16408 14501 16420 14535
rect 19168 14532 19196 14563
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 21269 14603 21327 14609
rect 21269 14600 21281 14603
rect 20772 14572 21281 14600
rect 20772 14560 20778 14572
rect 21269 14569 21281 14572
rect 21315 14569 21327 14603
rect 21269 14563 21327 14569
rect 21726 14560 21732 14612
rect 21784 14600 21790 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21784 14572 21925 14600
rect 21784 14560 21790 14572
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 21913 14563 21971 14569
rect 22002 14560 22008 14612
rect 22060 14560 22066 14612
rect 22097 14603 22155 14609
rect 22097 14569 22109 14603
rect 22143 14600 22155 14603
rect 22278 14600 22284 14612
rect 22143 14572 22284 14600
rect 22143 14569 22155 14572
rect 22097 14563 22155 14569
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 24118 14560 24124 14612
rect 24176 14600 24182 14612
rect 24305 14603 24363 14609
rect 24305 14600 24317 14603
rect 24176 14572 24317 14600
rect 24176 14560 24182 14572
rect 24305 14569 24317 14572
rect 24351 14569 24363 14603
rect 24305 14563 24363 14569
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 25958 14600 25964 14612
rect 24912 14572 25964 14600
rect 24912 14560 24918 14572
rect 25958 14560 25964 14572
rect 26016 14560 26022 14612
rect 31297 14603 31355 14609
rect 31297 14600 31309 14603
rect 26059 14572 31309 14600
rect 19490 14535 19548 14541
rect 19490 14532 19502 14535
rect 19168 14504 19502 14532
rect 16362 14495 16420 14501
rect 19490 14501 19502 14504
rect 19536 14501 19548 14535
rect 22020 14532 22048 14560
rect 19490 14495 19548 14501
rect 21836 14504 22048 14532
rect 22373 14535 22431 14541
rect 13081 14467 13139 14473
rect 13081 14433 13093 14467
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 13265 14467 13323 14473
rect 13265 14433 13277 14467
rect 13311 14433 13323 14467
rect 13265 14427 13323 14433
rect 13449 14467 13507 14473
rect 13449 14433 13461 14467
rect 13495 14433 13507 14467
rect 13449 14427 13507 14433
rect 11020 14368 11468 14396
rect 11020 14356 11026 14368
rect 11514 14356 11520 14408
rect 11572 14396 11578 14408
rect 13096 14396 13124 14427
rect 11572 14368 13124 14396
rect 13280 14396 13308 14427
rect 13722 14424 13728 14476
rect 13780 14424 13786 14476
rect 13814 14424 13820 14476
rect 13872 14424 13878 14476
rect 13909 14467 13967 14473
rect 13909 14433 13921 14467
rect 13955 14433 13967 14467
rect 13909 14427 13967 14433
rect 13924 14396 13952 14427
rect 13998 14424 14004 14476
rect 14056 14424 14062 14476
rect 14090 14424 14096 14476
rect 14148 14424 14154 14476
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 14240 14436 15485 14464
rect 14240 14424 14246 14436
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 16206 14464 16212 14476
rect 16163 14436 16212 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 13280 14368 13952 14396
rect 14108 14396 14136 14424
rect 14826 14396 14832 14408
rect 14108 14368 14832 14396
rect 11572 14356 11578 14368
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 11425 14331 11483 14337
rect 11425 14328 11437 14331
rect 11112 14300 11437 14328
rect 11112 14288 11118 14300
rect 11425 14297 11437 14300
rect 11471 14297 11483 14331
rect 11425 14291 11483 14297
rect 10376 14232 10916 14260
rect 10376 14220 10382 14232
rect 11330 14220 11336 14272
rect 11388 14220 11394 14272
rect 12526 14220 12532 14272
rect 12584 14260 12590 14272
rect 13280 14260 13308 14368
rect 12584 14232 13308 14260
rect 13924 14260 13952 14368
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 16132 14396 16160 14427
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 18969 14467 19027 14473
rect 18969 14433 18981 14467
rect 19015 14464 19027 14467
rect 19150 14464 19156 14476
rect 19015 14436 19156 14464
rect 19015 14433 19027 14436
rect 18969 14427 19027 14433
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 19245 14467 19303 14473
rect 19245 14433 19257 14467
rect 19291 14464 19303 14467
rect 19291 14436 20300 14464
rect 19291 14433 19303 14436
rect 19245 14427 19303 14433
rect 14936 14368 16160 14396
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 14936 14328 14964 14368
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 18782 14396 18788 14408
rect 17644 14368 18788 14396
rect 17644 14356 17650 14368
rect 18782 14356 18788 14368
rect 18840 14396 18846 14408
rect 19260 14396 19288 14427
rect 18840 14368 19288 14396
rect 18840 14356 18846 14368
rect 14700 14300 14964 14328
rect 14700 14288 14706 14300
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 15746 14328 15752 14340
rect 15528 14300 15752 14328
rect 15528 14288 15534 14300
rect 15746 14288 15752 14300
rect 15804 14288 15810 14340
rect 20272 14328 20300 14436
rect 21266 14424 21272 14476
rect 21324 14464 21330 14476
rect 21637 14467 21695 14473
rect 21637 14464 21649 14467
rect 21324 14436 21649 14464
rect 21324 14424 21330 14436
rect 21637 14433 21649 14436
rect 21683 14433 21695 14467
rect 21637 14427 21695 14433
rect 21545 14399 21603 14405
rect 21545 14365 21557 14399
rect 21591 14396 21603 14399
rect 21836 14396 21864 14504
rect 22373 14501 22385 14535
rect 22419 14532 22431 14535
rect 26059 14532 26087 14572
rect 31297 14569 31309 14572
rect 31343 14569 31355 14603
rect 31297 14563 31355 14569
rect 22419 14504 26087 14532
rect 22419 14501 22431 14504
rect 22373 14495 22431 14501
rect 28810 14492 28816 14544
rect 28868 14492 28874 14544
rect 29086 14492 29092 14544
rect 29144 14492 29150 14544
rect 30162 14535 30220 14541
rect 30162 14532 30174 14535
rect 29196 14504 30174 14532
rect 29196 14476 29224 14504
rect 30162 14501 30174 14504
rect 30208 14501 30220 14535
rect 30162 14495 30220 14501
rect 22005 14467 22063 14473
rect 22005 14433 22017 14467
rect 22051 14433 22063 14467
rect 22005 14427 22063 14433
rect 21591 14368 21864 14396
rect 22020 14396 22048 14427
rect 22186 14424 22192 14476
rect 22244 14464 22250 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22244 14436 22293 14464
rect 22244 14424 22250 14436
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 22465 14467 22523 14473
rect 22465 14433 22477 14467
rect 22511 14464 22523 14467
rect 22554 14464 22560 14476
rect 22511 14436 22560 14464
rect 22511 14433 22523 14436
rect 22465 14427 22523 14433
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 22646 14424 22652 14476
rect 22704 14424 22710 14476
rect 24026 14424 24032 14476
rect 24084 14464 24090 14476
rect 25429 14467 25487 14473
rect 25429 14464 25441 14467
rect 24084 14436 25441 14464
rect 24084 14424 24090 14436
rect 25429 14433 25441 14436
rect 25475 14464 25487 14467
rect 26602 14464 26608 14476
rect 25475 14436 26608 14464
rect 25475 14433 25487 14436
rect 25429 14427 25487 14433
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 28626 14424 28632 14476
rect 28684 14424 28690 14476
rect 28718 14424 28724 14476
rect 28776 14464 28782 14476
rect 28997 14467 29055 14473
rect 28997 14464 29009 14467
rect 28776 14436 29009 14464
rect 28776 14424 28782 14436
rect 28997 14433 29009 14436
rect 29043 14433 29055 14467
rect 28997 14427 29055 14433
rect 29178 14424 29184 14476
rect 29236 14424 29242 14476
rect 29365 14467 29423 14473
rect 29365 14433 29377 14467
rect 29411 14464 29423 14467
rect 29641 14467 29699 14473
rect 29641 14464 29653 14467
rect 29411 14436 29653 14464
rect 29411 14433 29423 14436
rect 29365 14427 29423 14433
rect 29641 14433 29653 14436
rect 29687 14433 29699 14467
rect 29641 14427 29699 14433
rect 23382 14396 23388 14408
rect 22020 14368 23388 14396
rect 21591 14365 21603 14368
rect 21545 14359 21603 14365
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 25685 14399 25743 14405
rect 25685 14365 25697 14399
rect 25731 14396 25743 14399
rect 25866 14396 25872 14408
rect 25731 14368 25872 14396
rect 25731 14365 25743 14368
rect 25685 14359 25743 14365
rect 25866 14356 25872 14368
rect 25924 14356 25930 14408
rect 25958 14356 25964 14408
rect 26016 14396 26022 14408
rect 26697 14399 26755 14405
rect 26697 14396 26709 14399
rect 26016 14368 26709 14396
rect 26016 14356 26022 14368
rect 26697 14365 26709 14368
rect 26743 14396 26755 14399
rect 26743 14368 28120 14396
rect 26743 14365 26755 14368
rect 26697 14359 26755 14365
rect 23290 14328 23296 14340
rect 20272 14300 23296 14328
rect 23290 14288 23296 14300
rect 23348 14288 23354 14340
rect 18414 14260 18420 14272
rect 13924 14232 18420 14260
rect 12584 14220 12590 14232
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 20622 14220 20628 14272
rect 20680 14220 20686 14272
rect 21726 14220 21732 14272
rect 21784 14220 21790 14272
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 26786 14260 26792 14272
rect 24360 14232 26792 14260
rect 24360 14220 24366 14232
rect 26786 14220 26792 14232
rect 26844 14220 26850 14272
rect 26973 14263 27031 14269
rect 26973 14229 26985 14263
rect 27019 14260 27031 14263
rect 27982 14260 27988 14272
rect 27019 14232 27988 14260
rect 27019 14229 27031 14232
rect 26973 14223 27031 14229
rect 27982 14220 27988 14232
rect 28040 14220 28046 14272
rect 28092 14260 28120 14368
rect 28644 14328 28672 14424
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14365 29975 14399
rect 29917 14359 29975 14365
rect 29932 14328 29960 14359
rect 28644 14300 29960 14328
rect 28626 14260 28632 14272
rect 28092 14232 28632 14260
rect 28626 14220 28632 14232
rect 28684 14260 28690 14272
rect 29549 14263 29607 14269
rect 29549 14260 29561 14263
rect 28684 14232 29561 14260
rect 28684 14220 28690 14232
rect 29549 14229 29561 14232
rect 29595 14229 29607 14263
rect 29549 14223 29607 14229
rect 552 14170 31648 14192
rect 552 14118 4285 14170
rect 4337 14118 4349 14170
rect 4401 14118 4413 14170
rect 4465 14118 4477 14170
rect 4529 14118 4541 14170
rect 4593 14118 12059 14170
rect 12111 14118 12123 14170
rect 12175 14118 12187 14170
rect 12239 14118 12251 14170
rect 12303 14118 12315 14170
rect 12367 14118 19833 14170
rect 19885 14118 19897 14170
rect 19949 14118 19961 14170
rect 20013 14118 20025 14170
rect 20077 14118 20089 14170
rect 20141 14118 27607 14170
rect 27659 14118 27671 14170
rect 27723 14118 27735 14170
rect 27787 14118 27799 14170
rect 27851 14118 27863 14170
rect 27915 14118 31648 14170
rect 552 14096 31648 14118
rect 1394 14016 1400 14068
rect 1452 14016 1458 14068
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 7800 14028 8401 14056
rect 7800 14016 7806 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 9490 14016 9496 14068
rect 9548 14016 9554 14068
rect 9766 14016 9772 14068
rect 9824 14016 9830 14068
rect 10226 14016 10232 14068
rect 10284 14016 10290 14068
rect 10410 14016 10416 14068
rect 10468 14056 10474 14068
rect 10468 14028 10640 14056
rect 10468 14016 10474 14028
rect 1302 13948 1308 14000
rect 1360 13988 1366 14000
rect 3326 13988 3332 14000
rect 1360 13960 3332 13988
rect 1360 13948 1366 13960
rect 3326 13948 3332 13960
rect 3384 13948 3390 14000
rect 4154 13948 4160 14000
rect 4212 13948 4218 14000
rect 7009 13991 7067 13997
rect 7009 13957 7021 13991
rect 7055 13988 7067 13991
rect 9508 13988 9536 14016
rect 10244 13988 10272 14016
rect 7055 13960 9536 13988
rect 9784 13960 10272 13988
rect 7055 13957 7067 13960
rect 7009 13951 7067 13957
rect 1121 13923 1179 13929
rect 1121 13889 1133 13923
rect 1167 13920 1179 13923
rect 1670 13920 1676 13932
rect 1167 13892 1676 13920
rect 1167 13889 1179 13892
rect 1121 13883 1179 13889
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 4172 13920 4200 13948
rect 3988 13892 5304 13920
rect 1026 13812 1032 13864
rect 1084 13812 1090 13864
rect 3988 13861 4016 13892
rect 5276 13864 5304 13892
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5500 13892 5641 13920
rect 5500 13880 5506 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 4154 13812 4160 13864
rect 4212 13812 4218 13864
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 5166 13852 5172 13864
rect 4295 13824 5172 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 5644 13852 5672 13883
rect 6454 13852 6460 13864
rect 5644 13824 6460 13852
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 9784 13861 9812 13960
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 10275 13892 10425 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10413 13889 10425 13892
rect 10459 13889 10471 13923
rect 10612 13920 10640 14028
rect 11054 14016 11060 14068
rect 11112 14016 11118 14068
rect 11330 14016 11336 14068
rect 11388 14016 11394 14068
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 11664 14028 12434 14056
rect 11664 14016 11670 14028
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 10873 13991 10931 13997
rect 10873 13988 10885 13991
rect 10744 13960 10885 13988
rect 10744 13948 10750 13960
rect 10873 13957 10885 13960
rect 10919 13957 10931 13991
rect 10873 13951 10931 13957
rect 11072 13929 11100 14016
rect 11057 13923 11115 13929
rect 10612 13892 10732 13920
rect 10413 13883 10471 13889
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 9769 13855 9827 13861
rect 9631 13824 9720 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 5902 13793 5908 13796
rect 5896 13747 5908 13793
rect 5902 13744 5908 13747
rect 5960 13744 5966 13796
rect 3786 13676 3792 13728
rect 3844 13676 3850 13728
rect 9692 13716 9720 13824
rect 9769 13821 9781 13855
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10137 13855 10195 13861
rect 10137 13852 10149 13855
rect 10091 13824 10149 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10137 13821 10149 13824
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 10318 13812 10324 13864
rect 10376 13812 10382 13864
rect 10704 13861 10732 13892
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11348 13920 11376 14016
rect 12406 13988 12434 14028
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 14182 14016 14188 14068
rect 14240 14016 14246 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 17126 14056 17132 14068
rect 16071 14028 17132 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 18233 14059 18291 14065
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 18322 14056 18328 14068
rect 18279 14028 18328 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 20622 14016 20628 14068
rect 20680 14016 20686 14068
rect 21177 14059 21235 14065
rect 21177 14025 21189 14059
rect 21223 14056 21235 14059
rect 21726 14056 21732 14068
rect 21223 14028 21732 14056
rect 21223 14025 21235 14028
rect 21177 14019 21235 14025
rect 21726 14016 21732 14028
rect 21784 14016 21790 14068
rect 23566 14016 23572 14068
rect 23624 14016 23630 14068
rect 24213 14059 24271 14065
rect 24213 14025 24225 14059
rect 24259 14056 24271 14059
rect 25038 14056 25044 14068
rect 24259 14028 25044 14056
rect 24259 14025 24271 14028
rect 24213 14019 24271 14025
rect 25038 14016 25044 14028
rect 25096 14016 25102 14068
rect 26050 14016 26056 14068
rect 26108 14016 26114 14068
rect 26786 14016 26792 14068
rect 26844 14056 26850 14068
rect 28074 14056 28080 14068
rect 26844 14028 28080 14056
rect 26844 14016 26850 14028
rect 28074 14016 28080 14028
rect 28132 14016 28138 14068
rect 28629 14059 28687 14065
rect 28629 14025 28641 14059
rect 28675 14056 28687 14059
rect 28718 14056 28724 14068
rect 28675 14028 28724 14056
rect 28675 14025 28687 14028
rect 28629 14019 28687 14025
rect 28718 14016 28724 14028
rect 28776 14016 28782 14068
rect 14200 13988 14228 14016
rect 12406 13960 14228 13988
rect 14369 13991 14427 13997
rect 14369 13957 14381 13991
rect 14415 13957 14427 13991
rect 14369 13951 14427 13957
rect 14384 13920 14412 13951
rect 20640 13920 20668 14016
rect 11348 13892 11468 13920
rect 14384 13892 14780 13920
rect 20640 13892 20944 13920
rect 11057 13883 11115 13889
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10735 13824 10793 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 10612 13784 10640 13815
rect 11330 13812 11336 13864
rect 11388 13812 11394 13864
rect 11440 13852 11468 13892
rect 11589 13855 11647 13861
rect 11589 13852 11601 13855
rect 11440 13824 11601 13852
rect 11589 13821 11601 13824
rect 11635 13821 11647 13855
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 11589 13815 11647 13821
rect 11716 13824 14197 13852
rect 10612 13756 10824 13784
rect 10796 13728 10824 13756
rect 10686 13716 10692 13728
rect 9692 13688 10692 13716
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 11716 13716 11744 13824
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 14642 13812 14648 13864
rect 14700 13812 14706 13864
rect 14752 13852 14780 13892
rect 14901 13855 14959 13861
rect 14901 13852 14913 13855
rect 14752 13824 14913 13852
rect 14901 13821 14913 13824
rect 14947 13821 14959 13855
rect 14901 13815 14959 13821
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13852 16911 13855
rect 17586 13852 17592 13864
rect 16899 13824 17592 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 20622 13812 20628 13864
rect 20680 13812 20686 13864
rect 20916 13861 20944 13892
rect 22094 13880 22100 13932
rect 22152 13920 22158 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 22152 13892 22201 13920
rect 22152 13880 22158 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 24581 13923 24639 13929
rect 24581 13889 24593 13923
rect 24627 13920 24639 13923
rect 25222 13920 25228 13932
rect 24627 13892 25228 13920
rect 24627 13889 24639 13892
rect 24581 13883 24639 13889
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 20901 13855 20959 13861
rect 20901 13821 20913 13855
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 20990 13812 20996 13864
rect 21048 13812 21054 13864
rect 23937 13855 23995 13861
rect 23937 13821 23949 13855
rect 23983 13821 23995 13855
rect 23937 13815 23995 13821
rect 17120 13787 17178 13793
rect 17120 13753 17132 13787
rect 17166 13784 17178 13787
rect 17678 13784 17684 13796
rect 17166 13756 17684 13784
rect 17166 13753 17178 13756
rect 17120 13747 17178 13753
rect 17678 13744 17684 13756
rect 17736 13744 17742 13796
rect 18414 13744 18420 13796
rect 18472 13784 18478 13796
rect 20809 13787 20867 13793
rect 20809 13784 20821 13787
rect 18472 13756 20821 13784
rect 18472 13744 18478 13756
rect 20809 13753 20821 13756
rect 20855 13753 20867 13787
rect 20809 13747 20867 13753
rect 10836 13688 11744 13716
rect 20824 13716 20852 13747
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22434 13787 22492 13793
rect 22434 13784 22446 13787
rect 22152 13756 22446 13784
rect 22152 13744 22158 13756
rect 22434 13753 22446 13756
rect 22480 13753 22492 13787
rect 22434 13747 22492 13753
rect 22554 13744 22560 13796
rect 22612 13744 22618 13796
rect 22572 13716 22600 13744
rect 20824 13688 22600 13716
rect 23952 13716 23980 13815
rect 24026 13812 24032 13864
rect 24084 13812 24090 13864
rect 24213 13855 24271 13861
rect 24213 13821 24225 13855
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 24228 13784 24256 13815
rect 24302 13812 24308 13864
rect 24360 13812 24366 13864
rect 26234 13812 26240 13864
rect 26292 13852 26298 13864
rect 26697 13855 26755 13861
rect 26697 13852 26709 13855
rect 26292 13824 26709 13852
rect 26292 13812 26298 13824
rect 26697 13821 26709 13824
rect 26743 13821 26755 13855
rect 28092 13852 28120 14016
rect 28813 13991 28871 13997
rect 28813 13957 28825 13991
rect 28859 13988 28871 13991
rect 28994 13988 29000 14000
rect 28859 13960 29000 13988
rect 28859 13957 28871 13960
rect 28813 13951 28871 13957
rect 28994 13948 29000 13960
rect 29052 13948 29058 14000
rect 29181 13855 29239 13861
rect 29181 13852 29193 13855
rect 28092 13824 29193 13852
rect 26697 13815 26755 13821
rect 29181 13821 29193 13824
rect 29227 13821 29239 13855
rect 29181 13815 29239 13821
rect 24228 13756 24992 13784
rect 24964 13728 24992 13756
rect 25590 13744 25596 13796
rect 25648 13744 25654 13796
rect 28445 13787 28503 13793
rect 28445 13753 28457 13787
rect 28491 13784 28503 13787
rect 28810 13784 28816 13796
rect 28491 13756 28816 13784
rect 28491 13753 28503 13756
rect 28445 13747 28503 13753
rect 28810 13744 28816 13756
rect 28868 13744 28874 13796
rect 29454 13744 29460 13796
rect 29512 13744 29518 13796
rect 30190 13744 30196 13796
rect 30248 13744 30254 13796
rect 24394 13716 24400 13728
rect 23952 13688 24400 13716
rect 10836 13676 10842 13688
rect 24394 13676 24400 13688
rect 24452 13676 24458 13728
rect 24946 13676 24952 13728
rect 25004 13676 25010 13728
rect 28655 13719 28713 13725
rect 28655 13685 28667 13719
rect 28701 13716 28713 13719
rect 29086 13716 29092 13728
rect 28701 13688 29092 13716
rect 28701 13685 28713 13688
rect 28655 13679 28713 13685
rect 29086 13676 29092 13688
rect 29144 13716 29150 13728
rect 30929 13719 30987 13725
rect 30929 13716 30941 13719
rect 29144 13688 30941 13716
rect 29144 13676 29150 13688
rect 30929 13685 30941 13688
rect 30975 13685 30987 13719
rect 30929 13679 30987 13685
rect 552 13626 31808 13648
rect 552 13574 8172 13626
rect 8224 13574 8236 13626
rect 8288 13574 8300 13626
rect 8352 13574 8364 13626
rect 8416 13574 8428 13626
rect 8480 13574 15946 13626
rect 15998 13574 16010 13626
rect 16062 13574 16074 13626
rect 16126 13574 16138 13626
rect 16190 13574 16202 13626
rect 16254 13574 23720 13626
rect 23772 13574 23784 13626
rect 23836 13574 23848 13626
rect 23900 13574 23912 13626
rect 23964 13574 23976 13626
rect 24028 13574 31494 13626
rect 31546 13574 31558 13626
rect 31610 13574 31622 13626
rect 31674 13574 31686 13626
rect 31738 13574 31750 13626
rect 31802 13574 31808 13626
rect 552 13552 31808 13574
rect 3234 13472 3240 13524
rect 3292 13472 3298 13524
rect 5166 13472 5172 13524
rect 5224 13512 5230 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5224 13484 6009 13512
rect 5224 13472 5230 13484
rect 5997 13481 6009 13484
rect 6043 13512 6055 13515
rect 6086 13512 6092 13524
rect 6043 13484 6092 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13481 7987 13515
rect 7929 13475 7987 13481
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11287 13484 12434 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 1302 13444 1308 13456
rect 1136 13416 1308 13444
rect 1136 13385 1164 13416
rect 1302 13404 1308 13416
rect 1360 13404 1366 13456
rect 3053 13447 3111 13453
rect 3053 13444 3065 13447
rect 2622 13416 3065 13444
rect 3053 13413 3065 13416
rect 3099 13413 3111 13447
rect 3053 13407 3111 13413
rect 1121 13379 1179 13385
rect 1121 13345 1133 13379
rect 1167 13345 1179 13379
rect 1121 13339 1179 13345
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13376 3203 13379
rect 3252 13376 3280 13472
rect 3697 13447 3755 13453
rect 3697 13413 3709 13447
rect 3743 13444 3755 13447
rect 3786 13444 3792 13456
rect 3743 13416 3792 13444
rect 3743 13413 3755 13416
rect 3697 13407 3755 13413
rect 3786 13404 3792 13416
rect 3844 13404 3850 13456
rect 4706 13404 4712 13456
rect 4764 13404 4770 13456
rect 6181 13447 6239 13453
rect 6181 13444 6193 13447
rect 5552 13416 6193 13444
rect 5552 13388 5580 13416
rect 6181 13413 6193 13416
rect 6227 13444 6239 13447
rect 7944 13444 7972 13475
rect 12406 13444 12434 13484
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 14056 13484 14105 13512
rect 14056 13472 14062 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 15562 13472 15568 13524
rect 15620 13472 15626 13524
rect 18874 13472 18880 13524
rect 18932 13472 18938 13524
rect 19702 13472 19708 13524
rect 19760 13512 19766 13524
rect 21913 13515 21971 13521
rect 21913 13512 21925 13515
rect 19760 13484 21925 13512
rect 19760 13472 19766 13484
rect 21913 13481 21925 13484
rect 21959 13481 21971 13515
rect 25130 13512 25136 13524
rect 21913 13475 21971 13481
rect 22296 13484 25136 13512
rect 14430 13447 14488 13453
rect 14430 13444 14442 13447
rect 6227 13416 6960 13444
rect 7944 13416 11468 13444
rect 12406 13416 14442 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 3191 13348 3280 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 5534 13336 5540 13388
rect 5592 13336 5598 13388
rect 5626 13336 5632 13388
rect 5684 13376 5690 13388
rect 5902 13376 5908 13388
rect 5684 13348 5908 13376
rect 5684 13336 5690 13348
rect 5902 13336 5908 13348
rect 5960 13376 5966 13388
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5960 13348 6101 13376
rect 5960 13336 5966 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6805 13379 6863 13385
rect 6805 13376 6817 13379
rect 6089 13339 6147 13345
rect 6380 13348 6817 13376
rect 1394 13268 1400 13320
rect 1452 13268 1458 13320
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 3384 13280 3433 13308
rect 3384 13268 3390 13280
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 6270 13200 6276 13252
rect 6328 13240 6334 13252
rect 6380 13249 6408 13348
rect 6805 13345 6817 13348
rect 6851 13345 6863 13379
rect 6932 13376 6960 13416
rect 8277 13379 8335 13385
rect 8277 13376 8289 13379
rect 6932 13348 8289 13376
rect 6805 13339 6863 13345
rect 8277 13345 8289 13348
rect 8323 13345 8335 13379
rect 8277 13339 8335 13345
rect 10686 13336 10692 13388
rect 10744 13376 10750 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10744 13348 11069 13376
rect 10744 13336 10750 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6512 13280 6561 13308
rect 6512 13268 6518 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 6365 13243 6423 13249
rect 6365 13240 6377 13243
rect 6328 13212 6377 13240
rect 6328 13200 6334 13212
rect 6365 13209 6377 13212
rect 6411 13209 6423 13243
rect 6365 13203 6423 13209
rect 2866 13132 2872 13184
rect 2924 13132 2930 13184
rect 5810 13132 5816 13184
rect 5868 13132 5874 13184
rect 6564 13172 6592 13271
rect 8036 13172 8064 13271
rect 11440 13240 11468 13416
rect 14430 13413 14442 13416
rect 14476 13413 14488 13447
rect 14430 13407 14488 13413
rect 14642 13404 14648 13456
rect 14700 13404 14706 13456
rect 17764 13447 17822 13453
rect 17764 13413 17776 13447
rect 17810 13444 17822 13447
rect 17954 13444 17960 13456
rect 17810 13416 17960 13444
rect 17810 13413 17822 13416
rect 17764 13407 17822 13413
rect 17954 13404 17960 13416
rect 18012 13404 18018 13456
rect 19058 13404 19064 13456
rect 19116 13444 19122 13456
rect 19116 13416 21496 13444
rect 19116 13404 19122 13416
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 12618 13376 12624 13388
rect 11664 13348 12624 13376
rect 11664 13336 11670 13348
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 12980 13379 13038 13385
rect 12980 13345 12992 13379
rect 13026 13376 13038 13379
rect 13354 13376 13360 13388
rect 13026 13348 13360 13376
rect 13026 13345 13038 13348
rect 12980 13339 13038 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 14185 13379 14243 13385
rect 14185 13345 14197 13379
rect 14231 13376 14243 13379
rect 14660 13376 14688 13404
rect 15010 13376 15016 13388
rect 14231 13348 15016 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 15010 13336 15016 13348
rect 15068 13336 15074 13388
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13376 17555 13379
rect 17586 13376 17592 13388
rect 17543 13348 17592 13376
rect 17543 13345 17555 13348
rect 17497 13339 17555 13345
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 21468 13385 21496 13416
rect 19521 13379 19579 13385
rect 19521 13345 19533 13379
rect 19567 13376 19579 13379
rect 21453 13379 21511 13385
rect 19567 13348 20852 13376
rect 19567 13345 19579 13348
rect 19521 13339 19579 13345
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 20824 13308 20852 13348
rect 21453 13345 21465 13379
rect 21499 13345 21511 13379
rect 21453 13339 21511 13345
rect 22094 13308 22100 13320
rect 20824 13280 22100 13308
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 12434 13240 12440 13252
rect 9416 13212 11376 13240
rect 11440 13212 12440 13240
rect 8294 13172 8300 13184
rect 6564 13144 8300 13172
rect 8294 13132 8300 13144
rect 8352 13172 8358 13184
rect 9306 13172 9312 13184
rect 8352 13144 9312 13172
rect 8352 13132 8358 13144
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9416 13181 9444 13212
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13141 9459 13175
rect 11348 13172 11376 13212
rect 12434 13200 12440 13212
rect 12492 13200 12498 13252
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 22296 13240 22324 13484
rect 25130 13472 25136 13484
rect 25188 13472 25194 13524
rect 25222 13472 25228 13524
rect 25280 13512 25286 13524
rect 25317 13515 25375 13521
rect 25317 13512 25329 13515
rect 25280 13484 25329 13512
rect 25280 13472 25286 13484
rect 25317 13481 25329 13484
rect 25363 13481 25375 13515
rect 25317 13475 25375 13481
rect 25590 13472 25596 13524
rect 25648 13472 25654 13524
rect 26513 13515 26571 13521
rect 26513 13481 26525 13515
rect 26559 13512 26571 13515
rect 26602 13512 26608 13524
rect 26559 13484 26608 13512
rect 26559 13481 26571 13484
rect 26513 13475 26571 13481
rect 24673 13447 24731 13453
rect 24673 13413 24685 13447
rect 24719 13444 24731 13447
rect 26528 13444 26556 13475
rect 26602 13472 26608 13484
rect 26660 13472 26666 13524
rect 28445 13515 28503 13521
rect 28445 13512 28457 13515
rect 27724 13484 28457 13512
rect 27724 13444 27752 13484
rect 28445 13481 28457 13484
rect 28491 13481 28503 13515
rect 28445 13475 28503 13481
rect 28810 13472 28816 13524
rect 28868 13472 28874 13524
rect 28994 13472 29000 13524
rect 29052 13472 29058 13524
rect 29454 13472 29460 13524
rect 29512 13472 29518 13524
rect 30190 13472 30196 13524
rect 30248 13512 30254 13524
rect 30285 13515 30343 13521
rect 30285 13512 30297 13515
rect 30248 13484 30297 13512
rect 30248 13472 30254 13484
rect 30285 13481 30297 13484
rect 30331 13481 30343 13515
rect 30285 13475 30343 13481
rect 24719 13416 25452 13444
rect 24719 13413 24731 13416
rect 24673 13407 24731 13413
rect 23037 13379 23095 13385
rect 23037 13345 23049 13379
rect 23083 13376 23095 13379
rect 24489 13379 24547 13385
rect 23083 13348 23704 13376
rect 23083 13345 23095 13348
rect 23037 13339 23095 13345
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 20404 13212 22324 13240
rect 20404 13200 20410 13212
rect 12986 13172 12992 13184
rect 11348 13144 12992 13172
rect 9401 13135 9459 13141
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 19889 13175 19947 13181
rect 19889 13141 19901 13175
rect 19935 13172 19947 13175
rect 20162 13172 20168 13184
rect 19935 13144 20168 13172
rect 19935 13141 19947 13144
rect 19889 13135 19947 13141
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 21358 13132 21364 13184
rect 21416 13132 21422 13184
rect 23014 13132 23020 13184
rect 23072 13172 23078 13184
rect 23308 13172 23336 13268
rect 23676 13184 23704 13348
rect 24489 13345 24501 13379
rect 24535 13376 24547 13379
rect 24535 13348 24716 13376
rect 24535 13345 24547 13348
rect 24489 13339 24547 13345
rect 24305 13311 24363 13317
rect 24305 13277 24317 13311
rect 24351 13308 24363 13311
rect 24394 13308 24400 13320
rect 24351 13280 24400 13308
rect 24351 13277 24363 13280
rect 24305 13271 24363 13277
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24688 13184 24716 13348
rect 24946 13336 24952 13388
rect 25004 13336 25010 13388
rect 25038 13336 25044 13388
rect 25096 13376 25102 13388
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 25096 13348 25237 13376
rect 25096 13336 25102 13348
rect 25225 13345 25237 13348
rect 25271 13345 25283 13379
rect 25225 13339 25283 13345
rect 25314 13336 25320 13388
rect 25372 13376 25378 13388
rect 25424 13385 25452 13416
rect 25552 13416 26556 13444
rect 27554 13416 27752 13444
rect 25409 13379 25467 13385
rect 25409 13376 25421 13379
rect 25372 13348 25421 13376
rect 25372 13336 25378 13348
rect 25409 13345 25421 13348
rect 25455 13345 25467 13379
rect 25409 13339 25467 13345
rect 23072 13144 23336 13172
rect 23072 13132 23078 13144
rect 23658 13132 23664 13184
rect 23716 13132 23722 13184
rect 24670 13132 24676 13184
rect 24728 13172 24734 13184
rect 24765 13175 24823 13181
rect 24765 13172 24777 13175
rect 24728 13144 24777 13172
rect 24728 13132 24734 13144
rect 24765 13141 24777 13144
rect 24811 13141 24823 13175
rect 24964 13172 24992 13336
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13308 25191 13311
rect 25552 13308 25580 13416
rect 27982 13404 27988 13456
rect 28040 13404 28046 13456
rect 28074 13404 28080 13456
rect 28132 13444 28138 13456
rect 29012 13444 29040 13472
rect 28132 13416 28304 13444
rect 29012 13416 29408 13444
rect 28132 13404 28138 13416
rect 28276 13385 28304 13416
rect 25685 13379 25743 13385
rect 25685 13345 25697 13379
rect 25731 13376 25743 13379
rect 28261 13379 28319 13385
rect 25731 13348 26004 13376
rect 25731 13345 25743 13348
rect 25685 13339 25743 13345
rect 25179 13280 25580 13308
rect 25179 13277 25191 13280
rect 25133 13271 25191 13277
rect 25976 13252 26004 13348
rect 28261 13345 28273 13379
rect 28307 13345 28319 13379
rect 28261 13339 28319 13345
rect 28534 13336 28540 13388
rect 28592 13336 28598 13388
rect 28718 13336 28724 13388
rect 28776 13336 28782 13388
rect 28994 13336 29000 13388
rect 29052 13336 29058 13388
rect 29104 13385 29132 13416
rect 29089 13379 29147 13385
rect 29089 13345 29101 13379
rect 29135 13345 29147 13379
rect 29089 13339 29147 13345
rect 29178 13336 29184 13388
rect 29236 13376 29242 13388
rect 29380 13385 29408 13416
rect 29273 13379 29331 13385
rect 29273 13376 29285 13379
rect 29236 13348 29285 13376
rect 29236 13336 29242 13348
rect 29273 13345 29285 13348
rect 29319 13345 29331 13379
rect 29273 13339 29331 13345
rect 29365 13379 29423 13385
rect 29365 13345 29377 13379
rect 29411 13345 29423 13379
rect 29365 13339 29423 13345
rect 29549 13379 29607 13385
rect 29549 13345 29561 13379
rect 29595 13345 29607 13379
rect 29549 13339 29607 13345
rect 26050 13268 26056 13320
rect 26108 13268 26114 13320
rect 25958 13200 25964 13252
rect 26016 13200 26022 13252
rect 26068 13172 26096 13268
rect 28736 13240 28764 13336
rect 29564 13308 29592 13339
rect 30098 13336 30104 13388
rect 30156 13376 30162 13388
rect 30193 13379 30251 13385
rect 30193 13376 30205 13379
rect 30156 13348 30205 13376
rect 30156 13336 30162 13348
rect 30193 13345 30205 13348
rect 30239 13345 30251 13379
rect 30193 13339 30251 13345
rect 29012 13280 29592 13308
rect 29012 13249 29040 13280
rect 28276 13212 28764 13240
rect 28997 13243 29055 13249
rect 28276 13184 28304 13212
rect 28997 13209 29009 13243
rect 29043 13209 29055 13243
rect 28997 13203 29055 13209
rect 24964 13144 26096 13172
rect 24765 13135 24823 13141
rect 28258 13132 28264 13184
rect 28316 13132 28322 13184
rect 28718 13132 28724 13184
rect 28776 13172 28782 13184
rect 29089 13175 29147 13181
rect 29089 13172 29101 13175
rect 28776 13144 29101 13172
rect 28776 13132 28782 13144
rect 29089 13141 29101 13144
rect 29135 13141 29147 13175
rect 29089 13135 29147 13141
rect 552 13082 31648 13104
rect 552 13030 4285 13082
rect 4337 13030 4349 13082
rect 4401 13030 4413 13082
rect 4465 13030 4477 13082
rect 4529 13030 4541 13082
rect 4593 13030 12059 13082
rect 12111 13030 12123 13082
rect 12175 13030 12187 13082
rect 12239 13030 12251 13082
rect 12303 13030 12315 13082
rect 12367 13030 19833 13082
rect 19885 13030 19897 13082
rect 19949 13030 19961 13082
rect 20013 13030 20025 13082
rect 20077 13030 20089 13082
rect 20141 13030 27607 13082
rect 27659 13030 27671 13082
rect 27723 13030 27735 13082
rect 27787 13030 27799 13082
rect 27851 13030 27863 13082
rect 27915 13030 31648 13082
rect 552 13008 31648 13030
rect 1394 12928 1400 12980
rect 1452 12928 1458 12980
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12937 2927 12971
rect 2869 12931 2927 12937
rect 3973 12971 4031 12977
rect 3973 12937 3985 12971
rect 4019 12968 4031 12971
rect 4154 12968 4160 12980
rect 4019 12940 4160 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 1029 12903 1087 12909
rect 1029 12869 1041 12903
rect 1075 12900 1087 12903
rect 1412 12900 1440 12928
rect 2685 12903 2743 12909
rect 2685 12900 2697 12903
rect 1075 12872 1440 12900
rect 1504 12872 2697 12900
rect 1075 12869 1087 12872
rect 1029 12863 1087 12869
rect 1504 12841 1532 12872
rect 2685 12869 2697 12872
rect 2731 12869 2743 12903
rect 2884 12900 2912 12931
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 4706 12968 4712 12980
rect 4479 12940 4712 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5258 12928 5264 12980
rect 5316 12928 5322 12980
rect 5626 12928 5632 12980
rect 5684 12928 5690 12980
rect 5810 12928 5816 12980
rect 5868 12928 5874 12980
rect 8205 12971 8263 12977
rect 8205 12937 8217 12971
rect 8251 12968 8263 12971
rect 12894 12968 12900 12980
rect 8251 12940 12900 12968
rect 8251 12937 8263 12940
rect 8205 12931 8263 12937
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 13357 12971 13415 12977
rect 13357 12937 13369 12971
rect 13403 12968 13415 12971
rect 13906 12968 13912 12980
rect 13403 12940 13912 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 19426 12928 19432 12980
rect 19484 12928 19490 12980
rect 20162 12928 20168 12980
rect 20220 12928 20226 12980
rect 21821 12971 21879 12977
rect 21821 12937 21833 12971
rect 21867 12968 21879 12971
rect 22094 12968 22100 12980
rect 21867 12940 22100 12968
rect 21867 12937 21879 12940
rect 21821 12931 21879 12937
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 22373 12971 22431 12977
rect 22373 12937 22385 12971
rect 22419 12968 22431 12971
rect 22922 12968 22928 12980
rect 22419 12940 22928 12968
rect 22419 12937 22431 12940
rect 22373 12931 22431 12937
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 24394 12928 24400 12980
rect 24452 12968 24458 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 24452 12940 24777 12968
rect 24452 12928 24458 12940
rect 24765 12937 24777 12940
rect 24811 12968 24823 12971
rect 24854 12968 24860 12980
rect 24811 12940 24860 12968
rect 24811 12937 24823 12940
rect 24765 12931 24823 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 26418 12968 26424 12980
rect 25056 12940 26424 12968
rect 2884 12872 3648 12900
rect 2685 12863 2743 12869
rect 1489 12835 1547 12841
rect 1489 12801 1501 12835
rect 1535 12801 1547 12835
rect 1489 12795 1547 12801
rect 3620 12776 3648 12872
rect 5644 12832 5672 12928
rect 3712 12804 5672 12832
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2866 12764 2872 12776
rect 1443 12736 2872 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2866 12724 2872 12736
rect 2924 12764 2930 12776
rect 2924 12736 3556 12764
rect 2924 12724 2930 12736
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 3418 12696 3424 12708
rect 3108 12668 3424 12696
rect 3108 12656 3114 12668
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 3528 12696 3556 12736
rect 3602 12724 3608 12776
rect 3660 12724 3666 12776
rect 3712 12773 3740 12804
rect 3697 12767 3755 12773
rect 3697 12733 3709 12767
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4798 12764 4804 12776
rect 4387 12736 4804 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 3712 12696 3740 12727
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 5166 12764 5172 12776
rect 4908 12736 5172 12764
rect 4908 12696 4936 12736
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12764 5411 12767
rect 5828 12764 5856 12928
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 11974 12900 11980 12912
rect 11931 12872 11980 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 17678 12860 17684 12912
rect 17736 12860 17742 12912
rect 18325 12903 18383 12909
rect 18325 12900 18337 12903
rect 17788 12872 18337 12900
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6512 12804 6837 12832
rect 6512 12792 6518 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 8352 12804 8861 12832
rect 8352 12792 8358 12804
rect 8849 12801 8861 12804
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 17788 12832 17816 12872
rect 18325 12869 18337 12872
rect 18371 12869 18383 12903
rect 18325 12863 18383 12869
rect 16163 12804 17816 12832
rect 18233 12835 18291 12841
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 18279 12804 18552 12832
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 5997 12767 6055 12773
rect 5997 12764 6009 12767
rect 5399 12736 6009 12764
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 5997 12733 6009 12736
rect 6043 12733 6055 12767
rect 5997 12727 6055 12733
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12764 10563 12767
rect 11330 12764 11336 12776
rect 10551 12736 11336 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 10980 12708 11008 12736
rect 11330 12724 11336 12736
rect 11388 12764 11394 12776
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 11388 12736 11989 12764
rect 11388 12724 11394 12736
rect 11977 12733 11989 12736
rect 12023 12764 12035 12767
rect 12710 12764 12716 12776
rect 12023 12736 12716 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 15838 12724 15844 12776
rect 15896 12724 15902 12776
rect 18322 12724 18328 12776
rect 18380 12724 18386 12776
rect 18524 12773 18552 12804
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 19444 12764 19472 12928
rect 20180 12832 20208 12928
rect 23201 12903 23259 12909
rect 23201 12900 23213 12903
rect 22296 12872 23213 12900
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 20180 12804 20361 12832
rect 20349 12801 20361 12804
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 18555 12736 19472 12764
rect 20073 12767 20131 12773
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 20073 12733 20085 12767
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 3528 12668 3740 12696
rect 3804 12668 4936 12696
rect 2866 12637 2872 12640
rect 2853 12631 2872 12637
rect 2853 12597 2865 12631
rect 2924 12628 2930 12640
rect 3804 12637 3832 12668
rect 5718 12656 5724 12708
rect 5776 12696 5782 12708
rect 5813 12699 5871 12705
rect 5813 12696 5825 12699
rect 5776 12668 5825 12696
rect 5776 12656 5782 12668
rect 5813 12665 5825 12668
rect 5859 12665 5871 12699
rect 5813 12659 5871 12665
rect 6362 12656 6368 12708
rect 6420 12656 6426 12708
rect 7092 12699 7150 12705
rect 7092 12665 7104 12699
rect 7138 12696 7150 12699
rect 7190 12696 7196 12708
rect 7138 12668 7196 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7190 12656 7196 12668
rect 7248 12656 7254 12708
rect 7282 12656 7288 12708
rect 7340 12696 7346 12708
rect 9094 12699 9152 12705
rect 9094 12696 9106 12699
rect 7340 12668 9106 12696
rect 7340 12656 7346 12668
rect 9094 12665 9106 12668
rect 9140 12665 9152 12699
rect 9094 12659 9152 12665
rect 9398 12656 9404 12708
rect 9456 12696 9462 12708
rect 10750 12699 10808 12705
rect 10750 12696 10762 12699
rect 9456 12668 10762 12696
rect 9456 12656 9462 12668
rect 10750 12665 10762 12668
rect 10796 12665 10808 12699
rect 10750 12659 10808 12665
rect 10962 12656 10968 12708
rect 11020 12656 11026 12708
rect 12244 12699 12302 12705
rect 12244 12665 12256 12699
rect 12290 12696 12302 12699
rect 13170 12696 13176 12708
rect 12290 12668 13176 12696
rect 12290 12665 12302 12668
rect 12244 12659 12302 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 16850 12656 16856 12708
rect 16908 12656 16914 12708
rect 17604 12668 18000 12696
rect 3789 12631 3847 12637
rect 3789 12628 3801 12631
rect 2924 12600 3801 12628
rect 2853 12591 2872 12597
rect 2866 12588 2872 12591
rect 2924 12588 2930 12600
rect 3789 12597 3801 12600
rect 3835 12597 3847 12631
rect 3789 12591 3847 12597
rect 6086 12588 6092 12640
rect 6144 12588 6150 12640
rect 6181 12631 6239 12637
rect 6181 12597 6193 12631
rect 6227 12628 6239 12631
rect 6730 12628 6736 12640
rect 6227 12600 6736 12628
rect 6227 12597 6239 12600
rect 6181 12591 6239 12597
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 11606 12628 11612 12640
rect 10275 12600 11612 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 17604 12637 17632 12668
rect 17972 12640 18000 12668
rect 18966 12656 18972 12708
rect 19024 12696 19030 12708
rect 20088 12696 20116 12727
rect 21358 12724 21364 12776
rect 21416 12764 21422 12776
rect 21416 12736 21482 12764
rect 21416 12724 21422 12736
rect 20346 12696 20352 12708
rect 19024 12668 20352 12696
rect 19024 12656 19030 12668
rect 20346 12656 20352 12668
rect 20404 12656 20410 12708
rect 22189 12699 22247 12705
rect 22189 12665 22201 12699
rect 22235 12696 22247 12699
rect 22296 12696 22324 12872
rect 23201 12869 23213 12872
rect 23247 12900 23259 12903
rect 24412 12900 24440 12928
rect 23247 12872 24440 12900
rect 23247 12869 23259 12872
rect 23201 12863 23259 12869
rect 22235 12668 22324 12696
rect 22388 12804 22968 12832
rect 22388 12705 22416 12804
rect 22940 12773 22968 12804
rect 22649 12767 22707 12773
rect 22649 12764 22661 12767
rect 22480 12736 22661 12764
rect 22388 12699 22447 12705
rect 22388 12668 22401 12699
rect 22235 12665 22247 12668
rect 22189 12659 22247 12665
rect 22389 12665 22401 12668
rect 22435 12665 22447 12699
rect 22389 12659 22447 12665
rect 17589 12631 17647 12637
rect 17589 12597 17601 12631
rect 17635 12597 17647 12631
rect 17589 12591 17647 12597
rect 17862 12588 17868 12640
rect 17920 12588 17926 12640
rect 17954 12588 17960 12640
rect 18012 12588 18018 12640
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12628 18107 12631
rect 18414 12628 18420 12640
rect 18095 12600 18420 12628
rect 18095 12597 18107 12600
rect 18049 12591 18107 12597
rect 18414 12588 18420 12600
rect 18472 12628 18478 12640
rect 22480 12628 22508 12736
rect 22649 12733 22661 12736
rect 22695 12733 22707 12767
rect 22649 12727 22707 12733
rect 22925 12767 22983 12773
rect 22925 12733 22937 12767
rect 22971 12764 22983 12767
rect 23293 12767 23351 12773
rect 23293 12764 23305 12767
rect 22971 12736 23305 12764
rect 22971 12733 22983 12736
rect 22925 12727 22983 12733
rect 23293 12733 23305 12736
rect 23339 12733 23351 12767
rect 23293 12727 23351 12733
rect 23474 12724 23480 12776
rect 23532 12724 23538 12776
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 25056 12773 25084 12940
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 29178 12928 29184 12980
rect 29236 12968 29242 12980
rect 30837 12971 30895 12977
rect 30837 12968 30849 12971
rect 29236 12940 30849 12968
rect 29236 12928 29242 12940
rect 30837 12937 30849 12940
rect 30883 12937 30895 12971
rect 30837 12931 30895 12937
rect 25501 12903 25559 12909
rect 25501 12869 25513 12903
rect 25547 12900 25559 12903
rect 27154 12900 27160 12912
rect 25547 12872 27160 12900
rect 25547 12869 25559 12872
rect 25501 12863 25559 12869
rect 27154 12860 27160 12872
rect 27212 12860 27218 12912
rect 28092 12872 28948 12900
rect 28092 12844 28120 12872
rect 25133 12835 25191 12841
rect 25133 12801 25145 12835
rect 25179 12832 25191 12835
rect 25179 12804 25544 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 25041 12767 25099 12773
rect 25041 12764 25053 12767
rect 23716 12736 25053 12764
rect 23716 12724 23722 12736
rect 24596 12705 24624 12736
rect 25041 12733 25053 12736
rect 25087 12733 25099 12767
rect 25041 12727 25099 12733
rect 25222 12724 25228 12776
rect 25280 12724 25286 12776
rect 25516 12773 25544 12804
rect 25958 12792 25964 12844
rect 26016 12832 26022 12844
rect 26016 12804 26924 12832
rect 26016 12792 26022 12804
rect 25317 12767 25375 12773
rect 25317 12733 25329 12767
rect 25363 12733 25375 12767
rect 25317 12727 25375 12733
rect 25501 12767 25559 12773
rect 25501 12733 25513 12767
rect 25547 12733 25559 12767
rect 25501 12727 25559 12733
rect 26145 12767 26203 12773
rect 26145 12733 26157 12767
rect 26191 12764 26203 12767
rect 26234 12764 26240 12776
rect 26191 12736 26240 12764
rect 26191 12733 26203 12736
rect 26145 12727 26203 12733
rect 23017 12699 23075 12705
rect 23017 12665 23029 12699
rect 23063 12665 23075 12699
rect 23017 12659 23075 12665
rect 24581 12699 24639 12705
rect 24581 12665 24593 12699
rect 24627 12665 24639 12699
rect 25332 12696 25360 12727
rect 26234 12724 26240 12736
rect 26292 12724 26298 12776
rect 26896 12773 26924 12804
rect 28074 12792 28080 12844
rect 28132 12792 28138 12844
rect 28718 12792 28724 12844
rect 28776 12832 28782 12844
rect 28776 12804 28856 12832
rect 28776 12792 28782 12804
rect 26881 12767 26939 12773
rect 26881 12733 26893 12767
rect 26927 12764 26939 12767
rect 28534 12764 28540 12776
rect 26927 12736 28540 12764
rect 26927 12733 26939 12736
rect 26881 12727 26939 12733
rect 28534 12724 28540 12736
rect 28592 12724 28598 12776
rect 28626 12724 28632 12776
rect 28684 12724 28690 12776
rect 28828 12773 28856 12804
rect 28813 12767 28871 12773
rect 28813 12733 28825 12767
rect 28859 12733 28871 12767
rect 28920 12764 28948 12872
rect 30098 12792 30104 12844
rect 30156 12832 30162 12844
rect 30156 12804 30972 12832
rect 30156 12792 30162 12804
rect 30944 12773 30972 12804
rect 29089 12767 29147 12773
rect 29089 12764 29101 12767
rect 28920 12736 29101 12764
rect 28813 12727 28871 12733
rect 29089 12733 29101 12736
rect 29135 12733 29147 12767
rect 29089 12727 29147 12733
rect 30929 12767 30987 12773
rect 30929 12733 30941 12767
rect 30975 12733 30987 12767
rect 30929 12727 30987 12733
rect 24581 12659 24639 12665
rect 24964 12668 25360 12696
rect 28721 12699 28779 12705
rect 18472 12600 22508 12628
rect 18472 12588 18478 12600
rect 22554 12588 22560 12640
rect 22612 12588 22618 12640
rect 22738 12588 22744 12640
rect 22796 12628 22802 12640
rect 22833 12631 22891 12637
rect 22833 12628 22845 12631
rect 22796 12600 22845 12628
rect 22796 12588 22802 12600
rect 22833 12597 22845 12600
rect 22879 12597 22891 12631
rect 22833 12591 22891 12597
rect 22922 12588 22928 12640
rect 22980 12628 22986 12640
rect 23032 12628 23060 12659
rect 24964 12640 24992 12668
rect 28721 12665 28733 12699
rect 28767 12696 28779 12699
rect 29365 12699 29423 12705
rect 29365 12696 29377 12699
rect 28767 12668 29377 12696
rect 28767 12665 28779 12668
rect 28721 12659 28779 12665
rect 29365 12665 29377 12668
rect 29411 12665 29423 12699
rect 31021 12699 31079 12705
rect 31021 12696 31033 12699
rect 30590 12668 31033 12696
rect 29365 12659 29423 12665
rect 31021 12665 31033 12668
rect 31067 12665 31079 12699
rect 31021 12659 31079 12665
rect 24670 12628 24676 12640
rect 22980 12600 24676 12628
rect 22980 12588 22986 12600
rect 24670 12588 24676 12600
rect 24728 12628 24734 12640
rect 24781 12631 24839 12637
rect 24781 12628 24793 12631
rect 24728 12600 24793 12628
rect 24728 12588 24734 12600
rect 24781 12597 24793 12600
rect 24827 12597 24839 12631
rect 24781 12591 24839 12597
rect 24946 12588 24952 12640
rect 25004 12588 25010 12640
rect 25130 12588 25136 12640
rect 25188 12628 25194 12640
rect 25961 12631 26019 12637
rect 25961 12628 25973 12631
rect 25188 12600 25973 12628
rect 25188 12588 25194 12600
rect 25961 12597 25973 12600
rect 26007 12628 26019 12631
rect 26786 12628 26792 12640
rect 26007 12600 26792 12628
rect 26007 12597 26019 12600
rect 25961 12591 26019 12597
rect 26786 12588 26792 12600
rect 26844 12588 26850 12640
rect 26970 12588 26976 12640
rect 27028 12588 27034 12640
rect 552 12538 31808 12560
rect 552 12486 8172 12538
rect 8224 12486 8236 12538
rect 8288 12486 8300 12538
rect 8352 12486 8364 12538
rect 8416 12486 8428 12538
rect 8480 12486 15946 12538
rect 15998 12486 16010 12538
rect 16062 12486 16074 12538
rect 16126 12486 16138 12538
rect 16190 12486 16202 12538
rect 16254 12486 23720 12538
rect 23772 12486 23784 12538
rect 23836 12486 23848 12538
rect 23900 12486 23912 12538
rect 23964 12486 23976 12538
rect 24028 12486 31494 12538
rect 31546 12486 31558 12538
rect 31610 12486 31622 12538
rect 31674 12486 31686 12538
rect 31738 12486 31750 12538
rect 31802 12486 31808 12538
rect 552 12464 31808 12486
rect 3050 12424 3056 12436
rect 2516 12396 3056 12424
rect 2516 12297 2544 12396
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3191 12396 3740 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3602 12356 3608 12368
rect 2792 12328 3608 12356
rect 2792 12297 2820 12328
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 3712 12365 3740 12396
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 5169 12427 5227 12433
rect 5169 12424 5181 12427
rect 4120 12396 5181 12424
rect 4120 12384 4126 12396
rect 5169 12393 5181 12396
rect 5215 12424 5227 12427
rect 5350 12424 5356 12436
rect 5215 12396 5356 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 5629 12427 5687 12433
rect 5629 12393 5641 12427
rect 5675 12424 5687 12427
rect 5675 12396 6040 12424
rect 5675 12393 5687 12396
rect 5629 12387 5687 12393
rect 3697 12359 3755 12365
rect 3697 12325 3709 12359
rect 3743 12325 3755 12359
rect 3697 12319 3755 12325
rect 4706 12316 4712 12368
rect 4764 12316 4770 12368
rect 5261 12359 5319 12365
rect 5261 12325 5273 12359
rect 5307 12325 5319 12359
rect 5261 12319 5319 12325
rect 5466 12359 5524 12365
rect 5466 12325 5478 12359
rect 5512 12356 5524 12359
rect 6012 12356 6040 12396
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6144 12396 6929 12424
rect 6144 12384 6150 12396
rect 6181 12359 6239 12365
rect 6181 12356 6193 12359
rect 5512 12328 5580 12356
rect 6012 12328 6193 12356
rect 5512 12325 5524 12328
rect 5466 12319 5524 12325
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12257 2375 12291
rect 2317 12251 2375 12257
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12257 2559 12291
rect 2501 12251 2559 12257
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 2332 12152 2360 12251
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 2455 12192 2697 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2685 12189 2697 12192
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 3384 12192 3433 12220
rect 3384 12180 3390 12192
rect 3421 12189 3433 12192
rect 3467 12189 3479 12223
rect 5276 12220 5304 12319
rect 5552 12288 5580 12328
rect 6181 12325 6193 12328
rect 6227 12325 6239 12359
rect 6181 12319 6239 12325
rect 6288 12288 6316 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 13078 12424 13084 12436
rect 12391 12396 13084 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 14461 12427 14519 12433
rect 14461 12393 14473 12427
rect 14507 12424 14519 12427
rect 14734 12424 14740 12436
rect 14507 12396 14740 12424
rect 14507 12393 14519 12396
rect 14461 12387 14519 12393
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15933 12427 15991 12433
rect 15933 12393 15945 12427
rect 15979 12424 15991 12427
rect 16390 12424 16396 12436
rect 15979 12396 16396 12424
rect 15979 12393 15991 12396
rect 15933 12387 15991 12393
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 16945 12427 17003 12433
rect 16945 12424 16957 12427
rect 16908 12396 16957 12424
rect 16908 12384 16914 12396
rect 16945 12393 16957 12396
rect 16991 12393 17003 12427
rect 16945 12387 17003 12393
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17828 12396 17877 12424
rect 17828 12384 17834 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 18049 12427 18107 12433
rect 18049 12393 18061 12427
rect 18095 12424 18107 12427
rect 18322 12424 18328 12436
rect 18095 12396 18328 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20530 12424 20536 12436
rect 20119 12396 20536 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 22646 12384 22652 12436
rect 22704 12384 22710 12436
rect 26418 12384 26424 12436
rect 26476 12384 26482 12436
rect 28810 12424 28816 12436
rect 28460 12396 28816 12424
rect 9232 12328 10456 12356
rect 5552 12260 6316 12288
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12288 7159 12291
rect 7190 12288 7196 12300
rect 7147 12260 7196 12288
rect 7147 12257 7159 12260
rect 7101 12251 7159 12257
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 7282 12248 7288 12300
rect 7340 12248 7346 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 9232 12297 9260 12328
rect 10428 12300 10456 12328
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 18233 12359 18291 12365
rect 18233 12356 18245 12359
rect 12768 12328 14596 12356
rect 12768 12316 12774 12328
rect 9033 12291 9091 12297
rect 9033 12288 9045 12291
rect 8076 12260 9045 12288
rect 8076 12248 8082 12260
rect 9033 12257 9045 12260
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12257 9275 12291
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9217 12251 9275 12257
rect 9324 12260 9597 12288
rect 6362 12220 6368 12232
rect 5276 12192 6368 12220
rect 3421 12183 3479 12189
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 9324 12220 9352 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 10410 12248 10416 12300
rect 10468 12288 10474 12300
rect 13096 12297 13124 12328
rect 11221 12291 11279 12297
rect 11221 12288 11233 12291
rect 10468 12260 11233 12288
rect 10468 12248 10474 12260
rect 11221 12257 11233 12260
rect 11267 12257 11279 12291
rect 11221 12251 11279 12257
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12257 13139 12291
rect 13081 12251 13139 12257
rect 13348 12291 13406 12297
rect 13348 12257 13360 12291
rect 13394 12288 13406 12291
rect 13722 12288 13728 12300
rect 13394 12260 13728 12288
rect 13394 12257 13406 12260
rect 13348 12251 13406 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14568 12297 14596 12328
rect 17880 12328 18245 12356
rect 17880 12300 17908 12328
rect 18233 12325 18245 12328
rect 18279 12356 18291 12359
rect 18938 12359 18996 12365
rect 18938 12356 18950 12359
rect 18279 12328 18950 12356
rect 18279 12325 18291 12328
rect 18233 12319 18291 12325
rect 18938 12325 18950 12328
rect 18984 12325 18996 12359
rect 18938 12319 18996 12325
rect 21284 12328 22048 12356
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12288 14611 12291
rect 14642 12288 14648 12300
rect 14599 12260 14648 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 14820 12291 14878 12297
rect 14820 12257 14832 12291
rect 14866 12288 14878 12291
rect 15194 12288 15200 12300
rect 14866 12260 15200 12288
rect 14866 12257 14878 12260
rect 14820 12251 14878 12257
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 17037 12291 17095 12297
rect 17037 12257 17049 12291
rect 17083 12257 17095 12291
rect 17037 12251 17095 12257
rect 6604 12192 9352 12220
rect 6604 12180 6610 12192
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 10962 12180 10968 12232
rect 11020 12180 11026 12232
rect 17052 12220 17080 12251
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 17405 12291 17463 12297
rect 17405 12288 17417 12291
rect 17276 12260 17417 12288
rect 17276 12248 17282 12260
rect 17405 12257 17417 12260
rect 17451 12257 17463 12291
rect 17405 12251 17463 12257
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 17862 12288 17868 12300
rect 17727 12260 17868 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 17052 12192 17356 12220
rect 2774 12152 2780 12164
rect 2332 12124 2780 12152
rect 2774 12112 2780 12124
rect 2832 12112 2838 12164
rect 9416 12152 9444 12180
rect 17328 12164 17356 12192
rect 5460 12124 6776 12152
rect 5460 12093 5488 12124
rect 6748 12096 6776 12124
rect 8956 12124 9444 12152
rect 8956 12096 8984 12124
rect 17310 12112 17316 12164
rect 17368 12112 17374 12164
rect 17420 12152 17448 12251
rect 17512 12220 17540 12251
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 17954 12248 17960 12300
rect 18012 12248 18018 12300
rect 18322 12248 18328 12300
rect 18380 12248 18386 12300
rect 21284 12297 21312 12328
rect 22020 12300 22048 12328
rect 22554 12316 22560 12368
rect 22612 12356 22618 12368
rect 23293 12359 23351 12365
rect 23293 12356 23305 12359
rect 22612 12328 23305 12356
rect 22612 12316 22618 12328
rect 23293 12325 23305 12328
rect 23339 12325 23351 12359
rect 23293 12319 23351 12325
rect 25590 12316 25596 12368
rect 25648 12316 25654 12368
rect 26878 12316 26884 12368
rect 26936 12316 26942 12368
rect 21542 12297 21548 12300
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12257 21327 12291
rect 21269 12251 21327 12257
rect 21536 12251 21548 12297
rect 21542 12248 21548 12251
rect 21600 12248 21606 12300
rect 22002 12248 22008 12300
rect 22060 12248 22066 12300
rect 24302 12248 24308 12300
rect 24360 12248 24366 12300
rect 28460 12297 28488 12396
rect 28810 12384 28816 12396
rect 28868 12424 28874 12436
rect 30745 12427 30803 12433
rect 30745 12424 30757 12427
rect 28868 12396 30757 12424
rect 28868 12384 28874 12396
rect 30745 12393 30757 12396
rect 30791 12393 30803 12427
rect 30745 12387 30803 12393
rect 30006 12316 30012 12368
rect 30064 12316 30070 12368
rect 28445 12291 28503 12297
rect 28445 12257 28457 12291
rect 28491 12257 28503 12291
rect 28445 12251 28503 12257
rect 17586 12220 17592 12232
rect 17512 12192 17592 12220
rect 17586 12180 17592 12192
rect 17644 12220 17650 12232
rect 18046 12220 18052 12232
rect 17644 12192 18052 12220
rect 17644 12180 17650 12192
rect 18046 12180 18052 12192
rect 18104 12220 18110 12232
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 18104 12192 18153 12220
rect 18104 12180 18110 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 18340 12152 18368 12248
rect 18690 12180 18696 12232
rect 18748 12180 18754 12232
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 27154 12180 27160 12232
rect 27212 12220 27218 12232
rect 27893 12223 27951 12229
rect 27893 12220 27905 12223
rect 27212 12192 27905 12220
rect 27212 12180 27218 12192
rect 27893 12189 27905 12192
rect 27939 12189 27951 12223
rect 27893 12183 27951 12189
rect 28169 12223 28227 12229
rect 28169 12189 28181 12223
rect 28215 12189 28227 12223
rect 28169 12183 28227 12189
rect 17420 12124 18368 12152
rect 26786 12112 26792 12164
rect 26844 12112 26850 12164
rect 28184 12152 28212 12183
rect 28258 12180 28264 12232
rect 28316 12220 28322 12232
rect 28353 12223 28411 12229
rect 28353 12220 28365 12223
rect 28316 12192 28365 12220
rect 28316 12180 28322 12192
rect 28353 12189 28365 12192
rect 28399 12189 28411 12223
rect 28997 12223 29055 12229
rect 28997 12220 29009 12223
rect 28353 12183 28411 12189
rect 28644 12192 29009 12220
rect 28644 12152 28672 12192
rect 28997 12189 29009 12192
rect 29043 12189 29055 12223
rect 29273 12223 29331 12229
rect 29273 12220 29285 12223
rect 28997 12183 29055 12189
rect 29104 12192 29285 12220
rect 28184 12124 28672 12152
rect 28813 12155 28871 12161
rect 5445 12087 5503 12093
rect 5445 12053 5457 12087
rect 5491 12053 5503 12087
rect 5445 12047 5503 12053
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6089 12087 6147 12093
rect 6089 12084 6101 12087
rect 6052 12056 6101 12084
rect 6052 12044 6058 12056
rect 6089 12053 6101 12056
rect 6135 12053 6147 12087
rect 6089 12047 6147 12053
rect 6730 12044 6736 12096
rect 6788 12044 6794 12096
rect 8938 12044 8944 12096
rect 8996 12044 9002 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 9456 12056 9689 12084
rect 9456 12044 9462 12056
rect 9677 12053 9689 12056
rect 9723 12084 9735 12087
rect 11146 12084 11152 12096
rect 9723 12056 11152 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 16850 12044 16856 12096
rect 16908 12084 16914 12096
rect 21634 12084 21640 12096
rect 16908 12056 21640 12084
rect 16908 12044 16914 12056
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 21910 12044 21916 12096
rect 21968 12084 21974 12096
rect 23385 12087 23443 12093
rect 23385 12084 23397 12087
rect 21968 12056 23397 12084
rect 21968 12044 21974 12056
rect 23385 12053 23397 12056
rect 23431 12084 23443 12087
rect 23474 12084 23480 12096
rect 23431 12056 23480 12084
rect 23431 12053 23443 12056
rect 23385 12047 23443 12053
rect 23474 12044 23480 12056
rect 23532 12044 23538 12096
rect 24670 12044 24676 12096
rect 24728 12084 24734 12096
rect 26053 12087 26111 12093
rect 26053 12084 26065 12087
rect 24728 12056 26065 12084
rect 24728 12044 24734 12056
rect 26053 12053 26065 12056
rect 26099 12053 26111 12087
rect 26804 12084 26832 12112
rect 28184 12084 28212 12124
rect 28813 12121 28825 12155
rect 28859 12152 28871 12155
rect 29104 12152 29132 12192
rect 29273 12189 29285 12192
rect 29319 12189 29331 12223
rect 29273 12183 29331 12189
rect 28859 12124 29132 12152
rect 28859 12121 28871 12124
rect 28813 12115 28871 12121
rect 26804 12056 28212 12084
rect 26053 12047 26111 12053
rect 552 11994 31648 12016
rect 552 11942 4285 11994
rect 4337 11942 4349 11994
rect 4401 11942 4413 11994
rect 4465 11942 4477 11994
rect 4529 11942 4541 11994
rect 4593 11942 12059 11994
rect 12111 11942 12123 11994
rect 12175 11942 12187 11994
rect 12239 11942 12251 11994
rect 12303 11942 12315 11994
rect 12367 11942 19833 11994
rect 19885 11942 19897 11994
rect 19949 11942 19961 11994
rect 20013 11942 20025 11994
rect 20077 11942 20089 11994
rect 20141 11942 27607 11994
rect 27659 11942 27671 11994
rect 27723 11942 27735 11994
rect 27787 11942 27799 11994
rect 27851 11942 27863 11994
rect 27915 11942 31648 11994
rect 552 11920 31648 11942
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 4706 11880 4712 11892
rect 4663 11852 4712 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 6362 11840 6368 11892
rect 6420 11880 6426 11892
rect 6733 11883 6791 11889
rect 6733 11880 6745 11883
rect 6420 11852 6745 11880
rect 6420 11840 6426 11852
rect 6733 11849 6745 11852
rect 6779 11880 6791 11883
rect 6779 11852 6914 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 6886 11812 6914 11852
rect 10410 11840 10416 11892
rect 10468 11840 10474 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 14829 11883 14887 11889
rect 14829 11880 14841 11883
rect 14700 11852 14841 11880
rect 14700 11840 14706 11852
rect 14829 11849 14841 11852
rect 14875 11849 14887 11883
rect 14829 11843 14887 11849
rect 15010 11840 15016 11892
rect 15068 11880 15074 11892
rect 15068 11852 16160 11880
rect 15068 11840 15074 11852
rect 8662 11812 8668 11824
rect 6886 11784 8668 11812
rect 7190 11744 7196 11756
rect 4632 11716 5120 11744
rect 4632 11688 4660 11716
rect 4614 11636 4620 11688
rect 4672 11636 4678 11688
rect 5092 11685 5120 11716
rect 6472 11716 7196 11744
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 5077 11679 5135 11685
rect 5077 11645 5089 11679
rect 5123 11645 5135 11679
rect 5077 11639 5135 11645
rect 4724 11608 4752 11639
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5994 11676 6000 11688
rect 5224 11648 6000 11676
rect 5224 11636 5230 11648
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6472 11685 6500 11716
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 8018 11744 8024 11756
rect 7392 11716 8024 11744
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11645 6331 11679
rect 6273 11639 6331 11645
rect 6457 11679 6515 11685
rect 6457 11645 6469 11679
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 5353 11611 5411 11617
rect 5353 11608 5365 11611
rect 4724 11580 5365 11608
rect 5353 11577 5365 11580
rect 5399 11608 5411 11611
rect 5718 11608 5724 11620
rect 5399 11580 5724 11608
rect 5399 11577 5411 11580
rect 5353 11571 5411 11577
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 6288 11608 6316 11639
rect 6917 11611 6975 11617
rect 6288 11580 6592 11608
rect 6564 11552 6592 11580
rect 6917 11577 6929 11611
rect 6963 11608 6975 11611
rect 7282 11608 7288 11620
rect 6963 11580 7288 11608
rect 6963 11577 6975 11580
rect 6917 11571 6975 11577
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 5810 11500 5816 11552
rect 5868 11500 5874 11552
rect 6546 11500 6552 11552
rect 6604 11500 6610 11552
rect 6730 11549 6736 11552
rect 6717 11543 6736 11549
rect 6717 11509 6729 11543
rect 6788 11540 6794 11552
rect 7392 11540 7420 11716
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8128 11753 8156 11784
rect 8662 11772 8668 11784
rect 8720 11772 8726 11824
rect 13630 11772 13636 11824
rect 13688 11812 13694 11824
rect 14093 11815 14151 11821
rect 14093 11812 14105 11815
rect 13688 11784 14105 11812
rect 13688 11772 13694 11784
rect 14093 11781 14105 11784
rect 14139 11812 14151 11815
rect 15194 11812 15200 11824
rect 14139 11784 15200 11812
rect 14139 11781 14151 11784
rect 14093 11775 14151 11781
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 9398 11744 9404 11756
rect 8113 11707 8171 11713
rect 8680 11716 9404 11744
rect 7466 11636 7472 11688
rect 7524 11636 7530 11688
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 7929 11679 7987 11685
rect 7699 11648 7788 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 7760 11617 7788 11648
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 8036 11676 8064 11704
rect 7975 11648 8064 11676
rect 8389 11679 8447 11685
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 8389 11645 8401 11679
rect 8435 11645 8447 11679
rect 8389 11639 8447 11645
rect 7745 11611 7803 11617
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 8404 11608 8432 11639
rect 8570 11636 8576 11688
rect 8628 11636 8634 11688
rect 8680 11685 8708 11716
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 15470 11744 15476 11756
rect 14936 11716 15476 11744
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11645 10747 11679
rect 10689 11639 10747 11645
rect 7791 11580 8432 11608
rect 8481 11611 8539 11617
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 8481 11577 8493 11611
rect 8527 11608 8539 11611
rect 8941 11611 8999 11617
rect 8941 11608 8953 11611
rect 8527 11580 8953 11608
rect 8527 11577 8539 11580
rect 8481 11571 8539 11577
rect 8941 11577 8953 11580
rect 8987 11577 8999 11611
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 10166 11580 10609 11608
rect 8941 11571 8999 11577
rect 10597 11577 10609 11580
rect 10643 11577 10655 11611
rect 10597 11571 10655 11577
rect 6788 11512 7420 11540
rect 6717 11503 6736 11509
rect 6730 11500 6736 11503
rect 6788 11500 6794 11512
rect 7558 11500 7564 11552
rect 7616 11500 7622 11552
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 10704 11540 10732 11639
rect 13354 11636 13360 11688
rect 13412 11676 13418 11688
rect 13814 11676 13820 11688
rect 13412 11648 13820 11676
rect 13412 11636 13418 11648
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 14936 11685 14964 11716
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15010 11636 15016 11688
rect 15068 11676 15074 11688
rect 16132 11685 16160 11852
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 18509 11883 18567 11889
rect 18509 11880 18521 11883
rect 17828 11852 18521 11880
rect 17828 11840 17834 11852
rect 18509 11849 18521 11852
rect 18555 11849 18567 11883
rect 18509 11843 18567 11849
rect 18690 11840 18696 11892
rect 18748 11840 18754 11892
rect 20533 11883 20591 11889
rect 20533 11849 20545 11883
rect 20579 11880 20591 11883
rect 20622 11880 20628 11892
rect 20579 11852 20628 11880
rect 20579 11849 20591 11852
rect 20533 11843 20591 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 21468 11852 22416 11880
rect 18708 11744 18736 11840
rect 19153 11747 19211 11753
rect 19153 11744 19165 11747
rect 18708 11716 19165 11744
rect 19153 11713 19165 11716
rect 19199 11713 19211 11747
rect 19153 11707 19211 11713
rect 15289 11679 15347 11685
rect 15289 11676 15301 11679
rect 15068 11648 15301 11676
rect 15068 11636 15074 11648
rect 15289 11645 15301 11648
rect 15335 11645 15347 11679
rect 15565 11679 15623 11685
rect 15565 11676 15577 11679
rect 15289 11639 15347 11645
rect 15488 11648 15577 11676
rect 11885 11611 11943 11617
rect 11885 11577 11897 11611
rect 11931 11608 11943 11611
rect 13541 11611 13599 11617
rect 13541 11608 13553 11611
rect 11931 11580 13553 11608
rect 11931 11577 11943 11580
rect 11885 11571 11943 11577
rect 13541 11577 13553 11580
rect 13587 11577 13599 11611
rect 13541 11571 13599 11577
rect 13722 11568 13728 11620
rect 13780 11568 13786 11620
rect 10560 11512 10732 11540
rect 10560 11500 10566 11512
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11112 11512 11805 11540
rect 11112 11500 11118 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 13446 11540 13452 11552
rect 13228 11512 13452 11540
rect 13228 11500 13234 11512
rect 13446 11500 13452 11512
rect 13504 11540 13510 11552
rect 15488 11549 15516 11648
rect 15565 11645 15577 11648
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11676 16175 11679
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 16163 11648 16221 11676
rect 16163 11645 16175 11648
rect 16117 11639 16175 11645
rect 16209 11645 16221 11648
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 16761 11679 16819 11685
rect 16761 11676 16773 11679
rect 16448 11648 16773 11676
rect 16448 11636 16454 11648
rect 16761 11645 16773 11648
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 19058 11676 19064 11688
rect 18923 11648 19064 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 15838 11568 15844 11620
rect 15896 11608 15902 11620
rect 16408 11608 16436 11636
rect 15896 11580 16436 11608
rect 15896 11568 15902 11580
rect 17034 11568 17040 11620
rect 17092 11568 17098 11620
rect 18785 11611 18843 11617
rect 18785 11608 18797 11611
rect 18262 11580 18797 11608
rect 18785 11577 18797 11580
rect 18831 11577 18843 11611
rect 18785 11571 18843 11577
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13504 11512 13921 11540
rect 13504 11500 13510 11512
rect 13909 11509 13921 11512
rect 13955 11509 13967 11543
rect 13909 11503 13967 11509
rect 15473 11543 15531 11549
rect 15473 11509 15485 11543
rect 15519 11509 15531 11543
rect 15473 11503 15531 11509
rect 15746 11500 15752 11552
rect 15804 11500 15810 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 18690 11540 18696 11552
rect 17368 11512 18696 11540
rect 17368 11500 17374 11512
rect 18690 11500 18696 11512
rect 18748 11540 18754 11552
rect 18892 11540 18920 11639
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 19168 11676 19196 11707
rect 21468 11685 21496 11852
rect 22388 11812 22416 11852
rect 22830 11840 22836 11892
rect 22888 11840 22894 11892
rect 23566 11840 23572 11892
rect 23624 11840 23630 11892
rect 24489 11883 24547 11889
rect 24489 11849 24501 11883
rect 24535 11880 24547 11883
rect 24578 11880 24584 11892
rect 24535 11852 24584 11880
rect 24535 11849 24547 11852
rect 24489 11843 24547 11849
rect 24578 11840 24584 11852
rect 24636 11840 24642 11892
rect 25501 11883 25559 11889
rect 25501 11849 25513 11883
rect 25547 11880 25559 11883
rect 25590 11880 25596 11892
rect 25547 11852 25596 11880
rect 25547 11849 25559 11852
rect 25501 11843 25559 11849
rect 25590 11840 25596 11852
rect 25648 11840 25654 11892
rect 28350 11880 28356 11892
rect 26206 11852 28356 11880
rect 23584 11812 23612 11840
rect 24670 11812 24676 11824
rect 22388 11784 22968 11812
rect 23584 11784 24676 11812
rect 22940 11756 22968 11784
rect 24670 11772 24676 11784
rect 24728 11812 24734 11824
rect 24728 11784 25176 11812
rect 24728 11772 24734 11784
rect 22922 11704 22928 11756
rect 22980 11704 22986 11756
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 23532 11716 24716 11744
rect 23532 11704 23538 11716
rect 24688 11688 24716 11716
rect 21453 11679 21511 11685
rect 21453 11676 21465 11679
rect 19168 11648 21465 11676
rect 21453 11645 21465 11648
rect 21499 11645 21511 11679
rect 21453 11639 21511 11645
rect 21542 11636 21548 11688
rect 21600 11636 21606 11688
rect 24670 11636 24676 11688
rect 24728 11636 24734 11688
rect 24946 11636 24952 11688
rect 25004 11636 25010 11688
rect 25148 11685 25176 11784
rect 25682 11772 25688 11824
rect 25740 11772 25746 11824
rect 25133 11679 25191 11685
rect 25133 11645 25145 11679
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 25593 11679 25651 11685
rect 25593 11645 25605 11679
rect 25639 11676 25651 11679
rect 25700 11676 25728 11772
rect 25639 11648 25728 11676
rect 25639 11645 25651 11648
rect 25593 11639 25651 11645
rect 19420 11611 19478 11617
rect 19420 11577 19432 11611
rect 19466 11608 19478 11611
rect 20806 11608 20812 11620
rect 19466 11580 20812 11608
rect 19466 11577 19478 11580
rect 19420 11571 19478 11577
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 21177 11611 21235 11617
rect 21177 11608 21189 11611
rect 20916 11580 21189 11608
rect 18748 11512 18920 11540
rect 18748 11500 18754 11512
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 20916 11540 20944 11580
rect 21177 11577 21189 11580
rect 21223 11608 21235 11611
rect 21560 11608 21588 11636
rect 21726 11617 21732 11620
rect 21720 11608 21732 11617
rect 21223 11580 21588 11608
rect 21687 11580 21732 11608
rect 21223 11577 21235 11580
rect 21177 11571 21235 11577
rect 21720 11571 21732 11580
rect 21726 11568 21732 11571
rect 21784 11568 21790 11620
rect 21818 11568 21824 11620
rect 21876 11608 21882 11620
rect 26206 11608 26234 11852
rect 28350 11840 28356 11852
rect 28408 11880 28414 11892
rect 28718 11880 28724 11892
rect 28408 11852 28724 11880
rect 28408 11840 28414 11852
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 30006 11840 30012 11892
rect 30064 11880 30070 11892
rect 30101 11883 30159 11889
rect 30101 11880 30113 11883
rect 30064 11852 30113 11880
rect 30064 11840 30070 11852
rect 30101 11849 30113 11852
rect 30147 11849 30159 11883
rect 30101 11843 30159 11849
rect 26786 11704 26792 11756
rect 26844 11744 26850 11756
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26844 11716 26985 11744
rect 26844 11704 26850 11716
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 28442 11704 28448 11756
rect 28500 11744 28506 11756
rect 30098 11744 30104 11756
rect 28500 11716 30104 11744
rect 28500 11704 28506 11716
rect 30024 11685 30052 11716
rect 30098 11704 30104 11716
rect 30156 11704 30162 11756
rect 26881 11679 26939 11685
rect 26881 11676 26893 11679
rect 21876 11580 26234 11608
rect 26712 11648 26893 11676
rect 21876 11568 21882 11580
rect 20680 11512 20944 11540
rect 20680 11500 20686 11512
rect 20990 11500 20996 11552
rect 21048 11500 21054 11552
rect 21082 11500 21088 11552
rect 21140 11500 21146 11552
rect 21361 11543 21419 11549
rect 21361 11509 21373 11543
rect 21407 11540 21419 11543
rect 22738 11540 22744 11552
rect 21407 11512 22744 11540
rect 21407 11509 21419 11512
rect 21361 11503 21419 11509
rect 22738 11500 22744 11512
rect 22796 11500 22802 11552
rect 26712 11540 26740 11648
rect 26881 11645 26893 11648
rect 26927 11645 26939 11679
rect 26881 11639 26939 11645
rect 30009 11679 30067 11685
rect 30009 11645 30021 11679
rect 30055 11645 30067 11679
rect 30009 11639 30067 11645
rect 26789 11611 26847 11617
rect 26789 11577 26801 11611
rect 26835 11608 26847 11611
rect 27249 11611 27307 11617
rect 27249 11608 27261 11611
rect 26835 11580 27261 11608
rect 26835 11577 26847 11580
rect 26789 11571 26847 11577
rect 27249 11577 27261 11580
rect 27295 11577 27307 11611
rect 28534 11608 28540 11620
rect 28474 11580 28540 11608
rect 27249 11571 27307 11577
rect 28534 11568 28540 11580
rect 28592 11568 28598 11620
rect 28258 11540 28264 11552
rect 26712 11512 28264 11540
rect 28258 11500 28264 11512
rect 28316 11540 28322 11552
rect 28721 11543 28779 11549
rect 28721 11540 28733 11543
rect 28316 11512 28733 11540
rect 28316 11500 28322 11512
rect 28721 11509 28733 11512
rect 28767 11509 28779 11543
rect 28721 11503 28779 11509
rect 552 11450 31808 11472
rect 552 11398 8172 11450
rect 8224 11398 8236 11450
rect 8288 11398 8300 11450
rect 8352 11398 8364 11450
rect 8416 11398 8428 11450
rect 8480 11398 15946 11450
rect 15998 11398 16010 11450
rect 16062 11398 16074 11450
rect 16126 11398 16138 11450
rect 16190 11398 16202 11450
rect 16254 11398 23720 11450
rect 23772 11398 23784 11450
rect 23836 11398 23848 11450
rect 23900 11398 23912 11450
rect 23964 11398 23976 11450
rect 24028 11398 31494 11450
rect 31546 11398 31558 11450
rect 31610 11398 31622 11450
rect 31674 11398 31686 11450
rect 31738 11398 31750 11450
rect 31802 11398 31808 11450
rect 552 11376 31808 11398
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 5077 11339 5135 11345
rect 5077 11336 5089 11339
rect 3476 11308 5089 11336
rect 3476 11296 3482 11308
rect 5077 11305 5089 11308
rect 5123 11336 5135 11339
rect 6270 11336 6276 11348
rect 5123 11308 6276 11336
rect 5123 11305 5135 11308
rect 5077 11299 5135 11305
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 7558 11296 7564 11348
rect 7616 11296 7622 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8934 11339 8992 11345
rect 8934 11336 8946 11339
rect 8628 11308 8946 11336
rect 8628 11296 8634 11308
rect 8934 11305 8946 11308
rect 8980 11305 8992 11339
rect 8934 11299 8992 11305
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 12897 11339 12955 11345
rect 12897 11305 12909 11339
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 13433 11339 13491 11345
rect 13433 11305 13445 11339
rect 13479 11336 13491 11339
rect 13814 11336 13820 11348
rect 13479 11308 13820 11336
rect 13479 11305 13491 11308
rect 13433 11299 13491 11305
rect 3436 11268 3464 11296
rect 5353 11271 5411 11277
rect 5353 11268 5365 11271
rect 2884 11240 3464 11268
rect 4830 11240 5365 11268
rect 2884 11209 2912 11240
rect 5353 11237 5365 11240
rect 5399 11237 5411 11271
rect 5353 11231 5411 11237
rect 5810 11228 5816 11280
rect 5868 11268 5874 11280
rect 6089 11271 6147 11277
rect 6089 11268 6101 11271
rect 5868 11240 6101 11268
rect 5868 11228 5874 11240
rect 6089 11237 6101 11240
rect 6135 11237 6147 11271
rect 6089 11231 6147 11237
rect 7098 11228 7104 11280
rect 7156 11228 7162 11280
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11169 2927 11203
rect 2869 11163 2927 11169
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 7576 11200 7604 11296
rect 8662 11228 8668 11280
rect 8720 11228 8726 11280
rect 9033 11271 9091 11277
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 10428 11268 10456 11296
rect 9079 11240 10456 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 12434 11228 12440 11280
rect 12492 11228 12498 11280
rect 12912 11268 12940 11299
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 15746 11296 15752 11348
rect 15804 11296 15810 11348
rect 16485 11339 16543 11345
rect 16485 11305 16497 11339
rect 16531 11336 16543 11339
rect 16761 11339 16819 11345
rect 16531 11308 16712 11336
rect 16531 11305 16543 11308
rect 16485 11299 16543 11305
rect 12912 11240 13400 11268
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 5491 11172 5764 11200
rect 7576 11172 7665 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 5736 11144 5764 11172
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 7653 11163 7711 11169
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11169 7895 11203
rect 8680 11200 8708 11228
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 8680 11172 8769 11200
rect 7837 11163 7895 11169
rect 8757 11169 8769 11172
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 8849 11203 8907 11209
rect 8849 11169 8861 11203
rect 8895 11200 8907 11203
rect 8938 11200 8944 11212
rect 8895 11172 8944 11200
rect 8895 11169 8907 11172
rect 8849 11163 8907 11169
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 3326 11092 3332 11144
rect 3384 11092 3390 11144
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 3436 11104 3617 11132
rect 3237 11067 3295 11073
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 3436 11064 3464 11104
rect 3605 11101 3617 11104
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 3752 11104 4660 11132
rect 3752 11092 3758 11104
rect 3283 11036 3464 11064
rect 4632 11064 4660 11104
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 6454 11132 6460 11144
rect 5859 11104 6460 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 5828 11064 5856 11095
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 7852 11132 7880 11163
rect 6604 11104 7880 11132
rect 8772 11132 8800 11163
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 11146 11160 11152 11212
rect 11204 11160 11210 11212
rect 13004 11209 13032 11240
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 13173 11203 13231 11209
rect 13035 11172 13069 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 13372 11200 13400 11240
rect 13630 11228 13636 11280
rect 13688 11228 13694 11280
rect 13722 11228 13728 11280
rect 13780 11228 13786 11280
rect 14826 11228 14832 11280
rect 14884 11228 14890 11280
rect 13740 11200 13768 11228
rect 13219 11172 13308 11200
rect 13372 11172 13768 11200
rect 15565 11203 15623 11209
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 11054 11132 11060 11144
rect 8772 11104 11060 11132
rect 6604 11092 6610 11104
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 4632 11036 5856 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 13280 11073 13308 11172
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 15654 11200 15660 11212
rect 15611 11172 15660 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 15580 11132 15608 11163
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 15764 11209 15792 11296
rect 16684 11277 16712 11308
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16850 11336 16856 11348
rect 16807 11308 16856 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 17092 11308 17509 11336
rect 17092 11296 17098 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 17497 11299 17555 11305
rect 17678 11296 17684 11348
rect 17736 11296 17742 11348
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 21542 11336 21548 11348
rect 21140 11308 21548 11336
rect 21140 11296 21146 11308
rect 21542 11296 21548 11308
rect 21600 11296 21606 11348
rect 21637 11339 21695 11345
rect 21637 11305 21649 11339
rect 21683 11336 21695 11339
rect 21726 11336 21732 11348
rect 21683 11308 21732 11336
rect 21683 11305 21695 11308
rect 21637 11299 21695 11305
rect 21726 11296 21732 11308
rect 21784 11336 21790 11348
rect 24305 11339 24363 11345
rect 21784 11308 23980 11336
rect 21784 11296 21790 11308
rect 16669 11271 16727 11277
rect 16669 11237 16681 11271
rect 16715 11237 16727 11271
rect 16669 11231 16727 11237
rect 17696 11209 17724 11296
rect 17954 11228 17960 11280
rect 18012 11268 18018 11280
rect 22005 11271 22063 11277
rect 22005 11268 22017 11271
rect 18012 11240 18276 11268
rect 18012 11228 18018 11240
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 16301 11203 16359 11209
rect 16301 11200 16313 11203
rect 15749 11163 15807 11169
rect 15948 11172 16313 11200
rect 13780 11104 15608 11132
rect 13780 11092 13786 11104
rect 15948 11073 15976 11172
rect 16301 11169 16313 11172
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 18046 11160 18052 11212
rect 18104 11160 18110 11212
rect 18248 11209 18276 11240
rect 20088 11240 22017 11268
rect 20088 11209 20116 11240
rect 22005 11237 22017 11240
rect 22051 11237 22063 11271
rect 22005 11231 22063 11237
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 20073 11203 20131 11209
rect 20073 11169 20085 11203
rect 20119 11169 20131 11203
rect 20073 11163 20131 11169
rect 20349 11203 20407 11209
rect 20349 11169 20361 11203
rect 20395 11200 20407 11203
rect 20622 11200 20628 11212
rect 20395 11172 20628 11200
rect 20395 11169 20407 11172
rect 20349 11163 20407 11169
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 20088 11132 20116 11163
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 21910 11200 21916 11212
rect 21499 11172 21916 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 21910 11160 21916 11172
rect 21968 11160 21974 11212
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11200 22155 11203
rect 22738 11200 22744 11212
rect 22143 11172 22744 11200
rect 22143 11169 22155 11172
rect 22097 11163 22155 11169
rect 22738 11160 22744 11172
rect 22796 11160 22802 11212
rect 23192 11203 23250 11209
rect 23192 11200 23204 11203
rect 22848 11172 23204 11200
rect 18003 11104 20116 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 22848 11132 22876 11172
rect 23192 11169 23204 11172
rect 23238 11200 23250 11203
rect 23474 11200 23480 11212
rect 23238 11172 23480 11200
rect 23238 11169 23250 11172
rect 23192 11163 23250 11169
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 21600 11104 22876 11132
rect 21600 11092 21606 11104
rect 22922 11092 22928 11144
rect 22980 11092 22986 11144
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 7248 11036 7573 11064
rect 7248 11024 7254 11036
rect 7561 11033 7573 11036
rect 7607 11033 7619 11067
rect 7561 11027 7619 11033
rect 13265 11067 13323 11073
rect 13265 11033 13277 11067
rect 13311 11064 13323 11067
rect 15933 11067 15991 11073
rect 13311 11036 14044 11064
rect 13311 11033 13323 11036
rect 13265 11027 13323 11033
rect 14016 11008 14044 11036
rect 15933 11033 15945 11067
rect 15979 11033 15991 11067
rect 15933 11027 15991 11033
rect 17865 11067 17923 11073
rect 17865 11033 17877 11067
rect 17911 11064 17923 11067
rect 18141 11067 18199 11073
rect 18141 11064 18153 11067
rect 17911 11036 18153 11064
rect 17911 11033 17923 11036
rect 17865 11027 17923 11033
rect 18141 11033 18153 11036
rect 18187 11033 18199 11067
rect 18141 11027 18199 11033
rect 20257 11067 20315 11073
rect 20257 11033 20269 11067
rect 20303 11064 20315 11067
rect 21269 11067 21327 11073
rect 21269 11064 21281 11067
rect 20303 11036 21281 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 21269 11033 21281 11036
rect 21315 11033 21327 11067
rect 21269 11027 21327 11033
rect 21821 11067 21879 11073
rect 21821 11033 21833 11067
rect 21867 11033 21879 11067
rect 23952 11064 23980 11308
rect 24305 11305 24317 11339
rect 24351 11336 24363 11339
rect 24762 11336 24768 11348
rect 24351 11308 24768 11336
rect 24351 11305 24363 11308
rect 24305 11299 24363 11305
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 28074 11296 28080 11348
rect 28132 11296 28138 11348
rect 28442 11296 28448 11348
rect 28500 11296 28506 11348
rect 28534 11296 28540 11348
rect 28592 11296 28598 11348
rect 24670 11228 24676 11280
rect 24728 11228 24734 11280
rect 27430 11228 27436 11280
rect 27488 11228 27494 11280
rect 28092 11268 28120 11296
rect 28092 11240 28212 11268
rect 24688 11200 24716 11228
rect 25225 11203 25283 11209
rect 25225 11200 25237 11203
rect 24688 11172 25237 11200
rect 25225 11169 25237 11172
rect 25271 11169 25283 11203
rect 25225 11163 25283 11169
rect 25406 11160 25412 11212
rect 25464 11160 25470 11212
rect 28184 11209 28212 11240
rect 25777 11203 25835 11209
rect 25777 11169 25789 11203
rect 25823 11169 25835 11203
rect 25777 11163 25835 11169
rect 28169 11203 28227 11209
rect 28169 11169 28181 11203
rect 28215 11169 28227 11203
rect 28460 11200 28488 11296
rect 28629 11203 28687 11209
rect 28629 11200 28641 11203
rect 28460 11172 28641 11200
rect 28169 11163 28227 11169
rect 28629 11169 28641 11172
rect 28675 11169 28687 11203
rect 28629 11163 28687 11169
rect 25317 11135 25375 11141
rect 25317 11101 25329 11135
rect 25363 11132 25375 11135
rect 25685 11135 25743 11141
rect 25685 11132 25697 11135
rect 25363 11104 25697 11132
rect 25363 11101 25375 11104
rect 25317 11095 25375 11101
rect 25685 11101 25697 11104
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 25792 11132 25820 11163
rect 26421 11135 26479 11141
rect 26421 11132 26433 11135
rect 25792 11104 26433 11132
rect 25792 11064 25820 11104
rect 26421 11101 26433 11104
rect 26467 11101 26479 11135
rect 27893 11135 27951 11141
rect 27893 11132 27905 11135
rect 26421 11095 26479 11101
rect 26896 11104 27905 11132
rect 23952 11036 25820 11064
rect 26145 11067 26203 11073
rect 21821 11027 21879 11033
rect 26145 11033 26157 11067
rect 26191 11064 26203 11067
rect 26896 11064 26924 11104
rect 27893 11101 27905 11104
rect 27939 11101 27951 11135
rect 28644 11132 28672 11163
rect 28718 11160 28724 11212
rect 28776 11200 28782 11212
rect 28905 11203 28963 11209
rect 28905 11200 28917 11203
rect 28776 11172 28917 11200
rect 28776 11160 28782 11172
rect 28905 11169 28917 11172
rect 28951 11169 28963 11203
rect 28905 11163 28963 11169
rect 29089 11135 29147 11141
rect 29089 11132 29101 11135
rect 28644 11104 29101 11132
rect 27893 11095 27951 11101
rect 29089 11101 29101 11104
rect 29135 11101 29147 11135
rect 29089 11095 29147 11101
rect 26191 11036 26924 11064
rect 26191 11033 26203 11036
rect 26145 11027 26203 11033
rect 7653 10999 7711 11005
rect 7653 10965 7665 10999
rect 7699 10996 7711 10999
rect 7742 10996 7748 11008
rect 7699 10968 7748 10996
rect 7699 10965 7711 10968
rect 7653 10959 7711 10965
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 13170 10956 13176 11008
rect 13228 10956 13234 11008
rect 13446 10956 13452 11008
rect 13504 10956 13510 11008
rect 13998 10956 14004 11008
rect 14056 10956 14062 11008
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 15301 10999 15359 11005
rect 15301 10996 15313 10999
rect 14148 10968 15313 10996
rect 14148 10956 14154 10968
rect 15301 10965 15313 10968
rect 15347 10965 15359 10999
rect 15301 10959 15359 10965
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19889 10999 19947 11005
rect 19889 10996 19901 10999
rect 19484 10968 19901 10996
rect 19484 10956 19490 10968
rect 19889 10965 19901 10968
rect 19935 10965 19947 10999
rect 19889 10959 19947 10965
rect 20806 10956 20812 11008
rect 20864 10996 20870 11008
rect 21726 10996 21732 11008
rect 20864 10968 21732 10996
rect 20864 10956 20870 10968
rect 21726 10956 21732 10968
rect 21784 10996 21790 11008
rect 21836 10996 21864 11027
rect 21784 10968 21864 10996
rect 21784 10956 21790 10968
rect 552 10906 31648 10928
rect 552 10854 4285 10906
rect 4337 10854 4349 10906
rect 4401 10854 4413 10906
rect 4465 10854 4477 10906
rect 4529 10854 4541 10906
rect 4593 10854 12059 10906
rect 12111 10854 12123 10906
rect 12175 10854 12187 10906
rect 12239 10854 12251 10906
rect 12303 10854 12315 10906
rect 12367 10854 19833 10906
rect 19885 10854 19897 10906
rect 19949 10854 19961 10906
rect 20013 10854 20025 10906
rect 20077 10854 20089 10906
rect 20141 10854 27607 10906
rect 27659 10854 27671 10906
rect 27723 10854 27735 10906
rect 27787 10854 27799 10906
rect 27851 10854 27863 10906
rect 27915 10854 31648 10906
rect 552 10832 31648 10854
rect 6181 10795 6239 10801
rect 6181 10761 6193 10795
rect 6227 10792 6239 10795
rect 7098 10792 7104 10804
rect 6227 10764 7104 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7524 10764 8217 10792
rect 7524 10752 7530 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11609 10795 11667 10801
rect 11609 10792 11621 10795
rect 11480 10764 11621 10792
rect 11480 10752 11486 10764
rect 11609 10761 11621 10764
rect 11655 10761 11667 10795
rect 11609 10755 11667 10761
rect 12161 10795 12219 10801
rect 12161 10761 12173 10795
rect 12207 10792 12219 10795
rect 12434 10792 12440 10804
rect 12207 10764 12440 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 12434 10752 12440 10764
rect 12492 10752 12498 10804
rect 14090 10752 14096 10804
rect 14148 10752 14154 10804
rect 14826 10752 14832 10804
rect 14884 10752 14890 10804
rect 20533 10795 20591 10801
rect 20533 10761 20545 10795
rect 20579 10792 20591 10795
rect 20622 10792 20628 10804
rect 20579 10764 20628 10792
rect 20579 10761 20591 10764
rect 20533 10755 20591 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 23474 10752 23480 10804
rect 23532 10752 23538 10804
rect 25406 10752 25412 10804
rect 25464 10792 25470 10804
rect 25685 10795 25743 10801
rect 25685 10792 25697 10795
rect 25464 10764 25697 10792
rect 25464 10752 25470 10764
rect 25685 10761 25697 10764
rect 25731 10761 25743 10795
rect 25685 10755 25743 10761
rect 27430 10752 27436 10804
rect 27488 10752 27494 10804
rect 13817 10727 13875 10733
rect 13817 10693 13829 10727
rect 13863 10693 13875 10727
rect 13817 10687 13875 10693
rect 6454 10616 6460 10668
rect 6512 10616 6518 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7742 10656 7748 10668
rect 6779 10628 7748 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 8662 10616 8668 10668
rect 8720 10656 8726 10668
rect 8849 10659 8907 10665
rect 8849 10656 8861 10659
rect 8720 10628 8861 10656
rect 8720 10616 8726 10628
rect 8849 10625 8861 10628
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 9355 10628 9689 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 11974 10656 11980 10668
rect 9677 10619 9735 10625
rect 10704 10628 11980 10656
rect 10704 10600 10732 10628
rect 11974 10616 11980 10628
rect 12032 10656 12038 10668
rect 12032 10628 13676 10656
rect 12032 10616 12038 10628
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 6089 10591 6147 10597
rect 6089 10588 6101 10591
rect 5776 10560 6101 10588
rect 5776 10548 5782 10560
rect 6089 10557 6101 10560
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 6104 10520 6132 10551
rect 8481 10523 8539 10529
rect 8481 10520 8493 10523
rect 6104 10492 6914 10520
rect 7958 10492 8493 10520
rect 6886 10452 6914 10492
rect 8481 10489 8493 10492
rect 8527 10489 8539 10523
rect 8481 10483 8539 10489
rect 8588 10464 8616 10551
rect 8938 10548 8944 10600
rect 8996 10548 9002 10600
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 10686 10548 10692 10600
rect 10744 10548 10750 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 12084 10597 12112 10628
rect 11425 10591 11483 10597
rect 11425 10588 11437 10591
rect 11112 10560 11437 10588
rect 11112 10548 11118 10560
rect 11425 10557 11437 10560
rect 11471 10557 11483 10591
rect 11425 10551 11483 10557
rect 11609 10591 11667 10597
rect 11609 10557 11621 10591
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 8570 10452 8576 10464
rect 6886 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 8956 10452 8984 10548
rect 10410 10480 10416 10532
rect 10468 10480 10474 10532
rect 11624 10520 11652 10551
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13541 10591 13599 10597
rect 13541 10588 13553 10591
rect 13504 10560 13553 10588
rect 13504 10548 13510 10560
rect 13541 10557 13553 10560
rect 13587 10557 13599 10591
rect 13541 10551 13599 10557
rect 13170 10520 13176 10532
rect 11624 10492 13176 10520
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 13648 10520 13676 10628
rect 13832 10588 13860 10687
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 19061 10659 19119 10665
rect 16448 10628 18828 10656
rect 16448 10616 16454 10628
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13832 10560 13921 10588
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 18800 10597 18828 10628
rect 19061 10625 19073 10659
rect 19107 10656 19119 10659
rect 19426 10656 19432 10668
rect 19107 10628 19432 10656
rect 19107 10625 19119 10628
rect 19061 10619 19119 10625
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 21174 10616 21180 10668
rect 21232 10616 21238 10668
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10656 21695 10659
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21683 10628 22017 10656
rect 21683 10625 21695 10628
rect 21637 10619 21695 10625
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 23937 10659 23995 10665
rect 23937 10625 23949 10659
rect 23983 10656 23995 10659
rect 24302 10656 24308 10668
rect 23983 10628 24308 10656
rect 23983 10625 23995 10628
rect 23937 10619 23995 10625
rect 24302 10616 24308 10628
rect 24360 10616 24366 10668
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 14056 10560 14105 10588
rect 14056 10548 14062 10560
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10557 14979 10591
rect 14921 10551 14979 10557
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 18785 10591 18843 10597
rect 18555 10560 18736 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 13648 10492 13768 10520
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 8956 10424 11161 10452
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 13630 10412 13636 10464
rect 13688 10412 13694 10464
rect 13740 10452 13768 10492
rect 13814 10480 13820 10532
rect 13872 10480 13878 10532
rect 14936 10452 14964 10551
rect 18708 10532 18736 10560
rect 18785 10557 18797 10591
rect 18831 10557 18843 10591
rect 18785 10551 18843 10557
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 21542 10588 21548 10600
rect 21315 10560 21548 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 16666 10480 16672 10532
rect 16724 10480 16730 10532
rect 18417 10523 18475 10529
rect 18417 10520 18429 10523
rect 17894 10492 18429 10520
rect 18417 10489 18429 10492
rect 18463 10489 18475 10523
rect 18417 10483 18475 10489
rect 18690 10480 18696 10532
rect 18748 10480 18754 10532
rect 15194 10452 15200 10464
rect 13740 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 18046 10452 18052 10464
rect 17736 10424 18052 10452
rect 17736 10412 17742 10424
rect 18046 10412 18052 10424
rect 18104 10452 18110 10464
rect 18141 10455 18199 10461
rect 18141 10452 18153 10455
rect 18104 10424 18153 10452
rect 18104 10412 18110 10424
rect 18141 10421 18153 10424
rect 18187 10421 18199 10455
rect 18800 10452 18828 10551
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 21729 10591 21787 10597
rect 21729 10557 21741 10591
rect 21775 10557 21787 10591
rect 21729 10551 21787 10557
rect 19794 10480 19800 10532
rect 19852 10480 19858 10532
rect 20346 10452 20352 10464
rect 18800 10424 20352 10452
rect 18141 10415 18199 10421
rect 20346 10412 20352 10424
rect 20404 10452 20410 10464
rect 21744 10452 21772 10551
rect 25682 10548 25688 10600
rect 25740 10588 25746 10600
rect 26053 10591 26111 10597
rect 26053 10588 26065 10591
rect 25740 10560 26065 10588
rect 25740 10548 25746 10560
rect 26053 10557 26065 10560
rect 26099 10588 26111 10591
rect 27525 10591 27583 10597
rect 27525 10588 27537 10591
rect 26099 10560 27537 10588
rect 26099 10557 26111 10560
rect 26053 10551 26111 10557
rect 27525 10557 27537 10560
rect 27571 10557 27583 10591
rect 27525 10551 27583 10557
rect 23014 10480 23020 10532
rect 23072 10480 23078 10532
rect 24210 10480 24216 10532
rect 24268 10480 24274 10532
rect 25961 10523 26019 10529
rect 25961 10520 25973 10523
rect 25438 10492 25973 10520
rect 25961 10489 25973 10492
rect 26007 10489 26019 10523
rect 25961 10483 26019 10489
rect 20404 10424 21772 10452
rect 20404 10412 20410 10424
rect 552 10362 31808 10384
rect 552 10310 8172 10362
rect 8224 10310 8236 10362
rect 8288 10310 8300 10362
rect 8352 10310 8364 10362
rect 8416 10310 8428 10362
rect 8480 10310 15946 10362
rect 15998 10310 16010 10362
rect 16062 10310 16074 10362
rect 16126 10310 16138 10362
rect 16190 10310 16202 10362
rect 16254 10310 23720 10362
rect 23772 10310 23784 10362
rect 23836 10310 23848 10362
rect 23900 10310 23912 10362
rect 23964 10310 23976 10362
rect 24028 10310 31494 10362
rect 31546 10310 31558 10362
rect 31610 10310 31622 10362
rect 31674 10310 31686 10362
rect 31738 10310 31750 10362
rect 31802 10310 31808 10362
rect 552 10288 31808 10310
rect 8570 10208 8576 10260
rect 8628 10208 8634 10260
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 10505 10251 10563 10257
rect 10505 10248 10517 10251
rect 10468 10220 10517 10248
rect 10468 10208 10474 10220
rect 10505 10217 10517 10220
rect 10551 10217 10563 10251
rect 10505 10211 10563 10217
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 13722 10248 13728 10260
rect 11204 10220 13728 10248
rect 11204 10208 11210 10220
rect 8588 10112 8616 10208
rect 10413 10115 10471 10121
rect 10413 10112 10425 10115
rect 8588 10084 10425 10112
rect 10413 10081 10425 10084
rect 10459 10112 10471 10115
rect 10502 10112 10508 10124
rect 10459 10084 10508 10112
rect 10459 10081 10471 10084
rect 10413 10075 10471 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 11256 10121 11284 10220
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15381 10251 15439 10257
rect 15381 10248 15393 10251
rect 15344 10220 15393 10248
rect 15344 10208 15350 10220
rect 15381 10217 15393 10220
rect 15427 10217 15439 10251
rect 15381 10211 15439 10217
rect 16666 10208 16672 10260
rect 16724 10208 16730 10260
rect 19794 10208 19800 10260
rect 19852 10208 19858 10260
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 21232 10220 21281 10248
rect 21232 10208 21238 10220
rect 21269 10217 21281 10220
rect 21315 10217 21327 10251
rect 22002 10248 22008 10260
rect 21269 10211 21327 10217
rect 21376 10220 22008 10248
rect 12526 10140 12532 10192
rect 12584 10140 12590 10192
rect 13265 10183 13323 10189
rect 13265 10149 13277 10183
rect 13311 10180 13323 10183
rect 13446 10180 13452 10192
rect 13311 10152 13452 10180
rect 13311 10149 13323 10152
rect 13265 10143 13323 10149
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 13740 10180 13768 10208
rect 15657 10183 15715 10189
rect 15657 10180 15669 10183
rect 13648 10152 13768 10180
rect 15134 10152 15669 10180
rect 13648 10121 13676 10152
rect 15657 10149 15669 10152
rect 15703 10149 15715 10183
rect 15657 10143 15715 10149
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 15565 10115 15623 10121
rect 15565 10112 15577 10115
rect 15252 10084 15577 10112
rect 15252 10072 15258 10084
rect 15565 10081 15577 10084
rect 15611 10081 15623 10115
rect 15565 10075 15623 10081
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 13906 10004 13912 10056
rect 13964 10004 13970 10056
rect 16684 10044 16712 10208
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 17865 10183 17923 10189
rect 17865 10180 17877 10183
rect 16908 10152 17877 10180
rect 16908 10140 16914 10152
rect 17865 10149 17877 10152
rect 17911 10149 17923 10183
rect 17865 10143 17923 10149
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10112 17187 10115
rect 17678 10112 17684 10124
rect 17175 10084 17684 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 18690 10072 18696 10124
rect 18748 10112 18754 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 18748 10084 19717 10112
rect 18748 10072 18754 10084
rect 19705 10081 19717 10084
rect 19751 10112 19763 10115
rect 21376 10112 21404 10220
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22925 10251 22983 10257
rect 22925 10217 22937 10251
rect 22971 10248 22983 10251
rect 23014 10248 23020 10260
rect 22971 10220 23020 10248
rect 22971 10217 22983 10220
rect 22925 10211 22983 10217
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 24210 10208 24216 10260
rect 24268 10208 24274 10260
rect 21437 10183 21495 10189
rect 21437 10149 21449 10183
rect 21483 10180 21495 10183
rect 21637 10183 21695 10189
rect 21483 10152 21588 10180
rect 21483 10149 21495 10152
rect 21437 10143 21495 10149
rect 19751 10084 21404 10112
rect 21560 10112 21588 10152
rect 21637 10149 21649 10183
rect 21683 10180 21695 10183
rect 21726 10180 21732 10192
rect 21683 10152 21732 10180
rect 21683 10149 21695 10152
rect 21637 10143 21695 10149
rect 21726 10140 21732 10152
rect 21784 10180 21790 10192
rect 21784 10152 23612 10180
rect 21784 10140 21790 10152
rect 21560 10084 21956 10112
rect 19751 10081 19763 10084
rect 19705 10075 19763 10081
rect 16761 10047 16819 10053
rect 16761 10044 16773 10047
rect 16684 10016 16773 10044
rect 16761 10013 16773 10016
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 17218 10004 17224 10056
rect 17276 10004 17282 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 18708 10044 18736 10072
rect 21928 10056 21956 10084
rect 22002 10072 22008 10124
rect 22060 10112 22066 10124
rect 23584 10121 23612 10152
rect 22833 10115 22891 10121
rect 22833 10112 22845 10115
rect 22060 10084 22845 10112
rect 22060 10072 22066 10084
rect 22833 10081 22845 10084
rect 22879 10081 22891 10115
rect 22833 10075 22891 10081
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10081 23627 10115
rect 23569 10075 23627 10081
rect 17635 10016 18736 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 21910 10004 21916 10056
rect 21968 10044 21974 10056
rect 23477 10047 23535 10053
rect 23477 10044 23489 10047
rect 21968 10016 23489 10044
rect 21968 10004 21974 10016
rect 23477 10013 23489 10016
rect 23523 10013 23535 10047
rect 23477 10007 23535 10013
rect 23584 9976 23612 10075
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10044 23995 10047
rect 24228 10044 24256 10208
rect 23983 10016 24256 10044
rect 23983 10013 23995 10016
rect 23937 10007 23995 10013
rect 25406 9976 25412 9988
rect 23584 9948 25412 9976
rect 25406 9936 25412 9948
rect 25464 9936 25470 9988
rect 21453 9911 21511 9917
rect 21453 9877 21465 9911
rect 21499 9908 21511 9911
rect 21634 9908 21640 9920
rect 21499 9880 21640 9908
rect 21499 9877 21511 9880
rect 21453 9871 21511 9877
rect 21634 9868 21640 9880
rect 21692 9868 21698 9920
rect 552 9818 31648 9840
rect 552 9766 4285 9818
rect 4337 9766 4349 9818
rect 4401 9766 4413 9818
rect 4465 9766 4477 9818
rect 4529 9766 4541 9818
rect 4593 9766 12059 9818
rect 12111 9766 12123 9818
rect 12175 9766 12187 9818
rect 12239 9766 12251 9818
rect 12303 9766 12315 9818
rect 12367 9766 19833 9818
rect 19885 9766 19897 9818
rect 19949 9766 19961 9818
rect 20013 9766 20025 9818
rect 20077 9766 20089 9818
rect 20141 9766 27607 9818
rect 27659 9766 27671 9818
rect 27723 9766 27735 9818
rect 27787 9766 27799 9818
rect 27851 9766 27863 9818
rect 27915 9766 31648 9818
rect 552 9744 31648 9766
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 11977 9707 12035 9713
rect 11977 9704 11989 9707
rect 11572 9676 11989 9704
rect 11572 9664 11578 9676
rect 11977 9673 11989 9676
rect 12023 9673 12035 9707
rect 11977 9667 12035 9673
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 14093 9707 14151 9713
rect 14093 9704 14105 9707
rect 13964 9676 14105 9704
rect 13964 9664 13970 9676
rect 14093 9673 14105 9676
rect 14139 9673 14151 9707
rect 14093 9667 14151 9673
rect 12345 9639 12403 9645
rect 12345 9605 12357 9639
rect 12391 9636 12403 9639
rect 12526 9636 12532 9648
rect 12391 9608 12532 9636
rect 12391 9605 12403 9608
rect 12345 9599 12403 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 13446 9568 13452 9580
rect 12084 9540 13452 9568
rect 11992 9432 12020 9528
rect 12084 9509 12112 9540
rect 13446 9528 13452 9540
rect 13504 9568 13510 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13504 9540 13829 9568
rect 13504 9528 13510 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 12069 9503 12127 9509
rect 12069 9469 12081 9503
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12268 9432 12296 9463
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13688 9472 13737 9500
rect 13688 9460 13694 9472
rect 13725 9469 13737 9472
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 11992 9404 12296 9432
rect 552 9274 31808 9296
rect 552 9222 8172 9274
rect 8224 9222 8236 9274
rect 8288 9222 8300 9274
rect 8352 9222 8364 9274
rect 8416 9222 8428 9274
rect 8480 9222 15946 9274
rect 15998 9222 16010 9274
rect 16062 9222 16074 9274
rect 16126 9222 16138 9274
rect 16190 9222 16202 9274
rect 16254 9222 23720 9274
rect 23772 9222 23784 9274
rect 23836 9222 23848 9274
rect 23900 9222 23912 9274
rect 23964 9222 23976 9274
rect 24028 9222 31494 9274
rect 31546 9222 31558 9274
rect 31610 9222 31622 9274
rect 31674 9222 31686 9274
rect 31738 9222 31750 9274
rect 31802 9222 31808 9274
rect 552 9200 31808 9222
rect 552 8730 31648 8752
rect 552 8678 4285 8730
rect 4337 8678 4349 8730
rect 4401 8678 4413 8730
rect 4465 8678 4477 8730
rect 4529 8678 4541 8730
rect 4593 8678 12059 8730
rect 12111 8678 12123 8730
rect 12175 8678 12187 8730
rect 12239 8678 12251 8730
rect 12303 8678 12315 8730
rect 12367 8678 19833 8730
rect 19885 8678 19897 8730
rect 19949 8678 19961 8730
rect 20013 8678 20025 8730
rect 20077 8678 20089 8730
rect 20141 8678 27607 8730
rect 27659 8678 27671 8730
rect 27723 8678 27735 8730
rect 27787 8678 27799 8730
rect 27851 8678 27863 8730
rect 27915 8678 31648 8730
rect 552 8656 31648 8678
rect 552 8186 31808 8208
rect 552 8134 8172 8186
rect 8224 8134 8236 8186
rect 8288 8134 8300 8186
rect 8352 8134 8364 8186
rect 8416 8134 8428 8186
rect 8480 8134 15946 8186
rect 15998 8134 16010 8186
rect 16062 8134 16074 8186
rect 16126 8134 16138 8186
rect 16190 8134 16202 8186
rect 16254 8134 23720 8186
rect 23772 8134 23784 8186
rect 23836 8134 23848 8186
rect 23900 8134 23912 8186
rect 23964 8134 23976 8186
rect 24028 8134 31494 8186
rect 31546 8134 31558 8186
rect 31610 8134 31622 8186
rect 31674 8134 31686 8186
rect 31738 8134 31750 8186
rect 31802 8134 31808 8186
rect 552 8112 31808 8134
rect 552 7642 31648 7664
rect 552 7590 4285 7642
rect 4337 7590 4349 7642
rect 4401 7590 4413 7642
rect 4465 7590 4477 7642
rect 4529 7590 4541 7642
rect 4593 7590 12059 7642
rect 12111 7590 12123 7642
rect 12175 7590 12187 7642
rect 12239 7590 12251 7642
rect 12303 7590 12315 7642
rect 12367 7590 19833 7642
rect 19885 7590 19897 7642
rect 19949 7590 19961 7642
rect 20013 7590 20025 7642
rect 20077 7590 20089 7642
rect 20141 7590 27607 7642
rect 27659 7590 27671 7642
rect 27723 7590 27735 7642
rect 27787 7590 27799 7642
rect 27851 7590 27863 7642
rect 27915 7590 31648 7642
rect 552 7568 31648 7590
rect 552 7098 31808 7120
rect 552 7046 8172 7098
rect 8224 7046 8236 7098
rect 8288 7046 8300 7098
rect 8352 7046 8364 7098
rect 8416 7046 8428 7098
rect 8480 7046 15946 7098
rect 15998 7046 16010 7098
rect 16062 7046 16074 7098
rect 16126 7046 16138 7098
rect 16190 7046 16202 7098
rect 16254 7046 23720 7098
rect 23772 7046 23784 7098
rect 23836 7046 23848 7098
rect 23900 7046 23912 7098
rect 23964 7046 23976 7098
rect 24028 7046 31494 7098
rect 31546 7046 31558 7098
rect 31610 7046 31622 7098
rect 31674 7046 31686 7098
rect 31738 7046 31750 7098
rect 31802 7046 31808 7098
rect 552 7024 31808 7046
rect 552 6554 31648 6576
rect 552 6502 4285 6554
rect 4337 6502 4349 6554
rect 4401 6502 4413 6554
rect 4465 6502 4477 6554
rect 4529 6502 4541 6554
rect 4593 6502 12059 6554
rect 12111 6502 12123 6554
rect 12175 6502 12187 6554
rect 12239 6502 12251 6554
rect 12303 6502 12315 6554
rect 12367 6502 19833 6554
rect 19885 6502 19897 6554
rect 19949 6502 19961 6554
rect 20013 6502 20025 6554
rect 20077 6502 20089 6554
rect 20141 6502 27607 6554
rect 27659 6502 27671 6554
rect 27723 6502 27735 6554
rect 27787 6502 27799 6554
rect 27851 6502 27863 6554
rect 27915 6502 31648 6554
rect 552 6480 31648 6502
rect 552 6010 31808 6032
rect 552 5958 8172 6010
rect 8224 5958 8236 6010
rect 8288 5958 8300 6010
rect 8352 5958 8364 6010
rect 8416 5958 8428 6010
rect 8480 5958 15946 6010
rect 15998 5958 16010 6010
rect 16062 5958 16074 6010
rect 16126 5958 16138 6010
rect 16190 5958 16202 6010
rect 16254 5958 23720 6010
rect 23772 5958 23784 6010
rect 23836 5958 23848 6010
rect 23900 5958 23912 6010
rect 23964 5958 23976 6010
rect 24028 5958 31494 6010
rect 31546 5958 31558 6010
rect 31610 5958 31622 6010
rect 31674 5958 31686 6010
rect 31738 5958 31750 6010
rect 31802 5958 31808 6010
rect 552 5936 31808 5958
rect 552 5466 31648 5488
rect 552 5414 4285 5466
rect 4337 5414 4349 5466
rect 4401 5414 4413 5466
rect 4465 5414 4477 5466
rect 4529 5414 4541 5466
rect 4593 5414 12059 5466
rect 12111 5414 12123 5466
rect 12175 5414 12187 5466
rect 12239 5414 12251 5466
rect 12303 5414 12315 5466
rect 12367 5414 19833 5466
rect 19885 5414 19897 5466
rect 19949 5414 19961 5466
rect 20013 5414 20025 5466
rect 20077 5414 20089 5466
rect 20141 5414 27607 5466
rect 27659 5414 27671 5466
rect 27723 5414 27735 5466
rect 27787 5414 27799 5466
rect 27851 5414 27863 5466
rect 27915 5414 31648 5466
rect 552 5392 31648 5414
rect 552 4922 31808 4944
rect 552 4870 8172 4922
rect 8224 4870 8236 4922
rect 8288 4870 8300 4922
rect 8352 4870 8364 4922
rect 8416 4870 8428 4922
rect 8480 4870 15946 4922
rect 15998 4870 16010 4922
rect 16062 4870 16074 4922
rect 16126 4870 16138 4922
rect 16190 4870 16202 4922
rect 16254 4870 23720 4922
rect 23772 4870 23784 4922
rect 23836 4870 23848 4922
rect 23900 4870 23912 4922
rect 23964 4870 23976 4922
rect 24028 4870 31494 4922
rect 31546 4870 31558 4922
rect 31610 4870 31622 4922
rect 31674 4870 31686 4922
rect 31738 4870 31750 4922
rect 31802 4870 31808 4922
rect 552 4848 31808 4870
rect 552 4378 31648 4400
rect 552 4326 4285 4378
rect 4337 4326 4349 4378
rect 4401 4326 4413 4378
rect 4465 4326 4477 4378
rect 4529 4326 4541 4378
rect 4593 4326 12059 4378
rect 12111 4326 12123 4378
rect 12175 4326 12187 4378
rect 12239 4326 12251 4378
rect 12303 4326 12315 4378
rect 12367 4326 19833 4378
rect 19885 4326 19897 4378
rect 19949 4326 19961 4378
rect 20013 4326 20025 4378
rect 20077 4326 20089 4378
rect 20141 4326 27607 4378
rect 27659 4326 27671 4378
rect 27723 4326 27735 4378
rect 27787 4326 27799 4378
rect 27851 4326 27863 4378
rect 27915 4326 31648 4378
rect 552 4304 31648 4326
rect 552 3834 31808 3856
rect 552 3782 8172 3834
rect 8224 3782 8236 3834
rect 8288 3782 8300 3834
rect 8352 3782 8364 3834
rect 8416 3782 8428 3834
rect 8480 3782 15946 3834
rect 15998 3782 16010 3834
rect 16062 3782 16074 3834
rect 16126 3782 16138 3834
rect 16190 3782 16202 3834
rect 16254 3782 23720 3834
rect 23772 3782 23784 3834
rect 23836 3782 23848 3834
rect 23900 3782 23912 3834
rect 23964 3782 23976 3834
rect 24028 3782 31494 3834
rect 31546 3782 31558 3834
rect 31610 3782 31622 3834
rect 31674 3782 31686 3834
rect 31738 3782 31750 3834
rect 31802 3782 31808 3834
rect 552 3760 31808 3782
rect 552 3290 31648 3312
rect 552 3238 4285 3290
rect 4337 3238 4349 3290
rect 4401 3238 4413 3290
rect 4465 3238 4477 3290
rect 4529 3238 4541 3290
rect 4593 3238 12059 3290
rect 12111 3238 12123 3290
rect 12175 3238 12187 3290
rect 12239 3238 12251 3290
rect 12303 3238 12315 3290
rect 12367 3238 19833 3290
rect 19885 3238 19897 3290
rect 19949 3238 19961 3290
rect 20013 3238 20025 3290
rect 20077 3238 20089 3290
rect 20141 3238 27607 3290
rect 27659 3238 27671 3290
rect 27723 3238 27735 3290
rect 27787 3238 27799 3290
rect 27851 3238 27863 3290
rect 27915 3238 31648 3290
rect 552 3216 31648 3238
rect 552 2746 31808 2768
rect 552 2694 8172 2746
rect 8224 2694 8236 2746
rect 8288 2694 8300 2746
rect 8352 2694 8364 2746
rect 8416 2694 8428 2746
rect 8480 2694 15946 2746
rect 15998 2694 16010 2746
rect 16062 2694 16074 2746
rect 16126 2694 16138 2746
rect 16190 2694 16202 2746
rect 16254 2694 23720 2746
rect 23772 2694 23784 2746
rect 23836 2694 23848 2746
rect 23900 2694 23912 2746
rect 23964 2694 23976 2746
rect 24028 2694 31494 2746
rect 31546 2694 31558 2746
rect 31610 2694 31622 2746
rect 31674 2694 31686 2746
rect 31738 2694 31750 2746
rect 31802 2694 31808 2746
rect 552 2672 31808 2694
rect 552 2202 31648 2224
rect 552 2150 4285 2202
rect 4337 2150 4349 2202
rect 4401 2150 4413 2202
rect 4465 2150 4477 2202
rect 4529 2150 4541 2202
rect 4593 2150 12059 2202
rect 12111 2150 12123 2202
rect 12175 2150 12187 2202
rect 12239 2150 12251 2202
rect 12303 2150 12315 2202
rect 12367 2150 19833 2202
rect 19885 2150 19897 2202
rect 19949 2150 19961 2202
rect 20013 2150 20025 2202
rect 20077 2150 20089 2202
rect 20141 2150 27607 2202
rect 27659 2150 27671 2202
rect 27723 2150 27735 2202
rect 27787 2150 27799 2202
rect 27851 2150 27863 2202
rect 27915 2150 31648 2202
rect 552 2128 31648 2150
rect 552 1658 31808 1680
rect 552 1606 8172 1658
rect 8224 1606 8236 1658
rect 8288 1606 8300 1658
rect 8352 1606 8364 1658
rect 8416 1606 8428 1658
rect 8480 1606 15946 1658
rect 15998 1606 16010 1658
rect 16062 1606 16074 1658
rect 16126 1606 16138 1658
rect 16190 1606 16202 1658
rect 16254 1606 23720 1658
rect 23772 1606 23784 1658
rect 23836 1606 23848 1658
rect 23900 1606 23912 1658
rect 23964 1606 23976 1658
rect 24028 1606 31494 1658
rect 31546 1606 31558 1658
rect 31610 1606 31622 1658
rect 31674 1606 31686 1658
rect 31738 1606 31750 1658
rect 31802 1606 31808 1658
rect 552 1584 31808 1606
rect 552 1114 31648 1136
rect 552 1062 4285 1114
rect 4337 1062 4349 1114
rect 4401 1062 4413 1114
rect 4465 1062 4477 1114
rect 4529 1062 4541 1114
rect 4593 1062 12059 1114
rect 12111 1062 12123 1114
rect 12175 1062 12187 1114
rect 12239 1062 12251 1114
rect 12303 1062 12315 1114
rect 12367 1062 19833 1114
rect 19885 1062 19897 1114
rect 19949 1062 19961 1114
rect 20013 1062 20025 1114
rect 20077 1062 20089 1114
rect 20141 1062 27607 1114
rect 27659 1062 27671 1114
rect 27723 1062 27735 1114
rect 27787 1062 27799 1114
rect 27851 1062 27863 1114
rect 27915 1062 31648 1114
rect 552 1040 31648 1062
rect 552 570 31808 592
rect 552 518 8172 570
rect 8224 518 8236 570
rect 8288 518 8300 570
rect 8352 518 8364 570
rect 8416 518 8428 570
rect 8480 518 15946 570
rect 15998 518 16010 570
rect 16062 518 16074 570
rect 16126 518 16138 570
rect 16190 518 16202 570
rect 16254 518 23720 570
rect 23772 518 23784 570
rect 23836 518 23848 570
rect 23900 518 23912 570
rect 23964 518 23976 570
rect 24028 518 31494 570
rect 31546 518 31558 570
rect 31610 518 31622 570
rect 31674 518 31686 570
rect 31738 518 31750 570
rect 31802 518 31808 570
rect 552 496 31808 518
<< via1 >>
rect 16304 21836 16356 21888
rect 23940 21836 23992 21888
rect 29368 21836 29420 21888
rect 4285 21734 4337 21786
rect 4349 21734 4401 21786
rect 4413 21734 4465 21786
rect 4477 21734 4529 21786
rect 4541 21734 4593 21786
rect 12059 21734 12111 21786
rect 12123 21734 12175 21786
rect 12187 21734 12239 21786
rect 12251 21734 12303 21786
rect 12315 21734 12367 21786
rect 19833 21734 19885 21786
rect 19897 21734 19949 21786
rect 19961 21734 20013 21786
rect 20025 21734 20077 21786
rect 20089 21734 20141 21786
rect 27607 21734 27659 21786
rect 27671 21734 27723 21786
rect 27735 21734 27787 21786
rect 27799 21734 27851 21786
rect 27863 21734 27915 21786
rect 848 21675 900 21684
rect 848 21641 857 21675
rect 857 21641 891 21675
rect 891 21641 900 21675
rect 848 21632 900 21641
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2320 21675 2372 21684
rect 2320 21641 2329 21675
rect 2329 21641 2363 21675
rect 2363 21641 2372 21675
rect 2320 21632 2372 21641
rect 3240 21675 3292 21684
rect 3240 21641 3249 21675
rect 3249 21641 3283 21675
rect 3283 21641 3292 21675
rect 3240 21632 3292 21641
rect 3792 21675 3844 21684
rect 3792 21641 3801 21675
rect 3801 21641 3835 21675
rect 3835 21641 3844 21675
rect 3792 21632 3844 21641
rect 4620 21632 4672 21684
rect 5264 21675 5316 21684
rect 5264 21641 5273 21675
rect 5273 21641 5307 21675
rect 5307 21641 5316 21675
rect 5264 21632 5316 21641
rect 6000 21675 6052 21684
rect 6000 21641 6009 21675
rect 6009 21641 6043 21675
rect 6043 21641 6052 21675
rect 6000 21632 6052 21641
rect 6736 21675 6788 21684
rect 6736 21641 6745 21675
rect 6745 21641 6779 21675
rect 6779 21641 6788 21675
rect 6736 21632 6788 21641
rect 7472 21675 7524 21684
rect 7472 21641 7481 21675
rect 7481 21641 7515 21675
rect 7515 21641 7524 21675
rect 7472 21632 7524 21641
rect 8208 21675 8260 21684
rect 8208 21641 8217 21675
rect 8217 21641 8251 21675
rect 8251 21641 8260 21675
rect 8208 21632 8260 21641
rect 8760 21675 8812 21684
rect 8760 21641 8769 21675
rect 8769 21641 8803 21675
rect 8803 21641 8812 21675
rect 8760 21632 8812 21641
rect 9680 21675 9732 21684
rect 9680 21641 9689 21675
rect 9689 21641 9723 21675
rect 9723 21641 9732 21675
rect 9680 21632 9732 21641
rect 10416 21675 10468 21684
rect 10416 21641 10425 21675
rect 10425 21641 10459 21675
rect 10459 21641 10468 21675
rect 10416 21632 10468 21641
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 16304 21632 16356 21684
rect 23940 21632 23992 21684
rect 6644 21428 6696 21480
rect 11520 21471 11572 21480
rect 11520 21437 11529 21471
rect 11529 21437 11563 21471
rect 11563 21437 11572 21471
rect 14648 21564 14700 21616
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 16672 21496 16724 21548
rect 11520 21428 11572 21437
rect 11428 21360 11480 21412
rect 8760 21292 8812 21344
rect 16304 21428 16356 21480
rect 13820 21403 13872 21412
rect 13820 21369 13829 21403
rect 13829 21369 13863 21403
rect 13863 21369 13872 21403
rect 13820 21360 13872 21369
rect 18236 21428 18288 21480
rect 20996 21428 21048 21480
rect 21456 21471 21508 21480
rect 21456 21437 21465 21471
rect 21465 21437 21499 21471
rect 21499 21437 21508 21471
rect 21456 21428 21508 21437
rect 23020 21564 23072 21616
rect 27160 21632 27212 21684
rect 25412 21564 25464 21616
rect 27344 21564 27396 21616
rect 19064 21360 19116 21412
rect 22192 21360 22244 21412
rect 25228 21471 25280 21480
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 24860 21403 24912 21412
rect 24860 21369 24869 21403
rect 24869 21369 24903 21403
rect 24903 21369 24912 21403
rect 24860 21360 24912 21369
rect 26884 21496 26936 21548
rect 25872 21471 25924 21480
rect 25872 21437 25881 21471
rect 25881 21437 25915 21471
rect 25915 21437 25924 21471
rect 25872 21428 25924 21437
rect 26792 21471 26844 21480
rect 26792 21437 26801 21471
rect 26801 21437 26835 21471
rect 26835 21437 26844 21471
rect 26792 21428 26844 21437
rect 28540 21471 28592 21480
rect 28540 21437 28549 21471
rect 28549 21437 28583 21471
rect 28583 21437 28592 21471
rect 28540 21428 28592 21437
rect 29000 21428 29052 21480
rect 29552 21471 29604 21480
rect 29552 21437 29561 21471
rect 29561 21437 29595 21471
rect 29595 21437 29604 21471
rect 29552 21428 29604 21437
rect 30012 21471 30064 21480
rect 30012 21437 30021 21471
rect 30021 21437 30055 21471
rect 30055 21437 30064 21471
rect 30012 21428 30064 21437
rect 27252 21360 27304 21412
rect 28080 21360 28132 21412
rect 14372 21292 14424 21344
rect 14648 21292 14700 21344
rect 15016 21335 15068 21344
rect 15016 21301 15025 21335
rect 15025 21301 15059 21335
rect 15059 21301 15068 21335
rect 15016 21292 15068 21301
rect 15844 21292 15896 21344
rect 18696 21335 18748 21344
rect 18696 21301 18705 21335
rect 18705 21301 18739 21335
rect 18739 21301 18748 21335
rect 18696 21292 18748 21301
rect 22652 21292 22704 21344
rect 22744 21292 22796 21344
rect 24584 21335 24636 21344
rect 24584 21301 24593 21335
rect 24593 21301 24627 21335
rect 24627 21301 24636 21335
rect 24584 21292 24636 21301
rect 24676 21292 24728 21344
rect 25504 21292 25556 21344
rect 26056 21335 26108 21344
rect 26056 21301 26065 21335
rect 26065 21301 26099 21335
rect 26099 21301 26108 21335
rect 26056 21292 26108 21301
rect 26148 21292 26200 21344
rect 28264 21292 28316 21344
rect 29736 21335 29788 21344
rect 29736 21301 29745 21335
rect 29745 21301 29779 21335
rect 29779 21301 29788 21335
rect 29736 21292 29788 21301
rect 8172 21190 8224 21242
rect 8236 21190 8288 21242
rect 8300 21190 8352 21242
rect 8364 21190 8416 21242
rect 8428 21190 8480 21242
rect 15946 21190 15998 21242
rect 16010 21190 16062 21242
rect 16074 21190 16126 21242
rect 16138 21190 16190 21242
rect 16202 21190 16254 21242
rect 23720 21190 23772 21242
rect 23784 21190 23836 21242
rect 23848 21190 23900 21242
rect 23912 21190 23964 21242
rect 23976 21190 24028 21242
rect 31494 21190 31546 21242
rect 31558 21190 31610 21242
rect 31622 21190 31674 21242
rect 31686 21190 31738 21242
rect 31750 21190 31802 21242
rect 11428 21131 11480 21140
rect 11428 21097 11437 21131
rect 11437 21097 11471 21131
rect 11471 21097 11480 21131
rect 11428 21088 11480 21097
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13360 21088 13412 21097
rect 14372 21088 14424 21140
rect 15752 21088 15804 21140
rect 8852 20952 8904 21004
rect 9864 20952 9916 21004
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 11060 20952 11112 21004
rect 11888 20995 11940 21004
rect 11888 20961 11897 20995
rect 11897 20961 11931 20995
rect 11931 20961 11940 20995
rect 11888 20952 11940 20961
rect 8760 20927 8812 20936
rect 8760 20893 8769 20927
rect 8769 20893 8803 20927
rect 8803 20893 8812 20927
rect 8760 20884 8812 20893
rect 14188 20952 14240 21004
rect 16672 21131 16724 21140
rect 16672 21097 16681 21131
rect 16681 21097 16715 21131
rect 16715 21097 16724 21131
rect 16672 21088 16724 21097
rect 19064 21131 19116 21140
rect 19064 21097 19073 21131
rect 19073 21097 19107 21131
rect 19107 21097 19116 21131
rect 19064 21088 19116 21097
rect 21180 21088 21232 21140
rect 21456 21088 21508 21140
rect 17960 21020 18012 21072
rect 13544 20884 13596 20936
rect 16304 20995 16356 21004
rect 16304 20961 16313 20995
rect 16313 20961 16347 20995
rect 16347 20961 16356 20995
rect 16304 20952 16356 20961
rect 16856 20952 16908 21004
rect 18328 20952 18380 21004
rect 20444 21020 20496 21072
rect 22192 21131 22244 21140
rect 22192 21097 22201 21131
rect 22201 21097 22235 21131
rect 22235 21097 22244 21131
rect 22192 21088 22244 21097
rect 24584 21088 24636 21140
rect 24860 21088 24912 21140
rect 25228 21088 25280 21140
rect 25504 21088 25556 21140
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 18236 20884 18288 20936
rect 19248 20952 19300 21004
rect 20352 20884 20404 20936
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 10876 20748 10928 20800
rect 12808 20791 12860 20800
rect 12808 20757 12817 20791
rect 12817 20757 12851 20791
rect 12851 20757 12860 20791
rect 12808 20748 12860 20757
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 14556 20748 14608 20800
rect 16580 20748 16632 20800
rect 16948 20748 17000 20800
rect 23020 20995 23072 21004
rect 23020 20961 23029 20995
rect 23029 20961 23063 20995
rect 23063 20961 23072 20995
rect 23020 20952 23072 20961
rect 24676 20859 24728 20868
rect 18144 20791 18196 20800
rect 18144 20757 18153 20791
rect 18153 20757 18187 20791
rect 18187 20757 18196 20791
rect 18144 20748 18196 20757
rect 20536 20748 20588 20800
rect 21456 20748 21508 20800
rect 24676 20825 24685 20859
rect 24685 20825 24719 20859
rect 24719 20825 24728 20859
rect 24676 20816 24728 20825
rect 24400 20791 24452 20800
rect 24400 20757 24409 20791
rect 24409 20757 24443 20791
rect 24443 20757 24452 20791
rect 24400 20748 24452 20757
rect 25412 20952 25464 21004
rect 29368 21088 29420 21140
rect 29736 21088 29788 21140
rect 25504 20816 25556 20868
rect 27068 20995 27120 21004
rect 27068 20961 27077 20995
rect 27077 20961 27111 20995
rect 27111 20961 27120 20995
rect 27068 20952 27120 20961
rect 27252 20995 27304 21004
rect 27252 20961 27261 20995
rect 27261 20961 27295 20995
rect 27295 20961 27304 20995
rect 27252 20952 27304 20961
rect 27528 20995 27580 21004
rect 27528 20961 27537 20995
rect 27537 20961 27571 20995
rect 27571 20961 27580 20995
rect 27528 20952 27580 20961
rect 27988 20952 28040 21004
rect 28080 20952 28132 21004
rect 26424 20859 26476 20868
rect 26424 20825 26433 20859
rect 26433 20825 26467 20859
rect 26467 20825 26476 20859
rect 26424 20816 26476 20825
rect 27436 20927 27488 20936
rect 27436 20893 27445 20927
rect 27445 20893 27479 20927
rect 27479 20893 27488 20927
rect 27436 20884 27488 20893
rect 29276 20927 29328 20936
rect 29276 20893 29285 20927
rect 29285 20893 29319 20927
rect 29319 20893 29328 20927
rect 29276 20884 29328 20893
rect 25964 20791 26016 20800
rect 25964 20757 25973 20791
rect 25973 20757 26007 20791
rect 26007 20757 26016 20791
rect 25964 20748 26016 20757
rect 26608 20816 26660 20868
rect 30012 20952 30064 21004
rect 27252 20748 27304 20800
rect 4285 20646 4337 20698
rect 4349 20646 4401 20698
rect 4413 20646 4465 20698
rect 4477 20646 4529 20698
rect 4541 20646 4593 20698
rect 12059 20646 12111 20698
rect 12123 20646 12175 20698
rect 12187 20646 12239 20698
rect 12251 20646 12303 20698
rect 12315 20646 12367 20698
rect 19833 20646 19885 20698
rect 19897 20646 19949 20698
rect 19961 20646 20013 20698
rect 20025 20646 20077 20698
rect 20089 20646 20141 20698
rect 27607 20646 27659 20698
rect 27671 20646 27723 20698
rect 27735 20646 27787 20698
rect 27799 20646 27851 20698
rect 27863 20646 27915 20698
rect 8852 20587 8904 20596
rect 8852 20553 8861 20587
rect 8861 20553 8895 20587
rect 8895 20553 8904 20587
rect 8852 20544 8904 20553
rect 5080 20340 5132 20392
rect 8760 20408 8812 20460
rect 11520 20544 11572 20596
rect 12808 20587 12860 20596
rect 12808 20553 12817 20587
rect 12817 20553 12851 20587
rect 12851 20553 12860 20587
rect 12808 20544 12860 20553
rect 13544 20519 13596 20528
rect 13544 20485 13553 20519
rect 13553 20485 13587 20519
rect 13587 20485 13596 20519
rect 13544 20476 13596 20485
rect 15476 20544 15528 20596
rect 13912 20476 13964 20528
rect 8852 20340 8904 20392
rect 9404 20340 9456 20392
rect 9864 20383 9916 20392
rect 9864 20349 9873 20383
rect 9873 20349 9907 20383
rect 9907 20349 9916 20383
rect 9864 20340 9916 20349
rect 10232 20383 10284 20392
rect 10232 20349 10266 20383
rect 10266 20349 10284 20383
rect 10232 20340 10284 20349
rect 11428 20383 11480 20392
rect 11428 20349 11437 20383
rect 11437 20349 11471 20383
rect 11471 20349 11480 20383
rect 11428 20340 11480 20349
rect 11704 20383 11756 20392
rect 11704 20349 11713 20383
rect 11713 20349 11747 20383
rect 11747 20349 11756 20383
rect 11704 20340 11756 20349
rect 13636 20340 13688 20392
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 14096 20408 14148 20417
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 15752 20408 15804 20460
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 6460 20272 6512 20324
rect 7196 20272 7248 20324
rect 15016 20340 15068 20392
rect 15108 20383 15160 20392
rect 15108 20349 15117 20383
rect 15117 20349 15151 20383
rect 15151 20349 15160 20383
rect 15108 20340 15160 20349
rect 15292 20383 15344 20392
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 16580 20340 16632 20392
rect 17316 20340 17368 20392
rect 17960 20544 18012 20596
rect 18972 20544 19024 20596
rect 20628 20544 20680 20596
rect 20812 20544 20864 20596
rect 27528 20544 27580 20596
rect 17960 20408 18012 20460
rect 18052 20383 18104 20392
rect 18052 20349 18092 20383
rect 18092 20349 18104 20383
rect 18052 20340 18104 20349
rect 19064 20383 19116 20392
rect 19064 20349 19068 20383
rect 19068 20349 19102 20383
rect 19102 20349 19116 20383
rect 19064 20340 19116 20349
rect 19340 20383 19392 20392
rect 19340 20349 19385 20383
rect 19385 20349 19392 20383
rect 19340 20340 19392 20349
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 5172 20204 5224 20256
rect 5448 20204 5500 20256
rect 6184 20247 6236 20256
rect 6184 20213 6193 20247
rect 6193 20213 6227 20247
rect 6227 20213 6236 20247
rect 6184 20204 6236 20213
rect 9036 20247 9088 20256
rect 9036 20213 9045 20247
rect 9045 20213 9079 20247
rect 9079 20213 9088 20247
rect 9036 20204 9088 20213
rect 9772 20247 9824 20256
rect 9772 20213 9781 20247
rect 9781 20213 9815 20247
rect 9815 20213 9824 20247
rect 9772 20204 9824 20213
rect 11612 20247 11664 20256
rect 11612 20213 11621 20247
rect 11621 20213 11655 20247
rect 11655 20213 11664 20247
rect 11612 20204 11664 20213
rect 13452 20204 13504 20256
rect 18972 20272 19024 20324
rect 20168 20340 20220 20392
rect 21456 20408 21508 20460
rect 24492 20519 24544 20528
rect 24492 20485 24501 20519
rect 24501 20485 24535 20519
rect 24535 20485 24544 20519
rect 24492 20476 24544 20485
rect 24676 20476 24728 20528
rect 30012 20544 30064 20596
rect 20536 20383 20588 20392
rect 20536 20349 20539 20383
rect 20539 20349 20573 20383
rect 20573 20349 20588 20383
rect 20536 20340 20588 20349
rect 20720 20383 20772 20392
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 21088 20340 21140 20392
rect 21824 20340 21876 20392
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 22468 20340 22520 20392
rect 22744 20383 22796 20392
rect 22744 20349 22753 20383
rect 22753 20349 22787 20383
rect 22787 20349 22796 20383
rect 22744 20340 22796 20349
rect 22928 20383 22980 20392
rect 22928 20349 22973 20383
rect 22973 20349 22980 20383
rect 22928 20340 22980 20349
rect 23112 20383 23164 20392
rect 23112 20349 23121 20383
rect 23121 20349 23155 20383
rect 23155 20349 23164 20383
rect 23112 20340 23164 20349
rect 24860 20340 24912 20392
rect 18696 20204 18748 20256
rect 22836 20315 22888 20324
rect 22836 20281 22845 20315
rect 22845 20281 22879 20315
rect 22879 20281 22888 20315
rect 22836 20272 22888 20281
rect 23388 20272 23440 20324
rect 24584 20272 24636 20324
rect 19984 20204 20036 20256
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 20260 20204 20312 20256
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 20628 20204 20680 20256
rect 24768 20204 24820 20256
rect 26424 20383 26476 20392
rect 26424 20349 26458 20383
rect 26458 20349 26476 20383
rect 26424 20340 26476 20349
rect 27436 20408 27488 20460
rect 26884 20383 26936 20392
rect 26884 20349 26893 20383
rect 26893 20349 26927 20383
rect 26927 20349 26936 20383
rect 26884 20340 26936 20349
rect 27252 20272 27304 20324
rect 26240 20247 26292 20256
rect 26240 20213 26249 20247
rect 26249 20213 26283 20247
rect 26283 20213 26292 20247
rect 26240 20204 26292 20213
rect 27160 20247 27212 20256
rect 27160 20213 27169 20247
rect 27169 20213 27203 20247
rect 27203 20213 27212 20247
rect 27160 20204 27212 20213
rect 27620 20383 27672 20392
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 28632 20408 28684 20460
rect 28080 20383 28132 20392
rect 28080 20349 28089 20383
rect 28089 20349 28123 20383
rect 28123 20349 28132 20383
rect 28080 20340 28132 20349
rect 28356 20315 28408 20324
rect 28356 20281 28365 20315
rect 28365 20281 28399 20315
rect 28399 20281 28408 20315
rect 28356 20272 28408 20281
rect 27988 20204 28040 20256
rect 29276 20340 29328 20392
rect 28816 20272 28868 20324
rect 29920 20272 29972 20324
rect 8172 20102 8224 20154
rect 8236 20102 8288 20154
rect 8300 20102 8352 20154
rect 8364 20102 8416 20154
rect 8428 20102 8480 20154
rect 15946 20102 15998 20154
rect 16010 20102 16062 20154
rect 16074 20102 16126 20154
rect 16138 20102 16190 20154
rect 16202 20102 16254 20154
rect 23720 20102 23772 20154
rect 23784 20102 23836 20154
rect 23848 20102 23900 20154
rect 23912 20102 23964 20154
rect 23976 20102 24028 20154
rect 31494 20102 31546 20154
rect 31558 20102 31610 20154
rect 31622 20102 31674 20154
rect 31686 20102 31738 20154
rect 31750 20102 31802 20154
rect 2964 19907 3016 19916
rect 2964 19873 2973 19907
rect 2973 19873 3007 19907
rect 3007 19873 3016 19907
rect 2964 19864 3016 19873
rect 3332 19864 3384 19916
rect 6184 20000 6236 20052
rect 6460 20043 6512 20052
rect 6460 20009 6469 20043
rect 6469 20009 6503 20043
rect 6503 20009 6512 20043
rect 6460 20000 6512 20009
rect 5908 19932 5960 19984
rect 9772 20000 9824 20052
rect 10048 20000 10100 20052
rect 10600 20000 10652 20052
rect 9220 19932 9272 19984
rect 9956 19932 10008 19984
rect 10968 19932 11020 19984
rect 4712 19728 4764 19780
rect 5080 19907 5132 19916
rect 5080 19873 5089 19907
rect 5089 19873 5123 19907
rect 5123 19873 5132 19907
rect 5080 19864 5132 19873
rect 5356 19907 5408 19916
rect 5356 19873 5365 19907
rect 5365 19873 5399 19907
rect 5399 19873 5408 19907
rect 5356 19864 5408 19873
rect 6368 19864 6420 19916
rect 6644 19864 6696 19916
rect 8852 19907 8904 19916
rect 8852 19873 8861 19907
rect 8861 19873 8895 19907
rect 8895 19873 8904 19907
rect 8852 19864 8904 19873
rect 9036 19907 9088 19916
rect 9036 19873 9045 19907
rect 9045 19873 9079 19907
rect 9079 19873 9088 19907
rect 9036 19864 9088 19873
rect 9404 19864 9456 19916
rect 5632 19839 5684 19848
rect 5632 19805 5641 19839
rect 5641 19805 5675 19839
rect 5675 19805 5684 19839
rect 5632 19796 5684 19805
rect 8668 19839 8720 19848
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 5448 19771 5500 19780
rect 5448 19737 5457 19771
rect 5457 19737 5491 19771
rect 5491 19737 5500 19771
rect 5448 19728 5500 19737
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 10416 19864 10468 19916
rect 13544 19975 13596 19984
rect 13544 19941 13553 19975
rect 13553 19941 13587 19975
rect 13587 19941 13596 19975
rect 13544 19932 13596 19941
rect 13176 19907 13228 19916
rect 13176 19873 13185 19907
rect 13185 19873 13219 19907
rect 13219 19873 13228 19907
rect 13176 19864 13228 19873
rect 13268 19907 13320 19916
rect 13268 19873 13278 19907
rect 13278 19873 13312 19907
rect 13312 19873 13320 19907
rect 13268 19864 13320 19873
rect 13452 19907 13504 19916
rect 13452 19873 13461 19907
rect 13461 19873 13495 19907
rect 13495 19873 13504 19907
rect 13452 19864 13504 19873
rect 13728 19864 13780 19916
rect 15108 20000 15160 20052
rect 15476 20000 15528 20052
rect 16672 20000 16724 20052
rect 16856 20043 16908 20052
rect 16856 20009 16865 20043
rect 16865 20009 16899 20043
rect 16899 20009 16908 20043
rect 16856 20000 16908 20009
rect 17500 20000 17552 20052
rect 18236 20000 18288 20052
rect 19340 20000 19392 20052
rect 20444 20000 20496 20052
rect 22928 20000 22980 20052
rect 24400 20000 24452 20052
rect 16948 19975 17000 19984
rect 16948 19941 16957 19975
rect 16957 19941 16991 19975
rect 16991 19941 17000 19975
rect 16948 19932 17000 19941
rect 15108 19864 15160 19916
rect 16488 19907 16540 19916
rect 16488 19873 16497 19907
rect 16497 19873 16531 19907
rect 16531 19873 16540 19907
rect 16488 19864 16540 19873
rect 17684 19932 17736 19984
rect 3700 19660 3752 19712
rect 4160 19660 4212 19712
rect 4620 19660 4672 19712
rect 5264 19703 5316 19712
rect 5264 19669 5273 19703
rect 5273 19669 5307 19703
rect 5307 19669 5316 19703
rect 5264 19660 5316 19669
rect 6092 19703 6144 19712
rect 6092 19669 6101 19703
rect 6101 19669 6135 19703
rect 6135 19669 6144 19703
rect 6092 19660 6144 19669
rect 8576 19703 8628 19712
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 9680 19728 9732 19780
rect 9772 19771 9824 19780
rect 9772 19737 9781 19771
rect 9781 19737 9815 19771
rect 9815 19737 9824 19771
rect 9772 19728 9824 19737
rect 9864 19728 9916 19780
rect 10784 19660 10836 19712
rect 14004 19839 14056 19848
rect 14004 19805 14013 19839
rect 14013 19805 14047 19839
rect 14047 19805 14056 19839
rect 14004 19796 14056 19805
rect 14280 19796 14332 19848
rect 19156 19864 19208 19916
rect 19248 19864 19300 19916
rect 13176 19728 13228 19780
rect 13820 19728 13872 19780
rect 11520 19660 11572 19712
rect 12716 19703 12768 19712
rect 12716 19669 12725 19703
rect 12725 19669 12759 19703
rect 12759 19669 12768 19703
rect 12716 19660 12768 19669
rect 13728 19660 13780 19712
rect 17500 19796 17552 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 20536 19932 20588 19984
rect 23112 19932 23164 19984
rect 24768 20000 24820 20052
rect 24860 20000 24912 20052
rect 25688 20000 25740 20052
rect 26148 20000 26200 20052
rect 27160 20000 27212 20052
rect 27620 20000 27672 20052
rect 20444 19907 20496 19916
rect 20444 19873 20453 19907
rect 20453 19873 20487 19907
rect 20487 19873 20496 19907
rect 20444 19864 20496 19873
rect 20904 19864 20956 19916
rect 22100 19864 22152 19916
rect 23296 19864 23348 19916
rect 15844 19660 15896 19712
rect 15936 19703 15988 19712
rect 15936 19669 15945 19703
rect 15945 19669 15979 19703
rect 15979 19669 15988 19703
rect 15936 19660 15988 19669
rect 20444 19771 20496 19780
rect 20444 19737 20453 19771
rect 20453 19737 20487 19771
rect 20487 19737 20496 19771
rect 20444 19728 20496 19737
rect 20812 19796 20864 19848
rect 20996 19796 21048 19848
rect 22744 19839 22796 19848
rect 22744 19805 22753 19839
rect 22753 19805 22787 19839
rect 22787 19805 22796 19839
rect 22744 19796 22796 19805
rect 24308 19864 24360 19916
rect 20076 19660 20128 19712
rect 21180 19728 21232 19780
rect 24860 19907 24912 19916
rect 24860 19873 24869 19907
rect 24869 19873 24903 19907
rect 24903 19873 24912 19907
rect 24860 19864 24912 19873
rect 28356 20000 28408 20052
rect 28816 20000 28868 20052
rect 29920 20043 29972 20052
rect 29920 20009 29929 20043
rect 29929 20009 29963 20043
rect 29963 20009 29972 20043
rect 29920 20000 29972 20009
rect 29368 19932 29420 19984
rect 29644 19932 29696 19984
rect 26056 19864 26108 19916
rect 28264 19864 28316 19916
rect 28356 19907 28408 19916
rect 28356 19873 28365 19907
rect 28365 19873 28399 19907
rect 28399 19873 28408 19907
rect 28356 19864 28408 19873
rect 20628 19660 20680 19712
rect 23664 19660 23716 19712
rect 24124 19703 24176 19712
rect 24124 19669 24133 19703
rect 24133 19669 24167 19703
rect 24167 19669 24176 19703
rect 24124 19660 24176 19669
rect 24216 19703 24268 19712
rect 24216 19669 24225 19703
rect 24225 19669 24259 19703
rect 24259 19669 24268 19703
rect 24216 19660 24268 19669
rect 26700 19703 26752 19712
rect 26700 19669 26709 19703
rect 26709 19669 26743 19703
rect 26743 19669 26752 19703
rect 26700 19660 26752 19669
rect 29092 19864 29144 19916
rect 29368 19728 29420 19780
rect 29276 19703 29328 19712
rect 29276 19669 29285 19703
rect 29285 19669 29319 19703
rect 29319 19669 29328 19703
rect 29276 19660 29328 19669
rect 4285 19558 4337 19610
rect 4349 19558 4401 19610
rect 4413 19558 4465 19610
rect 4477 19558 4529 19610
rect 4541 19558 4593 19610
rect 12059 19558 12111 19610
rect 12123 19558 12175 19610
rect 12187 19558 12239 19610
rect 12251 19558 12303 19610
rect 12315 19558 12367 19610
rect 19833 19558 19885 19610
rect 19897 19558 19949 19610
rect 19961 19558 20013 19610
rect 20025 19558 20077 19610
rect 20089 19558 20141 19610
rect 27607 19558 27659 19610
rect 27671 19558 27723 19610
rect 27735 19558 27787 19610
rect 27799 19558 27851 19610
rect 27863 19558 27915 19610
rect 2964 19456 3016 19508
rect 3332 19456 3384 19508
rect 4620 19456 4672 19508
rect 5632 19456 5684 19508
rect 8668 19456 8720 19508
rect 9312 19456 9364 19508
rect 9772 19456 9824 19508
rect 11060 19456 11112 19508
rect 11244 19499 11296 19508
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 11428 19456 11480 19508
rect 12716 19456 12768 19508
rect 14004 19456 14056 19508
rect 3608 19388 3660 19440
rect 5908 19388 5960 19440
rect 3700 19295 3752 19304
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 4160 19252 4212 19304
rect 4804 19252 4856 19304
rect 4988 19252 5040 19304
rect 5172 19295 5224 19304
rect 5172 19261 5206 19295
rect 5206 19261 5224 19295
rect 5172 19252 5224 19261
rect 6092 19252 6144 19304
rect 6460 19252 6512 19304
rect 6736 19252 6788 19304
rect 6920 19295 6972 19304
rect 6920 19261 6929 19295
rect 6929 19261 6963 19295
rect 6963 19261 6972 19295
rect 6920 19252 6972 19261
rect 9680 19388 9732 19440
rect 7472 19320 7524 19372
rect 8024 19252 8076 19304
rect 8576 19252 8628 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 8852 19295 8904 19304
rect 8852 19261 8861 19295
rect 8861 19261 8895 19295
rect 8895 19261 8904 19295
rect 8852 19252 8904 19261
rect 5264 19184 5316 19236
rect 9312 19252 9364 19304
rect 9404 19295 9456 19304
rect 9404 19261 9413 19295
rect 9413 19261 9447 19295
rect 9447 19261 9456 19295
rect 9404 19252 9456 19261
rect 9588 19295 9640 19304
rect 9588 19261 9597 19295
rect 9597 19261 9631 19295
rect 9631 19261 9640 19295
rect 9588 19252 9640 19261
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 9772 19295 9824 19304
rect 9772 19261 9781 19295
rect 9781 19261 9815 19295
rect 9815 19261 9824 19295
rect 9772 19252 9824 19261
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 4344 19116 4396 19168
rect 6460 19159 6512 19168
rect 6460 19125 6469 19159
rect 6469 19125 6503 19159
rect 6503 19125 6512 19159
rect 6460 19116 6512 19125
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 7104 19159 7156 19168
rect 7104 19125 7113 19159
rect 7113 19125 7147 19159
rect 7147 19125 7156 19159
rect 7104 19116 7156 19125
rect 9496 19184 9548 19236
rect 8944 19116 8996 19168
rect 9864 19116 9916 19168
rect 10048 19363 10100 19372
rect 10048 19329 10057 19363
rect 10057 19329 10091 19363
rect 10091 19329 10100 19363
rect 10048 19320 10100 19329
rect 11060 19320 11112 19372
rect 13268 19388 13320 19440
rect 16488 19456 16540 19508
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 19248 19456 19300 19508
rect 20076 19456 20128 19508
rect 20168 19456 20220 19508
rect 11520 19252 11572 19304
rect 10876 19227 10928 19236
rect 10876 19193 10885 19227
rect 10885 19193 10919 19227
rect 10919 19193 10928 19227
rect 10876 19184 10928 19193
rect 10968 19227 11020 19236
rect 10968 19193 10977 19227
rect 10977 19193 11011 19227
rect 11011 19193 11020 19227
rect 10968 19184 11020 19193
rect 13820 19184 13872 19236
rect 14740 19184 14792 19236
rect 15752 19320 15804 19372
rect 15936 19320 15988 19372
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 19064 19388 19116 19440
rect 17776 19320 17828 19329
rect 18236 19320 18288 19372
rect 17684 19295 17736 19304
rect 17684 19261 17693 19295
rect 17693 19261 17727 19295
rect 17727 19261 17736 19295
rect 17684 19252 17736 19261
rect 18512 19252 18564 19304
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 13544 19116 13596 19168
rect 15016 19116 15068 19168
rect 17132 19116 17184 19168
rect 17960 19227 18012 19236
rect 17960 19193 17969 19227
rect 17969 19193 18003 19227
rect 18003 19193 18012 19227
rect 17960 19184 18012 19193
rect 18328 19227 18380 19236
rect 18328 19193 18337 19227
rect 18337 19193 18371 19227
rect 18371 19193 18380 19227
rect 18328 19184 18380 19193
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 20168 19295 20220 19304
rect 20168 19261 20177 19295
rect 20177 19261 20211 19295
rect 20211 19261 20220 19295
rect 20168 19252 20220 19261
rect 20260 19252 20312 19304
rect 20904 19499 20956 19508
rect 20904 19465 20913 19499
rect 20913 19465 20947 19499
rect 20947 19465 20956 19499
rect 20904 19456 20956 19465
rect 20996 19456 21048 19508
rect 22100 19499 22152 19508
rect 22100 19465 22109 19499
rect 22109 19465 22143 19499
rect 22143 19465 22152 19499
rect 22100 19456 22152 19465
rect 23664 19499 23716 19508
rect 23664 19465 23673 19499
rect 23673 19465 23707 19499
rect 23707 19465 23716 19499
rect 23664 19456 23716 19465
rect 24676 19499 24728 19508
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 24768 19456 24820 19508
rect 27252 19456 27304 19508
rect 29000 19456 29052 19508
rect 20812 19388 20864 19440
rect 20904 19252 20956 19304
rect 29092 19388 29144 19440
rect 26056 19320 26108 19372
rect 18144 19116 18196 19168
rect 19156 19116 19208 19168
rect 19892 19116 19944 19168
rect 20168 19116 20220 19168
rect 23756 19252 23808 19304
rect 24124 19295 24176 19304
rect 24124 19261 24133 19295
rect 24133 19261 24167 19295
rect 24167 19261 24176 19295
rect 24124 19252 24176 19261
rect 24492 19295 24544 19304
rect 24492 19261 24501 19295
rect 24501 19261 24535 19295
rect 24535 19261 24544 19295
rect 24492 19252 24544 19261
rect 24952 19295 25004 19304
rect 24952 19261 24961 19295
rect 24961 19261 24995 19295
rect 24995 19261 25004 19295
rect 24952 19252 25004 19261
rect 25044 19295 25096 19304
rect 25044 19261 25053 19295
rect 25053 19261 25087 19295
rect 25087 19261 25096 19295
rect 25044 19252 25096 19261
rect 26700 19252 26752 19304
rect 29368 19320 29420 19372
rect 23020 19184 23072 19236
rect 24308 19227 24360 19236
rect 24308 19193 24317 19227
rect 24317 19193 24351 19227
rect 24351 19193 24360 19227
rect 24308 19184 24360 19193
rect 22284 19116 22336 19168
rect 25228 19159 25280 19168
rect 25228 19125 25237 19159
rect 25237 19125 25271 19159
rect 25271 19125 25280 19159
rect 25228 19116 25280 19125
rect 25780 19116 25832 19168
rect 27344 19252 27396 19304
rect 27068 19184 27120 19236
rect 28540 19252 28592 19304
rect 29460 19294 29512 19346
rect 29000 19227 29052 19236
rect 29000 19193 29009 19227
rect 29009 19193 29043 19227
rect 29043 19193 29052 19227
rect 29000 19184 29052 19193
rect 29368 19227 29420 19236
rect 29368 19193 29377 19227
rect 29377 19193 29411 19227
rect 29411 19193 29420 19227
rect 29368 19184 29420 19193
rect 29552 19230 29604 19282
rect 26884 19116 26936 19168
rect 26976 19116 27028 19168
rect 27160 19159 27212 19168
rect 27160 19125 27169 19159
rect 27169 19125 27203 19159
rect 27203 19125 27212 19159
rect 27160 19116 27212 19125
rect 27436 19159 27488 19168
rect 27436 19125 27445 19159
rect 27445 19125 27479 19159
rect 27479 19125 27488 19159
rect 27436 19116 27488 19125
rect 29092 19116 29144 19168
rect 29460 19116 29512 19168
rect 29552 19116 29604 19168
rect 29920 19159 29972 19168
rect 29920 19125 29929 19159
rect 29929 19125 29963 19159
rect 29963 19125 29972 19159
rect 29920 19116 29972 19125
rect 30472 19159 30524 19168
rect 30472 19125 30481 19159
rect 30481 19125 30515 19159
rect 30515 19125 30524 19159
rect 30472 19116 30524 19125
rect 8172 19014 8224 19066
rect 8236 19014 8288 19066
rect 8300 19014 8352 19066
rect 8364 19014 8416 19066
rect 8428 19014 8480 19066
rect 15946 19014 15998 19066
rect 16010 19014 16062 19066
rect 16074 19014 16126 19066
rect 16138 19014 16190 19066
rect 16202 19014 16254 19066
rect 23720 19014 23772 19066
rect 23784 19014 23836 19066
rect 23848 19014 23900 19066
rect 23912 19014 23964 19066
rect 23976 19014 24028 19066
rect 31494 19014 31546 19066
rect 31558 19014 31610 19066
rect 31622 19014 31674 19066
rect 31686 19014 31738 19066
rect 31750 19014 31802 19066
rect 2412 18776 2464 18828
rect 5448 18912 5500 18964
rect 3976 18819 4028 18828
rect 3976 18785 3985 18819
rect 3985 18785 4019 18819
rect 4019 18785 4028 18819
rect 3976 18776 4028 18785
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 5632 18887 5684 18896
rect 5632 18853 5641 18887
rect 5641 18853 5675 18887
rect 5675 18853 5684 18887
rect 5632 18844 5684 18853
rect 7104 18912 7156 18964
rect 9404 18912 9456 18964
rect 9036 18844 9088 18896
rect 10968 18912 11020 18964
rect 13820 18912 13872 18964
rect 14648 18955 14700 18964
rect 14648 18921 14657 18955
rect 14657 18921 14691 18955
rect 14691 18921 14700 18955
rect 14648 18912 14700 18921
rect 17776 18912 17828 18964
rect 17960 18912 18012 18964
rect 18328 18912 18380 18964
rect 4712 18776 4764 18828
rect 5172 18776 5224 18828
rect 5356 18819 5408 18828
rect 4620 18708 4672 18760
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 5080 18708 5132 18760
rect 5356 18785 5365 18819
rect 5365 18785 5399 18819
rect 5399 18785 5408 18819
rect 5356 18776 5408 18785
rect 6000 18819 6052 18828
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 6184 18819 6236 18828
rect 6184 18785 6193 18819
rect 6193 18785 6227 18819
rect 6227 18785 6236 18819
rect 6184 18776 6236 18785
rect 6552 18819 6604 18828
rect 6552 18785 6561 18819
rect 6561 18785 6595 18819
rect 6595 18785 6604 18819
rect 6552 18776 6604 18785
rect 6276 18751 6328 18760
rect 6276 18717 6285 18751
rect 6285 18717 6319 18751
rect 6319 18717 6328 18751
rect 6276 18708 6328 18717
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 9404 18776 9456 18828
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 9864 18798 9916 18850
rect 13360 18844 13412 18896
rect 14556 18844 14608 18896
rect 15200 18844 15252 18896
rect 4068 18572 4120 18624
rect 5264 18640 5316 18692
rect 6736 18683 6788 18692
rect 6736 18649 6745 18683
rect 6745 18649 6779 18683
rect 6779 18649 6788 18683
rect 6736 18640 6788 18649
rect 6828 18640 6880 18692
rect 8484 18683 8536 18692
rect 8484 18649 8493 18683
rect 8493 18649 8527 18683
rect 8527 18649 8536 18683
rect 8484 18640 8536 18649
rect 9220 18683 9272 18692
rect 9220 18649 9229 18683
rect 9229 18649 9263 18683
rect 9263 18649 9272 18683
rect 9220 18640 9272 18649
rect 9956 18708 10008 18760
rect 9496 18640 9548 18692
rect 4712 18572 4764 18624
rect 4896 18572 4948 18624
rect 6368 18572 6420 18624
rect 9036 18572 9088 18624
rect 10324 18819 10376 18828
rect 10324 18785 10333 18819
rect 10333 18785 10367 18819
rect 10367 18785 10376 18819
rect 10324 18776 10376 18785
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 11704 18776 11756 18828
rect 12808 18819 12860 18828
rect 12808 18785 12818 18819
rect 12818 18785 12852 18819
rect 12852 18785 12860 18819
rect 12808 18776 12860 18785
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 13176 18819 13228 18828
rect 13176 18785 13190 18819
rect 13190 18785 13224 18819
rect 13224 18785 13228 18819
rect 13176 18776 13228 18785
rect 13452 18819 13504 18828
rect 13452 18785 13461 18819
rect 13461 18785 13495 18819
rect 13495 18785 13504 18819
rect 13452 18776 13504 18785
rect 13544 18819 13596 18828
rect 13544 18785 13554 18819
rect 13554 18785 13588 18819
rect 13588 18785 13596 18819
rect 13544 18776 13596 18785
rect 12992 18708 13044 18760
rect 11152 18640 11204 18692
rect 13912 18776 13964 18828
rect 14188 18819 14240 18828
rect 14188 18785 14197 18819
rect 14197 18785 14231 18819
rect 14231 18785 14240 18819
rect 14188 18776 14240 18785
rect 14740 18708 14792 18760
rect 18236 18776 18288 18828
rect 20076 18844 20128 18896
rect 23020 18955 23072 18964
rect 23020 18921 23029 18955
rect 23029 18921 23063 18955
rect 23063 18921 23072 18955
rect 23020 18912 23072 18921
rect 23480 18912 23532 18964
rect 24952 18912 25004 18964
rect 26148 18912 26200 18964
rect 26884 18912 26936 18964
rect 24400 18887 24452 18896
rect 24400 18853 24409 18887
rect 24409 18853 24443 18887
rect 24443 18853 24452 18887
rect 24400 18844 24452 18853
rect 25044 18844 25096 18896
rect 18512 18776 18564 18828
rect 18972 18776 19024 18828
rect 19156 18776 19208 18828
rect 19248 18708 19300 18760
rect 19432 18776 19484 18828
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 19892 18776 19944 18828
rect 20996 18776 21048 18828
rect 14648 18640 14700 18692
rect 19524 18640 19576 18692
rect 20812 18683 20864 18692
rect 10048 18572 10100 18624
rect 10324 18572 10376 18624
rect 10876 18572 10928 18624
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 13452 18572 13504 18624
rect 15016 18572 15068 18624
rect 17592 18615 17644 18624
rect 17592 18581 17601 18615
rect 17601 18581 17635 18615
rect 17635 18581 17644 18615
rect 17592 18572 17644 18581
rect 18880 18615 18932 18624
rect 18880 18581 18889 18615
rect 18889 18581 18923 18615
rect 18923 18581 18932 18615
rect 18880 18572 18932 18581
rect 19064 18572 19116 18624
rect 19892 18572 19944 18624
rect 20812 18649 20821 18683
rect 20821 18649 20855 18683
rect 20855 18649 20864 18683
rect 20812 18640 20864 18649
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 20996 18572 21048 18624
rect 22652 18708 22704 18760
rect 25872 18819 25924 18828
rect 25872 18785 25881 18819
rect 25881 18785 25915 18819
rect 25915 18785 25924 18819
rect 25872 18776 25924 18785
rect 26056 18776 26108 18828
rect 26976 18844 27028 18896
rect 27436 18912 27488 18964
rect 29000 18912 29052 18964
rect 29368 18912 29420 18964
rect 30472 18912 30524 18964
rect 27436 18776 27488 18828
rect 27988 18776 28040 18828
rect 28724 18819 28776 18828
rect 28724 18785 28733 18819
rect 28733 18785 28767 18819
rect 28767 18785 28776 18819
rect 28724 18776 28776 18785
rect 28908 18819 28960 18828
rect 28908 18785 28917 18819
rect 28917 18785 28951 18819
rect 28951 18785 28960 18819
rect 28908 18776 28960 18785
rect 29000 18819 29052 18828
rect 29000 18785 29009 18819
rect 29009 18785 29043 18819
rect 29043 18785 29052 18819
rect 29000 18776 29052 18785
rect 29184 18819 29236 18828
rect 29184 18785 29193 18819
rect 29193 18785 29227 18819
rect 29227 18785 29236 18819
rect 29184 18776 29236 18785
rect 29460 18776 29512 18828
rect 23572 18708 23624 18760
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 22560 18640 22612 18692
rect 23020 18640 23072 18692
rect 23204 18640 23256 18692
rect 23848 18640 23900 18692
rect 25044 18640 25096 18692
rect 26056 18640 26108 18692
rect 27436 18640 27488 18692
rect 28356 18640 28408 18692
rect 28816 18640 28868 18692
rect 29000 18640 29052 18692
rect 24492 18572 24544 18624
rect 25412 18572 25464 18624
rect 25780 18572 25832 18624
rect 25872 18572 25924 18624
rect 27252 18615 27304 18624
rect 27252 18581 27261 18615
rect 27261 18581 27295 18615
rect 27295 18581 27304 18615
rect 27252 18572 27304 18581
rect 29552 18615 29604 18624
rect 29552 18581 29561 18615
rect 29561 18581 29595 18615
rect 29595 18581 29604 18615
rect 29552 18572 29604 18581
rect 4285 18470 4337 18522
rect 4349 18470 4401 18522
rect 4413 18470 4465 18522
rect 4477 18470 4529 18522
rect 4541 18470 4593 18522
rect 12059 18470 12111 18522
rect 12123 18470 12175 18522
rect 12187 18470 12239 18522
rect 12251 18470 12303 18522
rect 12315 18470 12367 18522
rect 19833 18470 19885 18522
rect 19897 18470 19949 18522
rect 19961 18470 20013 18522
rect 20025 18470 20077 18522
rect 20089 18470 20141 18522
rect 27607 18470 27659 18522
rect 27671 18470 27723 18522
rect 27735 18470 27787 18522
rect 27799 18470 27851 18522
rect 27863 18470 27915 18522
rect 4252 18368 4304 18420
rect 4436 18275 4488 18284
rect 4436 18241 4445 18275
rect 4445 18241 4479 18275
rect 4479 18241 4488 18275
rect 4436 18232 4488 18241
rect 9312 18368 9364 18420
rect 9404 18368 9456 18420
rect 9772 18368 9824 18420
rect 10232 18411 10284 18420
rect 4068 18164 4120 18216
rect 4344 18207 4396 18216
rect 4344 18173 4353 18207
rect 4353 18173 4387 18207
rect 4387 18173 4396 18207
rect 4344 18164 4396 18173
rect 4896 18164 4948 18216
rect 5908 18232 5960 18284
rect 6092 18232 6144 18284
rect 6920 18232 6972 18284
rect 5448 18207 5500 18216
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 6460 18207 6512 18216
rect 6460 18173 6469 18207
rect 6469 18173 6503 18207
rect 6503 18173 6512 18207
rect 6460 18164 6512 18173
rect 7932 18232 7984 18284
rect 7564 18164 7616 18216
rect 9864 18300 9916 18352
rect 10232 18377 10241 18411
rect 10241 18377 10275 18411
rect 10275 18377 10284 18411
rect 10232 18368 10284 18377
rect 10508 18368 10560 18420
rect 10324 18343 10376 18352
rect 10324 18309 10333 18343
rect 10333 18309 10367 18343
rect 10367 18309 10376 18343
rect 10324 18300 10376 18309
rect 10876 18300 10928 18352
rect 13084 18368 13136 18420
rect 10140 18275 10192 18284
rect 10140 18241 10149 18275
rect 10149 18241 10183 18275
rect 10183 18241 10192 18275
rect 10140 18232 10192 18241
rect 10048 18207 10100 18216
rect 5080 18096 5132 18148
rect 5172 18096 5224 18148
rect 9588 18096 9640 18148
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 4804 18028 4856 18080
rect 5264 18028 5316 18080
rect 6276 18028 6328 18080
rect 7012 18028 7064 18080
rect 7472 18028 7524 18080
rect 7748 18028 7800 18080
rect 8024 18028 8076 18080
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10600 18232 10652 18284
rect 10784 18232 10836 18284
rect 10048 18164 10100 18173
rect 9772 18139 9824 18148
rect 9772 18105 9781 18139
rect 9781 18105 9815 18139
rect 9815 18105 9824 18139
rect 9772 18096 9824 18105
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 12440 18300 12492 18352
rect 16304 18368 16356 18420
rect 17684 18368 17736 18420
rect 16672 18300 16724 18352
rect 18236 18300 18288 18352
rect 14740 18232 14792 18284
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 19248 18368 19300 18420
rect 19708 18368 19760 18420
rect 26884 18368 26936 18420
rect 27252 18368 27304 18420
rect 27436 18368 27488 18420
rect 28724 18411 28776 18420
rect 20260 18343 20312 18352
rect 20260 18309 20269 18343
rect 20269 18309 20303 18343
rect 20303 18309 20312 18343
rect 20260 18300 20312 18309
rect 20812 18300 20864 18352
rect 19340 18232 19392 18284
rect 10968 18096 11020 18148
rect 11520 18096 11572 18148
rect 14556 18096 14608 18148
rect 17316 18096 17368 18148
rect 14924 18071 14976 18080
rect 14924 18037 14933 18071
rect 14933 18037 14967 18071
rect 14967 18037 14976 18071
rect 14924 18028 14976 18037
rect 18696 18139 18748 18148
rect 18696 18105 18705 18139
rect 18705 18105 18739 18139
rect 18739 18105 18748 18139
rect 18696 18096 18748 18105
rect 19248 18164 19300 18216
rect 19708 18164 19760 18216
rect 20260 18164 20312 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 20812 18164 20864 18216
rect 20904 18207 20956 18216
rect 20904 18173 20913 18207
rect 20913 18173 20947 18207
rect 20947 18173 20956 18207
rect 20904 18164 20956 18173
rect 22100 18164 22152 18216
rect 22652 18300 22704 18352
rect 24952 18300 25004 18352
rect 27344 18343 27396 18352
rect 27344 18309 27353 18343
rect 27353 18309 27387 18343
rect 27387 18309 27396 18343
rect 27344 18300 27396 18309
rect 23204 18232 23256 18284
rect 23848 18232 23900 18284
rect 28724 18377 28733 18411
rect 28733 18377 28767 18411
rect 28767 18377 28776 18411
rect 28724 18368 28776 18377
rect 29460 18368 29512 18420
rect 29552 18368 29604 18420
rect 29184 18300 29236 18352
rect 22560 18164 22612 18216
rect 22652 18207 22704 18216
rect 22652 18173 22661 18207
rect 22661 18173 22695 18207
rect 22695 18173 22704 18207
rect 22652 18164 22704 18173
rect 23020 18164 23072 18216
rect 23572 18164 23624 18216
rect 24400 18164 24452 18216
rect 18972 18028 19024 18080
rect 19432 18028 19484 18080
rect 24308 18096 24360 18148
rect 24952 18207 25004 18216
rect 24952 18173 24961 18207
rect 24961 18173 24995 18207
rect 24995 18173 25004 18207
rect 24952 18164 25004 18173
rect 26148 18164 26200 18216
rect 26424 18164 26476 18216
rect 26792 18207 26844 18216
rect 26792 18173 26801 18207
rect 26801 18173 26835 18207
rect 26835 18173 26844 18207
rect 26792 18164 26844 18173
rect 27160 18164 27212 18216
rect 28540 18207 28592 18216
rect 28540 18173 28549 18207
rect 28549 18173 28583 18207
rect 28583 18173 28592 18207
rect 28540 18164 28592 18173
rect 29460 18232 29512 18284
rect 24676 18096 24728 18148
rect 23204 18071 23256 18080
rect 23204 18037 23213 18071
rect 23213 18037 23247 18071
rect 23247 18037 23256 18071
rect 23204 18028 23256 18037
rect 23572 18028 23624 18080
rect 24952 18028 25004 18080
rect 29000 18139 29052 18148
rect 29000 18105 29009 18139
rect 29009 18105 29043 18139
rect 29043 18105 29052 18139
rect 29000 18096 29052 18105
rect 29092 18096 29144 18148
rect 29368 18164 29420 18216
rect 8172 17926 8224 17978
rect 8236 17926 8288 17978
rect 8300 17926 8352 17978
rect 8364 17926 8416 17978
rect 8428 17926 8480 17978
rect 15946 17926 15998 17978
rect 16010 17926 16062 17978
rect 16074 17926 16126 17978
rect 16138 17926 16190 17978
rect 16202 17926 16254 17978
rect 23720 17926 23772 17978
rect 23784 17926 23836 17978
rect 23848 17926 23900 17978
rect 23912 17926 23964 17978
rect 23976 17926 24028 17978
rect 31494 17926 31546 17978
rect 31558 17926 31610 17978
rect 31622 17926 31674 17978
rect 31686 17926 31738 17978
rect 31750 17926 31802 17978
rect 4252 17824 4304 17876
rect 4896 17824 4948 17876
rect 4988 17824 5040 17876
rect 5172 17824 5224 17876
rect 1216 17484 1268 17536
rect 4344 17688 4396 17740
rect 4528 17688 4580 17740
rect 4988 17731 5040 17740
rect 4988 17697 4997 17731
rect 4997 17697 5031 17731
rect 5031 17697 5040 17731
rect 4988 17688 5040 17697
rect 5080 17731 5132 17740
rect 5080 17697 5089 17731
rect 5089 17697 5123 17731
rect 5123 17697 5132 17731
rect 5080 17688 5132 17697
rect 5264 17688 5316 17740
rect 7196 17756 7248 17808
rect 5908 17688 5960 17740
rect 6092 17688 6144 17740
rect 6460 17620 6512 17672
rect 6736 17663 6788 17672
rect 6736 17629 6745 17663
rect 6745 17629 6779 17663
rect 6779 17629 6788 17663
rect 6736 17620 6788 17629
rect 7012 17731 7064 17740
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7380 17731 7432 17740
rect 7012 17688 7064 17697
rect 7380 17697 7389 17731
rect 7389 17697 7423 17731
rect 7423 17697 7432 17731
rect 7380 17688 7432 17697
rect 7748 17799 7800 17808
rect 7748 17765 7782 17799
rect 7782 17765 7800 17799
rect 7748 17756 7800 17765
rect 9772 17824 9824 17876
rect 10140 17824 10192 17876
rect 10692 17824 10744 17876
rect 10232 17756 10284 17808
rect 10416 17756 10468 17808
rect 11060 17824 11112 17876
rect 12808 17824 12860 17876
rect 13360 17824 13412 17876
rect 14924 17824 14976 17876
rect 17040 17824 17092 17876
rect 17500 17824 17552 17876
rect 18604 17824 18656 17876
rect 18696 17824 18748 17876
rect 7196 17620 7248 17672
rect 9404 17731 9456 17740
rect 9404 17697 9413 17731
rect 9413 17697 9447 17731
rect 9447 17697 9456 17731
rect 9404 17688 9456 17697
rect 9588 17688 9640 17740
rect 9956 17688 10008 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 5448 17552 5500 17604
rect 6920 17595 6972 17604
rect 6920 17561 6929 17595
rect 6929 17561 6963 17595
rect 6963 17561 6972 17595
rect 6920 17552 6972 17561
rect 7104 17552 7156 17604
rect 6460 17484 6512 17536
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 6828 17527 6880 17536
rect 6828 17493 6837 17527
rect 6837 17493 6871 17527
rect 6871 17493 6880 17527
rect 6828 17484 6880 17493
rect 11336 17731 11388 17740
rect 10692 17552 10744 17604
rect 7748 17484 7800 17536
rect 9404 17484 9456 17536
rect 9772 17484 9824 17536
rect 9864 17527 9916 17536
rect 9864 17493 9873 17527
rect 9873 17493 9907 17527
rect 9907 17493 9916 17527
rect 9864 17484 9916 17493
rect 10232 17484 10284 17536
rect 10416 17484 10468 17536
rect 11336 17697 11345 17731
rect 11345 17697 11379 17731
rect 11379 17697 11388 17731
rect 11336 17688 11388 17697
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 11704 17688 11756 17740
rect 12440 17620 12492 17672
rect 12900 17620 12952 17672
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 13268 17688 13320 17740
rect 13728 17688 13780 17740
rect 17040 17688 17092 17740
rect 17592 17756 17644 17808
rect 19708 17824 19760 17876
rect 22836 17824 22888 17876
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 14832 17663 14884 17672
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 14832 17620 14884 17629
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 18512 17620 18564 17672
rect 18880 17731 18932 17740
rect 18880 17697 18889 17731
rect 18889 17697 18923 17731
rect 18923 17697 18932 17731
rect 18880 17688 18932 17697
rect 19248 17731 19300 17740
rect 19248 17697 19257 17731
rect 19257 17697 19291 17731
rect 19291 17697 19300 17731
rect 19248 17688 19300 17697
rect 23204 17799 23256 17808
rect 19616 17731 19668 17740
rect 19616 17697 19625 17731
rect 19625 17697 19659 17731
rect 19659 17697 19668 17731
rect 19616 17688 19668 17697
rect 15108 17552 15160 17604
rect 13452 17527 13504 17536
rect 13452 17493 13461 17527
rect 13461 17493 13495 17527
rect 13495 17493 13504 17527
rect 13452 17484 13504 17493
rect 13820 17527 13872 17536
rect 13820 17493 13829 17527
rect 13829 17493 13863 17527
rect 13863 17493 13872 17527
rect 13820 17484 13872 17493
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 15660 17484 15712 17493
rect 19524 17552 19576 17604
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20260 17688 20312 17697
rect 23204 17765 23238 17799
rect 23238 17765 23256 17799
rect 23204 17756 23256 17765
rect 24860 17756 24912 17808
rect 20720 17688 20772 17740
rect 22928 17731 22980 17740
rect 22928 17697 22937 17731
rect 22937 17697 22971 17731
rect 22971 17697 22980 17731
rect 22928 17688 22980 17697
rect 26056 17824 26108 17876
rect 26792 17824 26844 17876
rect 29000 17824 29052 17876
rect 29460 17867 29512 17876
rect 29460 17833 29469 17867
rect 29469 17833 29503 17867
rect 29503 17833 29512 17867
rect 29460 17824 29512 17833
rect 25872 17756 25924 17808
rect 29920 17799 29972 17808
rect 29000 17731 29052 17740
rect 29000 17697 29009 17731
rect 29009 17697 29043 17731
rect 29043 17697 29052 17731
rect 29000 17688 29052 17697
rect 29092 17688 29144 17740
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 18512 17484 18564 17536
rect 20260 17552 20312 17604
rect 20444 17552 20496 17604
rect 24952 17620 25004 17672
rect 26608 17663 26660 17672
rect 26608 17629 26617 17663
rect 26617 17629 26651 17663
rect 26651 17629 26660 17663
rect 26608 17620 26660 17629
rect 27528 17663 27580 17672
rect 27528 17629 27537 17663
rect 27537 17629 27571 17663
rect 27571 17629 27580 17663
rect 27528 17620 27580 17629
rect 28816 17620 28868 17672
rect 29276 17688 29328 17740
rect 29920 17765 29954 17799
rect 29954 17765 29972 17799
rect 29920 17756 29972 17765
rect 29552 17731 29604 17740
rect 29552 17697 29561 17731
rect 29561 17697 29595 17731
rect 29595 17697 29604 17731
rect 29552 17688 29604 17697
rect 24860 17552 24912 17604
rect 27988 17552 28040 17604
rect 29460 17552 29512 17604
rect 21088 17527 21140 17536
rect 21088 17493 21097 17527
rect 21097 17493 21131 17527
rect 21131 17493 21140 17527
rect 21088 17484 21140 17493
rect 22652 17484 22704 17536
rect 23572 17484 23624 17536
rect 24400 17527 24452 17536
rect 24400 17493 24409 17527
rect 24409 17493 24443 17527
rect 24443 17493 24452 17527
rect 24400 17484 24452 17493
rect 26148 17484 26200 17536
rect 26332 17484 26384 17536
rect 28172 17484 28224 17536
rect 31024 17527 31076 17536
rect 31024 17493 31033 17527
rect 31033 17493 31067 17527
rect 31067 17493 31076 17527
rect 31024 17484 31076 17493
rect 4285 17382 4337 17434
rect 4349 17382 4401 17434
rect 4413 17382 4465 17434
rect 4477 17382 4529 17434
rect 4541 17382 4593 17434
rect 12059 17382 12111 17434
rect 12123 17382 12175 17434
rect 12187 17382 12239 17434
rect 12251 17382 12303 17434
rect 12315 17382 12367 17434
rect 19833 17382 19885 17434
rect 19897 17382 19949 17434
rect 19961 17382 20013 17434
rect 20025 17382 20077 17434
rect 20089 17382 20141 17434
rect 27607 17382 27659 17434
rect 27671 17382 27723 17434
rect 27735 17382 27787 17434
rect 27799 17382 27851 17434
rect 27863 17382 27915 17434
rect 6736 17280 6788 17332
rect 9588 17280 9640 17332
rect 9772 17280 9824 17332
rect 10508 17280 10560 17332
rect 10692 17280 10744 17332
rect 13452 17280 13504 17332
rect 13820 17280 13872 17332
rect 14372 17280 14424 17332
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 14832 17280 14884 17332
rect 18144 17323 18196 17332
rect 18144 17289 18153 17323
rect 18153 17289 18187 17323
rect 18187 17289 18196 17323
rect 18144 17280 18196 17289
rect 9956 17212 10008 17264
rect 10416 17212 10468 17264
rect 5080 17187 5132 17196
rect 1216 17119 1268 17128
rect 1216 17085 1225 17119
rect 1225 17085 1259 17119
rect 1259 17085 1268 17119
rect 1216 17076 1268 17085
rect 3332 17076 3384 17128
rect 5080 17153 5089 17187
rect 5089 17153 5123 17187
rect 5123 17153 5132 17187
rect 5080 17144 5132 17153
rect 6644 17144 6696 17196
rect 4988 17076 5040 17128
rect 7012 17119 7064 17128
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 7104 17076 7156 17128
rect 7656 17144 7708 17196
rect 7748 17076 7800 17128
rect 10508 17144 10560 17196
rect 10048 17076 10100 17128
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 13728 17212 13780 17264
rect 1492 17051 1544 17060
rect 1492 17017 1501 17051
rect 1501 17017 1535 17051
rect 1535 17017 1544 17051
rect 1492 17008 1544 17017
rect 2228 17008 2280 17060
rect 1400 16940 1452 16992
rect 7656 17008 7708 17060
rect 7104 16983 7156 16992
rect 7104 16949 7113 16983
rect 7113 16949 7147 16983
rect 7147 16949 7156 16983
rect 7104 16940 7156 16949
rect 10600 17008 10652 17060
rect 10876 17076 10928 17128
rect 11980 17144 12032 17196
rect 13176 17076 13228 17128
rect 16488 17212 16540 17264
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 16580 17187 16632 17196
rect 16580 17153 16589 17187
rect 16589 17153 16623 17187
rect 16623 17153 16632 17187
rect 16580 17144 16632 17153
rect 17316 17187 17368 17196
rect 17316 17153 17325 17187
rect 17325 17153 17359 17187
rect 17359 17153 17368 17187
rect 17316 17144 17368 17153
rect 12532 17008 12584 17060
rect 13636 16940 13688 16992
rect 15660 17076 15712 17128
rect 16396 17076 16448 17128
rect 17132 17076 17184 17128
rect 18236 17212 18288 17264
rect 19524 17280 19576 17332
rect 17684 17144 17736 17196
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 18512 17119 18564 17128
rect 18512 17085 18521 17119
rect 18521 17085 18555 17119
rect 18555 17085 18564 17119
rect 18512 17076 18564 17085
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 19248 17119 19300 17128
rect 19248 17085 19257 17119
rect 19257 17085 19291 17119
rect 19291 17085 19300 17119
rect 19248 17076 19300 17085
rect 19432 17076 19484 17128
rect 16304 16940 16356 16992
rect 17960 16940 18012 16992
rect 18696 16983 18748 16992
rect 18696 16949 18705 16983
rect 18705 16949 18739 16983
rect 18739 16949 18748 16983
rect 18696 16940 18748 16949
rect 18972 17051 19024 17060
rect 18972 17017 18981 17051
rect 18981 17017 19015 17051
rect 19015 17017 19024 17051
rect 18972 17008 19024 17017
rect 23204 17280 23256 17332
rect 24492 17323 24544 17332
rect 24492 17289 24501 17323
rect 24501 17289 24535 17323
rect 24535 17289 24544 17323
rect 24492 17280 24544 17289
rect 26608 17280 26660 17332
rect 29552 17280 29604 17332
rect 20260 17212 20312 17264
rect 24676 17212 24728 17264
rect 26700 17212 26752 17264
rect 20352 17076 20404 17128
rect 20996 17076 21048 17128
rect 21088 17076 21140 17128
rect 22284 17076 22336 17128
rect 22560 17076 22612 17128
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 22100 17008 22152 17060
rect 26332 17119 26384 17128
rect 26332 17085 26341 17119
rect 26341 17085 26375 17119
rect 26375 17085 26384 17119
rect 26332 17076 26384 17085
rect 26424 17076 26476 17128
rect 27804 17144 27856 17196
rect 30380 17144 30432 17196
rect 24768 17008 24820 17060
rect 21640 16983 21692 16992
rect 21640 16949 21649 16983
rect 21649 16949 21683 16983
rect 21683 16949 21692 16983
rect 21640 16940 21692 16949
rect 22468 16940 22520 16992
rect 22928 16940 22980 16992
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 24952 16940 25004 16992
rect 25320 16940 25372 16992
rect 27988 17008 28040 17060
rect 28080 17008 28132 17060
rect 28908 17076 28960 17128
rect 29092 17119 29144 17128
rect 29092 17085 29101 17119
rect 29101 17085 29135 17119
rect 29135 17085 29144 17119
rect 29092 17076 29144 17085
rect 29184 17008 29236 17060
rect 29276 17051 29328 17060
rect 29276 17017 29285 17051
rect 29285 17017 29319 17051
rect 29319 17017 29328 17051
rect 29276 17008 29328 17017
rect 26884 16983 26936 16992
rect 26884 16949 26893 16983
rect 26893 16949 26927 16983
rect 26927 16949 26936 16983
rect 26884 16940 26936 16949
rect 29000 16983 29052 16992
rect 29000 16949 29009 16983
rect 29009 16949 29043 16983
rect 29043 16949 29052 16983
rect 29000 16940 29052 16949
rect 29828 16940 29880 16992
rect 29920 16983 29972 16992
rect 29920 16949 29929 16983
rect 29929 16949 29963 16983
rect 29963 16949 29972 16983
rect 29920 16940 29972 16949
rect 8172 16838 8224 16890
rect 8236 16838 8288 16890
rect 8300 16838 8352 16890
rect 8364 16838 8416 16890
rect 8428 16838 8480 16890
rect 15946 16838 15998 16890
rect 16010 16838 16062 16890
rect 16074 16838 16126 16890
rect 16138 16838 16190 16890
rect 16202 16838 16254 16890
rect 23720 16838 23772 16890
rect 23784 16838 23836 16890
rect 23848 16838 23900 16890
rect 23912 16838 23964 16890
rect 23976 16838 24028 16890
rect 31494 16838 31546 16890
rect 31558 16838 31610 16890
rect 31622 16838 31674 16890
rect 31686 16838 31738 16890
rect 31750 16838 31802 16890
rect 1492 16736 1544 16788
rect 2228 16736 2280 16788
rect 1400 16600 1452 16652
rect 1308 16575 1360 16584
rect 1308 16541 1317 16575
rect 1317 16541 1351 16575
rect 1351 16541 1360 16575
rect 1308 16532 1360 16541
rect 2412 16643 2464 16652
rect 2412 16609 2421 16643
rect 2421 16609 2455 16643
rect 2455 16609 2464 16643
rect 2412 16600 2464 16609
rect 4804 16668 4856 16720
rect 7012 16736 7064 16788
rect 7656 16736 7708 16788
rect 9956 16736 10008 16788
rect 3332 16600 3384 16652
rect 3792 16643 3844 16652
rect 3792 16609 3826 16643
rect 3826 16609 3844 16643
rect 3792 16600 3844 16609
rect 7380 16600 7432 16652
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 10600 16736 10652 16788
rect 10692 16736 10744 16788
rect 13544 16736 13596 16788
rect 14004 16736 14056 16788
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 7840 16575 7892 16584
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 7564 16507 7616 16516
rect 7564 16473 7573 16507
rect 7573 16473 7607 16507
rect 7607 16473 7616 16507
rect 7564 16464 7616 16473
rect 10324 16600 10376 16652
rect 10784 16668 10836 16720
rect 10508 16600 10560 16652
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 12992 16532 13044 16584
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 13636 16668 13688 16720
rect 15108 16600 15160 16652
rect 10784 16464 10836 16516
rect 13176 16464 13228 16516
rect 13820 16532 13872 16584
rect 14280 16532 14332 16584
rect 14740 16532 14792 16584
rect 17684 16736 17736 16788
rect 16764 16668 16816 16720
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 17960 16600 18012 16652
rect 2596 16439 2648 16448
rect 2596 16405 2605 16439
rect 2605 16405 2639 16439
rect 2639 16405 2648 16439
rect 2596 16396 2648 16405
rect 7748 16396 7800 16448
rect 13268 16396 13320 16448
rect 15844 16532 15896 16584
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 17592 16532 17644 16584
rect 18144 16643 18196 16652
rect 18144 16609 18153 16643
rect 18153 16609 18187 16643
rect 18187 16609 18196 16643
rect 18144 16600 18196 16609
rect 18236 16643 18288 16652
rect 18236 16609 18245 16643
rect 18245 16609 18279 16643
rect 18279 16609 18288 16643
rect 18236 16600 18288 16609
rect 18880 16736 18932 16788
rect 18788 16668 18840 16720
rect 19340 16668 19392 16720
rect 19524 16736 19576 16788
rect 20996 16668 21048 16720
rect 22468 16736 22520 16788
rect 22560 16668 22612 16720
rect 22836 16711 22888 16720
rect 21548 16600 21600 16652
rect 21640 16643 21692 16652
rect 21640 16609 21649 16643
rect 21649 16609 21683 16643
rect 21683 16609 21692 16643
rect 21640 16600 21692 16609
rect 16580 16396 16632 16448
rect 18604 16532 18656 16584
rect 20996 16532 21048 16584
rect 22468 16600 22520 16652
rect 22836 16677 22845 16711
rect 22845 16677 22879 16711
rect 22879 16677 22888 16711
rect 22836 16668 22888 16677
rect 23112 16736 23164 16788
rect 23204 16736 23256 16788
rect 24860 16736 24912 16788
rect 22100 16532 22152 16584
rect 23204 16643 23256 16652
rect 23204 16609 23213 16643
rect 23213 16609 23247 16643
rect 23247 16609 23256 16643
rect 23204 16600 23256 16609
rect 23296 16600 23348 16652
rect 23572 16600 23624 16652
rect 26884 16736 26936 16788
rect 27436 16736 27488 16788
rect 24676 16600 24728 16652
rect 24768 16643 24820 16652
rect 24768 16609 24777 16643
rect 24777 16609 24811 16643
rect 24811 16609 24820 16643
rect 24768 16600 24820 16609
rect 25228 16643 25280 16652
rect 25228 16609 25232 16643
rect 25232 16609 25266 16643
rect 25266 16609 25280 16643
rect 25228 16600 25280 16609
rect 25320 16643 25372 16652
rect 25320 16609 25329 16643
rect 25329 16609 25363 16643
rect 25363 16609 25372 16643
rect 25320 16600 25372 16609
rect 25412 16643 25464 16652
rect 25412 16609 25421 16643
rect 25421 16609 25455 16643
rect 25455 16609 25464 16643
rect 25412 16600 25464 16609
rect 25504 16643 25556 16652
rect 25504 16609 25549 16643
rect 25549 16609 25556 16643
rect 25504 16600 25556 16609
rect 25688 16643 25740 16652
rect 25688 16609 25697 16643
rect 25697 16609 25731 16643
rect 25731 16609 25740 16643
rect 25688 16600 25740 16609
rect 28080 16779 28132 16788
rect 28080 16745 28089 16779
rect 28089 16745 28123 16779
rect 28123 16745 28132 16779
rect 28080 16736 28132 16745
rect 29092 16736 29144 16788
rect 29276 16736 29328 16788
rect 29920 16736 29972 16788
rect 31300 16779 31352 16788
rect 31300 16745 31309 16779
rect 31309 16745 31343 16779
rect 31343 16745 31352 16779
rect 31300 16736 31352 16745
rect 27436 16532 27488 16584
rect 27804 16600 27856 16652
rect 28908 16643 28960 16652
rect 25780 16507 25832 16516
rect 18236 16396 18288 16448
rect 25780 16473 25789 16507
rect 25789 16473 25823 16507
rect 25823 16473 25832 16507
rect 25780 16464 25832 16473
rect 27252 16507 27304 16516
rect 27252 16473 27261 16507
rect 27261 16473 27295 16507
rect 27295 16473 27304 16507
rect 27252 16464 27304 16473
rect 28908 16609 28917 16643
rect 28917 16609 28951 16643
rect 28951 16609 28960 16643
rect 28908 16600 28960 16609
rect 20444 16396 20496 16448
rect 22192 16439 22244 16448
rect 22192 16405 22201 16439
rect 22201 16405 22235 16439
rect 22235 16405 22244 16439
rect 22192 16396 22244 16405
rect 22560 16439 22612 16448
rect 22560 16405 22569 16439
rect 22569 16405 22603 16439
rect 22603 16405 22612 16439
rect 22560 16396 22612 16405
rect 23848 16439 23900 16448
rect 23848 16405 23857 16439
rect 23857 16405 23891 16439
rect 23891 16405 23900 16439
rect 23848 16396 23900 16405
rect 24216 16439 24268 16448
rect 24216 16405 24225 16439
rect 24225 16405 24259 16439
rect 24259 16405 24268 16439
rect 24216 16396 24268 16405
rect 29000 16507 29052 16516
rect 29000 16473 29009 16507
rect 29009 16473 29043 16507
rect 29043 16473 29052 16507
rect 29000 16464 29052 16473
rect 29552 16643 29604 16652
rect 29552 16609 29561 16643
rect 29561 16609 29595 16643
rect 29595 16609 29604 16643
rect 29552 16600 29604 16609
rect 29828 16600 29880 16652
rect 4285 16294 4337 16346
rect 4349 16294 4401 16346
rect 4413 16294 4465 16346
rect 4477 16294 4529 16346
rect 4541 16294 4593 16346
rect 12059 16294 12111 16346
rect 12123 16294 12175 16346
rect 12187 16294 12239 16346
rect 12251 16294 12303 16346
rect 12315 16294 12367 16346
rect 19833 16294 19885 16346
rect 19897 16294 19949 16346
rect 19961 16294 20013 16346
rect 20025 16294 20077 16346
rect 20089 16294 20141 16346
rect 27607 16294 27659 16346
rect 27671 16294 27723 16346
rect 27735 16294 27787 16346
rect 27799 16294 27851 16346
rect 27863 16294 27915 16346
rect 7748 16192 7800 16244
rect 7840 16192 7892 16244
rect 9680 16192 9732 16244
rect 1124 16056 1176 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 1216 16031 1268 16040
rect 1216 15997 1225 16031
rect 1225 15997 1259 16031
rect 1259 15997 1268 16031
rect 1216 15988 1268 15997
rect 4988 16031 5040 16040
rect 4988 15997 4997 16031
rect 4997 15997 5031 16031
rect 5031 15997 5040 16031
rect 4988 15988 5040 15997
rect 7104 15988 7156 16040
rect 2596 15920 2648 15972
rect 1308 15852 1360 15904
rect 2412 15852 2464 15904
rect 5080 15920 5132 15972
rect 8116 15988 8168 16040
rect 8668 15988 8720 16040
rect 9036 16031 9088 16040
rect 9036 15997 9070 16031
rect 9070 15997 9088 16031
rect 9036 15988 9088 15997
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 10324 15988 10376 16040
rect 12532 16056 12584 16108
rect 10784 15920 10836 15972
rect 10968 15920 11020 15972
rect 14188 16192 14240 16244
rect 15752 16192 15804 16244
rect 16764 16235 16816 16244
rect 16764 16201 16773 16235
rect 16773 16201 16807 16235
rect 16807 16201 16816 16235
rect 16764 16192 16816 16201
rect 18052 16192 18104 16244
rect 18328 16192 18380 16244
rect 20536 16192 20588 16244
rect 20812 16235 20864 16244
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 14464 16124 14516 16176
rect 14740 16124 14792 16176
rect 22376 16192 22428 16244
rect 22468 16192 22520 16244
rect 22652 16192 22704 16244
rect 13636 15988 13688 16040
rect 13728 15988 13780 16040
rect 14096 16056 14148 16108
rect 12532 15920 12584 15972
rect 13084 15963 13136 15972
rect 13084 15929 13093 15963
rect 13093 15929 13127 15963
rect 13127 15929 13136 15963
rect 13084 15920 13136 15929
rect 13820 15852 13872 15904
rect 14648 16056 14700 16108
rect 15568 16056 15620 16108
rect 14556 15988 14608 16040
rect 15108 15988 15160 16040
rect 14188 15963 14240 15972
rect 14188 15929 14197 15963
rect 14197 15929 14231 15963
rect 14231 15929 14240 15963
rect 14188 15920 14240 15929
rect 15292 15988 15344 16040
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 16304 16031 16356 16040
rect 16304 15997 16313 16031
rect 16313 15997 16347 16031
rect 16347 15997 16356 16031
rect 16304 15988 16356 15997
rect 16396 16031 16448 16040
rect 16396 15997 16405 16031
rect 16405 15997 16439 16031
rect 16439 15997 16448 16031
rect 16396 15988 16448 15997
rect 16580 15988 16632 16040
rect 17040 15988 17092 16040
rect 17500 15988 17552 16040
rect 18236 16056 18288 16108
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 18328 15988 18380 16040
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 20260 16056 20312 16108
rect 21364 16124 21416 16176
rect 21824 16056 21876 16108
rect 15568 15852 15620 15904
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 17592 15852 17644 15904
rect 18328 15895 18380 15904
rect 18328 15861 18337 15895
rect 18337 15861 18371 15895
rect 18371 15861 18380 15895
rect 18328 15852 18380 15861
rect 18420 15852 18472 15904
rect 20444 15963 20496 15972
rect 20444 15929 20453 15963
rect 20453 15929 20487 15963
rect 20487 15929 20496 15963
rect 20444 15920 20496 15929
rect 20904 15963 20956 15972
rect 20904 15929 20913 15963
rect 20913 15929 20947 15963
rect 20947 15929 20956 15963
rect 20904 15920 20956 15929
rect 21456 16031 21508 16040
rect 21456 15997 21465 16031
rect 21465 15997 21499 16031
rect 21499 15997 21508 16031
rect 21456 15988 21508 15997
rect 22468 16031 22520 16040
rect 22468 15997 22472 16031
rect 22472 15997 22506 16031
rect 22506 15997 22520 16031
rect 22468 15988 22520 15997
rect 22836 16031 22888 16040
rect 22836 15997 22844 16031
rect 22844 15997 22878 16031
rect 22878 15997 22888 16031
rect 22836 15988 22888 15997
rect 24400 16192 24452 16244
rect 25504 16235 25556 16244
rect 25504 16201 25513 16235
rect 25513 16201 25547 16235
rect 25547 16201 25556 16235
rect 25504 16192 25556 16201
rect 26332 16192 26384 16244
rect 23848 16124 23900 16176
rect 26700 16167 26752 16176
rect 26700 16133 26709 16167
rect 26709 16133 26743 16167
rect 26743 16133 26752 16167
rect 26700 16124 26752 16133
rect 23020 15988 23072 16040
rect 24032 15988 24084 16040
rect 28632 16124 28684 16176
rect 29000 16056 29052 16108
rect 22008 15920 22060 15972
rect 22284 15920 22336 15972
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 21548 15852 21600 15904
rect 23388 15963 23440 15972
rect 23388 15929 23397 15963
rect 23397 15929 23431 15963
rect 23431 15929 23440 15963
rect 23388 15920 23440 15929
rect 24124 15852 24176 15904
rect 27160 15920 27212 15972
rect 25872 15852 25924 15904
rect 29644 15920 29696 15972
rect 8172 15750 8224 15802
rect 8236 15750 8288 15802
rect 8300 15750 8352 15802
rect 8364 15750 8416 15802
rect 8428 15750 8480 15802
rect 15946 15750 15998 15802
rect 16010 15750 16062 15802
rect 16074 15750 16126 15802
rect 16138 15750 16190 15802
rect 16202 15750 16254 15802
rect 23720 15750 23772 15802
rect 23784 15750 23836 15802
rect 23848 15750 23900 15802
rect 23912 15750 23964 15802
rect 23976 15750 24028 15802
rect 31494 15750 31546 15802
rect 31558 15750 31610 15802
rect 31622 15750 31674 15802
rect 31686 15750 31738 15802
rect 31750 15750 31802 15802
rect 1216 15648 1268 15700
rect 1308 15648 1360 15700
rect 2412 15648 2464 15700
rect 3056 15648 3108 15700
rect 3700 15648 3752 15700
rect 7472 15648 7524 15700
rect 2044 15419 2096 15428
rect 2044 15385 2053 15419
rect 2053 15385 2087 15419
rect 2087 15385 2096 15419
rect 2964 15444 3016 15496
rect 3884 15555 3936 15564
rect 3884 15521 3893 15555
rect 3893 15521 3927 15555
rect 3927 15521 3936 15555
rect 3884 15512 3936 15521
rect 4712 15512 4764 15564
rect 5724 15512 5776 15564
rect 7380 15512 7432 15564
rect 7840 15555 7892 15564
rect 7840 15521 7849 15555
rect 7849 15521 7883 15555
rect 7883 15521 7892 15555
rect 7840 15512 7892 15521
rect 8024 15512 8076 15564
rect 6552 15444 6604 15496
rect 7656 15444 7708 15496
rect 8668 15512 8720 15564
rect 9312 15512 9364 15564
rect 10416 15512 10468 15564
rect 14188 15648 14240 15700
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 14464 15648 14516 15700
rect 15476 15648 15528 15700
rect 18512 15691 18564 15700
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 20904 15648 20956 15700
rect 21456 15648 21508 15700
rect 22284 15648 22336 15700
rect 12624 15512 12676 15564
rect 13636 15580 13688 15632
rect 10232 15444 10284 15496
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 12808 15444 12860 15496
rect 13176 15555 13228 15564
rect 13176 15521 13185 15555
rect 13185 15521 13219 15555
rect 13219 15521 13228 15555
rect 13176 15512 13228 15521
rect 13268 15555 13320 15564
rect 13268 15521 13313 15555
rect 13313 15521 13320 15555
rect 13268 15512 13320 15521
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 2044 15376 2096 15385
rect 1676 15308 1728 15360
rect 3884 15376 3936 15428
rect 5080 15376 5132 15428
rect 3424 15351 3476 15360
rect 3424 15317 3433 15351
rect 3433 15317 3467 15351
rect 3467 15317 3476 15351
rect 3424 15308 3476 15317
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 12440 15308 12492 15360
rect 13176 15376 13228 15428
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 13728 15512 13780 15521
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 13912 15555 13964 15564
rect 13912 15521 13921 15555
rect 13921 15521 13955 15555
rect 13955 15521 13964 15555
rect 13912 15512 13964 15521
rect 14096 15512 14148 15564
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 14004 15444 14056 15496
rect 15016 15512 15068 15564
rect 15200 15376 15252 15428
rect 15476 15512 15528 15564
rect 17776 15555 17828 15564
rect 17776 15521 17785 15555
rect 17785 15521 17819 15555
rect 17819 15521 17828 15555
rect 17776 15512 17828 15521
rect 18144 15555 18196 15564
rect 18144 15521 18153 15555
rect 18153 15521 18187 15555
rect 18187 15521 18196 15555
rect 18144 15512 18196 15521
rect 18972 15512 19024 15564
rect 15752 15444 15804 15496
rect 16304 15444 16356 15496
rect 17040 15444 17092 15496
rect 18788 15444 18840 15496
rect 21364 15555 21416 15564
rect 21364 15521 21373 15555
rect 21373 15521 21407 15555
rect 21407 15521 21416 15555
rect 21364 15512 21416 15521
rect 22100 15580 22152 15632
rect 22376 15580 22428 15632
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 22560 15512 22612 15564
rect 23572 15512 23624 15564
rect 25228 15580 25280 15632
rect 25780 15580 25832 15632
rect 25872 15580 25924 15632
rect 25964 15623 26016 15632
rect 25964 15589 25982 15623
rect 25982 15589 26016 15623
rect 25964 15580 26016 15589
rect 27160 15691 27212 15700
rect 27160 15657 27169 15691
rect 27169 15657 27203 15691
rect 27203 15657 27212 15691
rect 27160 15648 27212 15657
rect 29092 15648 29144 15700
rect 30380 15648 30432 15700
rect 27252 15512 27304 15564
rect 27988 15512 28040 15564
rect 28356 15512 28408 15564
rect 28816 15512 28868 15564
rect 24676 15444 24728 15496
rect 15384 15308 15436 15360
rect 24400 15419 24452 15428
rect 24400 15385 24409 15419
rect 24409 15385 24443 15419
rect 24443 15385 24452 15419
rect 24400 15376 24452 15385
rect 20720 15308 20772 15360
rect 22192 15308 22244 15360
rect 22468 15308 22520 15360
rect 23020 15308 23072 15360
rect 24492 15308 24544 15360
rect 28632 15308 28684 15360
rect 4285 15206 4337 15258
rect 4349 15206 4401 15258
rect 4413 15206 4465 15258
rect 4477 15206 4529 15258
rect 4541 15206 4593 15258
rect 12059 15206 12111 15258
rect 12123 15206 12175 15258
rect 12187 15206 12239 15258
rect 12251 15206 12303 15258
rect 12315 15206 12367 15258
rect 19833 15206 19885 15258
rect 19897 15206 19949 15258
rect 19961 15206 20013 15258
rect 20025 15206 20077 15258
rect 20089 15206 20141 15258
rect 27607 15206 27659 15258
rect 27671 15206 27723 15258
rect 27735 15206 27787 15258
rect 27799 15206 27851 15258
rect 27863 15206 27915 15258
rect 5080 15147 5132 15156
rect 5080 15113 5089 15147
rect 5089 15113 5123 15147
rect 5123 15113 5132 15147
rect 5080 15104 5132 15113
rect 7932 15104 7984 15156
rect 7840 15079 7892 15088
rect 7840 15045 7849 15079
rect 7849 15045 7883 15079
rect 7883 15045 7892 15079
rect 7840 15036 7892 15045
rect 4988 14968 5040 15020
rect 5448 15011 5500 15020
rect 5448 14977 5457 15011
rect 5457 14977 5491 15011
rect 5491 14977 5500 15011
rect 5448 14968 5500 14977
rect 7380 14968 7432 15020
rect 2964 14900 3016 14952
rect 3056 14943 3108 14952
rect 3056 14909 3065 14943
rect 3065 14909 3099 14943
rect 3099 14909 3108 14943
rect 3056 14900 3108 14909
rect 3332 14943 3384 14952
rect 3332 14909 3341 14943
rect 3341 14909 3375 14943
rect 3375 14909 3384 14943
rect 3332 14900 3384 14909
rect 5540 14900 5592 14952
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 7748 14943 7800 14952
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 7748 14900 7800 14909
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 3608 14875 3660 14884
rect 3608 14841 3617 14875
rect 3617 14841 3651 14875
rect 3651 14841 3660 14875
rect 3608 14832 3660 14841
rect 4344 14832 4396 14884
rect 2872 14764 2924 14816
rect 3056 14807 3108 14816
rect 3056 14773 3065 14807
rect 3065 14773 3099 14807
rect 3099 14773 3108 14807
rect 3056 14764 3108 14773
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7472 14807 7524 14816
rect 7472 14773 7481 14807
rect 7481 14773 7515 14807
rect 7515 14773 7524 14807
rect 7472 14764 7524 14773
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 9680 15104 9732 15156
rect 10508 15104 10560 15156
rect 13820 15104 13872 15156
rect 14188 15104 14240 15156
rect 15200 15147 15252 15156
rect 15200 15113 15209 15147
rect 15209 15113 15243 15147
rect 15243 15113 15252 15147
rect 15200 15104 15252 15113
rect 15292 15104 15344 15156
rect 16488 15104 16540 15156
rect 13176 15036 13228 15088
rect 9312 14900 9364 14952
rect 10968 14900 11020 14952
rect 12440 14900 12492 14952
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 13636 14943 13688 14952
rect 13636 14909 13646 14943
rect 13646 14909 13680 14943
rect 13680 14909 13688 14943
rect 13636 14900 13688 14909
rect 14096 14900 14148 14952
rect 14188 14900 14240 14952
rect 9220 14764 9272 14816
rect 10232 14832 10284 14884
rect 9496 14764 9548 14816
rect 13728 14764 13780 14816
rect 13912 14875 13964 14884
rect 13912 14841 13921 14875
rect 13921 14841 13955 14875
rect 13955 14841 13964 14875
rect 13912 14832 13964 14841
rect 14832 14943 14884 14952
rect 14832 14909 14846 14943
rect 14846 14909 14880 14943
rect 14880 14909 14884 14943
rect 14832 14900 14884 14909
rect 14740 14875 14792 14884
rect 14740 14841 14749 14875
rect 14749 14841 14783 14875
rect 14783 14841 14792 14875
rect 14740 14832 14792 14841
rect 15384 14968 15436 15020
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 16304 14900 16356 14952
rect 15200 14764 15252 14816
rect 15660 14832 15712 14884
rect 15936 14832 15988 14884
rect 17776 15104 17828 15156
rect 17040 14943 17092 14952
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 17592 14968 17644 15020
rect 17500 14943 17552 14952
rect 17500 14909 17514 14943
rect 17514 14909 17548 14943
rect 17548 14909 17552 14943
rect 17500 14900 17552 14909
rect 17316 14875 17368 14884
rect 17316 14841 17325 14875
rect 17325 14841 17359 14875
rect 17359 14841 17368 14875
rect 17316 14832 17368 14841
rect 17408 14875 17460 14884
rect 17408 14841 17417 14875
rect 17417 14841 17451 14875
rect 17451 14841 17460 14875
rect 17408 14832 17460 14841
rect 18420 14900 18472 14952
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 18880 14943 18932 14952
rect 18880 14909 18887 14943
rect 18887 14909 18932 14943
rect 18880 14900 18932 14909
rect 20168 14900 20220 14952
rect 20352 15011 20404 15020
rect 20352 14977 20361 15011
rect 20361 14977 20395 15011
rect 20395 14977 20404 15011
rect 20352 14968 20404 14977
rect 22192 14900 22244 14952
rect 22468 14900 22520 14952
rect 25228 15147 25280 15156
rect 25228 15113 25237 15147
rect 25237 15113 25271 15147
rect 25271 15113 25280 15147
rect 25228 15104 25280 15113
rect 27528 15104 27580 15156
rect 22928 14943 22980 14952
rect 22928 14909 22937 14943
rect 22937 14909 22971 14943
rect 22971 14909 22980 14943
rect 22928 14900 22980 14909
rect 19708 14832 19760 14884
rect 20352 14764 20404 14816
rect 22100 14832 22152 14884
rect 21732 14807 21784 14816
rect 21732 14773 21741 14807
rect 21741 14773 21775 14807
rect 21775 14773 21784 14807
rect 21732 14764 21784 14773
rect 22008 14764 22060 14816
rect 23296 14764 23348 14816
rect 28632 15011 28684 15020
rect 28632 14977 28641 15011
rect 28641 14977 28675 15011
rect 28675 14977 28684 15011
rect 28632 14968 28684 14977
rect 24492 14900 24544 14952
rect 25872 14900 25924 14952
rect 23480 14832 23532 14884
rect 26056 14875 26108 14884
rect 26056 14841 26090 14875
rect 26090 14841 26108 14875
rect 26056 14832 26108 14841
rect 28724 14832 28776 14884
rect 8172 14662 8224 14714
rect 8236 14662 8288 14714
rect 8300 14662 8352 14714
rect 8364 14662 8416 14714
rect 8428 14662 8480 14714
rect 15946 14662 15998 14714
rect 16010 14662 16062 14714
rect 16074 14662 16126 14714
rect 16138 14662 16190 14714
rect 16202 14662 16254 14714
rect 23720 14662 23772 14714
rect 23784 14662 23836 14714
rect 23848 14662 23900 14714
rect 23912 14662 23964 14714
rect 23976 14662 24028 14714
rect 31494 14662 31546 14714
rect 31558 14662 31610 14714
rect 31622 14662 31674 14714
rect 31686 14662 31738 14714
rect 31750 14662 31802 14714
rect 3056 14560 3108 14612
rect 1308 14492 1360 14544
rect 3608 14560 3660 14612
rect 4344 14560 4396 14612
rect 4804 14560 4856 14612
rect 7472 14560 7524 14612
rect 7564 14560 7616 14612
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 3240 14288 3292 14340
rect 3424 14424 3476 14476
rect 8668 14492 8720 14544
rect 4160 14356 4212 14408
rect 5448 14424 5500 14476
rect 6092 14467 6144 14476
rect 6092 14433 6126 14467
rect 6126 14433 6144 14467
rect 6092 14424 6144 14433
rect 7656 14424 7708 14476
rect 10232 14560 10284 14612
rect 13544 14560 13596 14612
rect 14188 14560 14240 14612
rect 15108 14560 15160 14612
rect 11336 14492 11388 14544
rect 11520 14492 11572 14544
rect 9404 14424 9456 14476
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 7196 14331 7248 14340
rect 7196 14297 7205 14331
rect 7205 14297 7239 14331
rect 7239 14297 7248 14331
rect 7196 14288 7248 14297
rect 9220 14288 9272 14340
rect 1032 14220 1084 14272
rect 2044 14220 2096 14272
rect 2872 14263 2924 14272
rect 2872 14229 2881 14263
rect 2881 14229 2915 14263
rect 2915 14229 2924 14263
rect 2872 14220 2924 14229
rect 9404 14220 9456 14272
rect 10416 14288 10468 14340
rect 10784 14288 10836 14340
rect 10232 14263 10284 14272
rect 10232 14229 10241 14263
rect 10241 14229 10275 14263
rect 10275 14229 10284 14263
rect 10232 14220 10284 14229
rect 10324 14220 10376 14272
rect 11244 14424 11296 14476
rect 10968 14356 11020 14408
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 12532 14424 12584 14476
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 14372 14492 14424 14544
rect 15844 14492 15896 14544
rect 17408 14560 17460 14612
rect 20720 14560 20772 14612
rect 21732 14560 21784 14612
rect 22008 14560 22060 14612
rect 22284 14560 22336 14612
rect 24124 14560 24176 14612
rect 24860 14560 24912 14612
rect 25964 14560 26016 14612
rect 11520 14356 11572 14408
rect 13728 14467 13780 14476
rect 13728 14433 13737 14467
rect 13737 14433 13771 14467
rect 13771 14433 13780 14467
rect 13728 14424 13780 14433
rect 13820 14424 13872 14476
rect 14004 14467 14056 14476
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 14188 14424 14240 14476
rect 11060 14288 11112 14340
rect 11336 14263 11388 14272
rect 11336 14229 11345 14263
rect 11345 14229 11379 14263
rect 11379 14229 11388 14263
rect 11336 14220 11388 14229
rect 12532 14220 12584 14272
rect 14832 14356 14884 14408
rect 16212 14424 16264 14476
rect 19156 14424 19208 14476
rect 14648 14288 14700 14340
rect 17592 14356 17644 14408
rect 18788 14356 18840 14408
rect 15476 14288 15528 14340
rect 15752 14288 15804 14340
rect 21272 14424 21324 14476
rect 28816 14535 28868 14544
rect 28816 14501 28825 14535
rect 28825 14501 28859 14535
rect 28859 14501 28868 14535
rect 28816 14492 28868 14501
rect 29092 14535 29144 14544
rect 29092 14501 29101 14535
rect 29101 14501 29135 14535
rect 29135 14501 29144 14535
rect 29092 14492 29144 14501
rect 22192 14424 22244 14476
rect 22560 14424 22612 14476
rect 22652 14467 22704 14476
rect 22652 14433 22661 14467
rect 22661 14433 22695 14467
rect 22695 14433 22704 14467
rect 22652 14424 22704 14433
rect 24032 14424 24084 14476
rect 26608 14467 26660 14476
rect 26608 14433 26617 14467
rect 26617 14433 26651 14467
rect 26651 14433 26660 14467
rect 26608 14424 26660 14433
rect 28632 14424 28684 14476
rect 28724 14424 28776 14476
rect 29184 14467 29236 14476
rect 29184 14433 29193 14467
rect 29193 14433 29227 14467
rect 29227 14433 29236 14467
rect 29184 14424 29236 14433
rect 23388 14356 23440 14408
rect 25872 14356 25924 14408
rect 25964 14356 26016 14408
rect 23296 14288 23348 14340
rect 18420 14220 18472 14272
rect 20628 14263 20680 14272
rect 20628 14229 20637 14263
rect 20637 14229 20671 14263
rect 20671 14229 20680 14263
rect 20628 14220 20680 14229
rect 21732 14263 21784 14272
rect 21732 14229 21741 14263
rect 21741 14229 21775 14263
rect 21775 14229 21784 14263
rect 21732 14220 21784 14229
rect 24308 14220 24360 14272
rect 26792 14220 26844 14272
rect 27988 14220 28040 14272
rect 28632 14220 28684 14272
rect 4285 14118 4337 14170
rect 4349 14118 4401 14170
rect 4413 14118 4465 14170
rect 4477 14118 4529 14170
rect 4541 14118 4593 14170
rect 12059 14118 12111 14170
rect 12123 14118 12175 14170
rect 12187 14118 12239 14170
rect 12251 14118 12303 14170
rect 12315 14118 12367 14170
rect 19833 14118 19885 14170
rect 19897 14118 19949 14170
rect 19961 14118 20013 14170
rect 20025 14118 20077 14170
rect 20089 14118 20141 14170
rect 27607 14118 27659 14170
rect 27671 14118 27723 14170
rect 27735 14118 27787 14170
rect 27799 14118 27851 14170
rect 27863 14118 27915 14170
rect 1400 14059 1452 14068
rect 1400 14025 1409 14059
rect 1409 14025 1443 14059
rect 1443 14025 1452 14059
rect 1400 14016 1452 14025
rect 7748 14016 7800 14068
rect 9496 14016 9548 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 10232 14016 10284 14068
rect 10416 14016 10468 14068
rect 1308 13948 1360 14000
rect 3332 13948 3384 14000
rect 4160 13948 4212 14000
rect 1676 13880 1728 13932
rect 1032 13855 1084 13864
rect 1032 13821 1041 13855
rect 1041 13821 1075 13855
rect 1075 13821 1084 13855
rect 1032 13812 1084 13821
rect 5448 13880 5500 13932
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 5172 13812 5224 13864
rect 5264 13812 5316 13864
rect 6460 13812 6512 13864
rect 11060 14016 11112 14068
rect 11336 14016 11388 14068
rect 11612 14016 11664 14068
rect 10692 13948 10744 14000
rect 5908 13787 5960 13796
rect 5908 13753 5942 13787
rect 5942 13753 5960 13787
rect 5908 13744 5960 13753
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 14188 14016 14240 14068
rect 17132 14016 17184 14068
rect 18328 14016 18380 14068
rect 20628 14016 20680 14068
rect 21732 14016 21784 14068
rect 23572 14059 23624 14068
rect 23572 14025 23581 14059
rect 23581 14025 23615 14059
rect 23615 14025 23624 14059
rect 23572 14016 23624 14025
rect 25044 14016 25096 14068
rect 26056 14059 26108 14068
rect 26056 14025 26065 14059
rect 26065 14025 26099 14059
rect 26099 14025 26108 14059
rect 26056 14016 26108 14025
rect 26792 14059 26844 14068
rect 26792 14025 26801 14059
rect 26801 14025 26835 14059
rect 26835 14025 26844 14059
rect 26792 14016 26844 14025
rect 28080 14016 28132 14068
rect 28724 14016 28776 14068
rect 11336 13855 11388 13864
rect 11336 13821 11345 13855
rect 11345 13821 11379 13855
rect 11379 13821 11388 13855
rect 11336 13812 11388 13821
rect 10692 13719 10744 13728
rect 10692 13685 10701 13719
rect 10701 13685 10735 13719
rect 10735 13685 10744 13719
rect 10692 13676 10744 13685
rect 10784 13719 10836 13728
rect 10784 13685 10793 13719
rect 10793 13685 10827 13719
rect 10827 13685 10836 13719
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 17592 13812 17644 13864
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 22100 13880 22152 13932
rect 25228 13880 25280 13932
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 17684 13744 17736 13796
rect 18420 13744 18472 13796
rect 22100 13744 22152 13796
rect 22560 13744 22612 13796
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24032 13812 24084 13821
rect 24308 13855 24360 13864
rect 24308 13821 24317 13855
rect 24317 13821 24351 13855
rect 24351 13821 24360 13855
rect 24308 13812 24360 13821
rect 26240 13812 26292 13864
rect 29000 13948 29052 14000
rect 25596 13744 25648 13796
rect 28816 13744 28868 13796
rect 29460 13787 29512 13796
rect 29460 13753 29469 13787
rect 29469 13753 29503 13787
rect 29503 13753 29512 13787
rect 29460 13744 29512 13753
rect 30196 13744 30248 13796
rect 10784 13676 10836 13685
rect 24400 13676 24452 13728
rect 24952 13676 25004 13728
rect 29092 13676 29144 13728
rect 8172 13574 8224 13626
rect 8236 13574 8288 13626
rect 8300 13574 8352 13626
rect 8364 13574 8416 13626
rect 8428 13574 8480 13626
rect 15946 13574 15998 13626
rect 16010 13574 16062 13626
rect 16074 13574 16126 13626
rect 16138 13574 16190 13626
rect 16202 13574 16254 13626
rect 23720 13574 23772 13626
rect 23784 13574 23836 13626
rect 23848 13574 23900 13626
rect 23912 13574 23964 13626
rect 23976 13574 24028 13626
rect 31494 13574 31546 13626
rect 31558 13574 31610 13626
rect 31622 13574 31674 13626
rect 31686 13574 31738 13626
rect 31750 13574 31802 13626
rect 3240 13472 3292 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 6092 13472 6144 13524
rect 1308 13404 1360 13456
rect 3792 13404 3844 13456
rect 4712 13404 4764 13456
rect 14004 13472 14056 13524
rect 15568 13515 15620 13524
rect 15568 13481 15577 13515
rect 15577 13481 15611 13515
rect 15611 13481 15620 13515
rect 15568 13472 15620 13481
rect 18880 13515 18932 13524
rect 18880 13481 18889 13515
rect 18889 13481 18923 13515
rect 18923 13481 18932 13515
rect 18880 13472 18932 13481
rect 19708 13472 19760 13524
rect 5540 13336 5592 13388
rect 5632 13336 5684 13388
rect 5908 13336 5960 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 3332 13268 3384 13320
rect 6276 13200 6328 13252
rect 10692 13336 10744 13388
rect 6460 13268 6512 13320
rect 2872 13175 2924 13184
rect 2872 13141 2881 13175
rect 2881 13141 2915 13175
rect 2915 13141 2924 13175
rect 2872 13132 2924 13141
rect 5816 13175 5868 13184
rect 5816 13141 5825 13175
rect 5825 13141 5859 13175
rect 5859 13141 5868 13175
rect 5816 13132 5868 13141
rect 14648 13404 14700 13456
rect 17960 13404 18012 13456
rect 19064 13404 19116 13456
rect 11612 13336 11664 13388
rect 12624 13336 12676 13388
rect 13360 13336 13412 13388
rect 15016 13336 15068 13388
rect 17592 13336 17644 13388
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 22100 13268 22152 13320
rect 8300 13132 8352 13184
rect 9312 13132 9364 13184
rect 12440 13200 12492 13252
rect 20352 13200 20404 13252
rect 25136 13472 25188 13524
rect 25228 13472 25280 13524
rect 25596 13515 25648 13524
rect 25596 13481 25605 13515
rect 25605 13481 25639 13515
rect 25639 13481 25648 13515
rect 25596 13472 25648 13481
rect 26608 13472 26660 13524
rect 28816 13515 28868 13524
rect 28816 13481 28825 13515
rect 28825 13481 28859 13515
rect 28859 13481 28868 13515
rect 28816 13472 28868 13481
rect 29000 13472 29052 13524
rect 29460 13515 29512 13524
rect 29460 13481 29469 13515
rect 29469 13481 29503 13515
rect 29503 13481 29512 13515
rect 29460 13472 29512 13481
rect 30196 13472 30248 13524
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 12992 13132 13044 13184
rect 20168 13132 20220 13184
rect 21364 13175 21416 13184
rect 21364 13141 21373 13175
rect 21373 13141 21407 13175
rect 21407 13141 21416 13175
rect 21364 13132 21416 13141
rect 23020 13132 23072 13184
rect 24400 13268 24452 13320
rect 24952 13379 25004 13388
rect 24952 13345 24961 13379
rect 24961 13345 24995 13379
rect 24995 13345 25004 13379
rect 24952 13336 25004 13345
rect 25044 13336 25096 13388
rect 25320 13336 25372 13388
rect 23664 13132 23716 13184
rect 24676 13132 24728 13184
rect 27988 13447 28040 13456
rect 27988 13413 27997 13447
rect 27997 13413 28031 13447
rect 28031 13413 28040 13447
rect 27988 13404 28040 13413
rect 28080 13404 28132 13456
rect 28540 13379 28592 13388
rect 28540 13345 28549 13379
rect 28549 13345 28583 13379
rect 28583 13345 28592 13379
rect 28540 13336 28592 13345
rect 28724 13379 28776 13388
rect 28724 13345 28733 13379
rect 28733 13345 28767 13379
rect 28767 13345 28776 13379
rect 28724 13336 28776 13345
rect 29000 13379 29052 13388
rect 29000 13345 29009 13379
rect 29009 13345 29043 13379
rect 29043 13345 29052 13379
rect 29000 13336 29052 13345
rect 29184 13336 29236 13388
rect 26056 13268 26108 13320
rect 25964 13200 26016 13252
rect 30104 13336 30156 13388
rect 28264 13132 28316 13184
rect 28724 13132 28776 13184
rect 4285 13030 4337 13082
rect 4349 13030 4401 13082
rect 4413 13030 4465 13082
rect 4477 13030 4529 13082
rect 4541 13030 4593 13082
rect 12059 13030 12111 13082
rect 12123 13030 12175 13082
rect 12187 13030 12239 13082
rect 12251 13030 12303 13082
rect 12315 13030 12367 13082
rect 19833 13030 19885 13082
rect 19897 13030 19949 13082
rect 19961 13030 20013 13082
rect 20025 13030 20077 13082
rect 20089 13030 20141 13082
rect 27607 13030 27659 13082
rect 27671 13030 27723 13082
rect 27735 13030 27787 13082
rect 27799 13030 27851 13082
rect 27863 13030 27915 13082
rect 1400 12928 1452 12980
rect 4160 12928 4212 12980
rect 4712 12928 4764 12980
rect 5264 12971 5316 12980
rect 5264 12937 5273 12971
rect 5273 12937 5307 12971
rect 5307 12937 5316 12971
rect 5264 12928 5316 12937
rect 5632 12928 5684 12980
rect 5816 12928 5868 12980
rect 12900 12928 12952 12980
rect 13912 12928 13964 12980
rect 19432 12928 19484 12980
rect 20168 12928 20220 12980
rect 22100 12928 22152 12980
rect 22928 12928 22980 12980
rect 24400 12928 24452 12980
rect 24860 12928 24912 12980
rect 2872 12724 2924 12776
rect 3056 12699 3108 12708
rect 3056 12665 3065 12699
rect 3065 12665 3099 12699
rect 3099 12665 3108 12699
rect 3424 12699 3476 12708
rect 3056 12656 3108 12665
rect 3424 12665 3433 12699
rect 3433 12665 3467 12699
rect 3467 12665 3476 12699
rect 3424 12656 3476 12665
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 4804 12724 4856 12776
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 11980 12860 12032 12912
rect 17684 12903 17736 12912
rect 17684 12869 17693 12903
rect 17693 12869 17727 12903
rect 17727 12869 17736 12903
rect 17684 12860 17736 12869
rect 6460 12792 6512 12844
rect 8300 12792 8352 12844
rect 11336 12724 11388 12776
rect 12716 12724 12768 12776
rect 15844 12767 15896 12776
rect 15844 12733 15853 12767
rect 15853 12733 15887 12767
rect 15887 12733 15896 12767
rect 15844 12724 15896 12733
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 2872 12631 2924 12640
rect 2872 12597 2899 12631
rect 2899 12597 2924 12631
rect 5724 12656 5776 12708
rect 6368 12699 6420 12708
rect 6368 12665 6377 12699
rect 6377 12665 6411 12699
rect 6411 12665 6420 12699
rect 6368 12656 6420 12665
rect 7196 12656 7248 12708
rect 7288 12656 7340 12708
rect 9404 12656 9456 12708
rect 10968 12656 11020 12708
rect 13176 12656 13228 12708
rect 16856 12656 16908 12708
rect 2872 12588 2924 12597
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 6736 12588 6788 12640
rect 11612 12588 11664 12640
rect 18972 12656 19024 12708
rect 21364 12724 21416 12776
rect 20352 12656 20404 12708
rect 17868 12631 17920 12640
rect 17868 12597 17877 12631
rect 17877 12597 17911 12631
rect 17911 12597 17920 12631
rect 17868 12588 17920 12597
rect 17960 12631 18012 12640
rect 17960 12597 17969 12631
rect 17969 12597 18003 12631
rect 18003 12597 18012 12631
rect 17960 12588 18012 12597
rect 18420 12588 18472 12640
rect 23480 12767 23532 12776
rect 23480 12733 23489 12767
rect 23489 12733 23523 12767
rect 23523 12733 23532 12767
rect 23480 12724 23532 12733
rect 23664 12767 23716 12776
rect 23664 12733 23673 12767
rect 23673 12733 23707 12767
rect 23707 12733 23716 12767
rect 26424 12928 26476 12980
rect 29184 12928 29236 12980
rect 27160 12860 27212 12912
rect 23664 12724 23716 12733
rect 25228 12767 25280 12776
rect 25228 12733 25237 12767
rect 25237 12733 25271 12767
rect 25271 12733 25280 12767
rect 25228 12724 25280 12733
rect 25964 12792 26016 12844
rect 26240 12724 26292 12776
rect 28080 12792 28132 12844
rect 28724 12792 28776 12844
rect 28540 12724 28592 12776
rect 28632 12767 28684 12776
rect 28632 12733 28641 12767
rect 28641 12733 28675 12767
rect 28675 12733 28684 12767
rect 28632 12724 28684 12733
rect 30104 12792 30156 12844
rect 22560 12631 22612 12640
rect 22560 12597 22569 12631
rect 22569 12597 22603 12631
rect 22603 12597 22612 12631
rect 22560 12588 22612 12597
rect 22744 12588 22796 12640
rect 22928 12588 22980 12640
rect 24676 12588 24728 12640
rect 24952 12631 25004 12640
rect 24952 12597 24961 12631
rect 24961 12597 24995 12631
rect 24995 12597 25004 12631
rect 24952 12588 25004 12597
rect 25136 12588 25188 12640
rect 26792 12588 26844 12640
rect 26976 12631 27028 12640
rect 26976 12597 26985 12631
rect 26985 12597 27019 12631
rect 27019 12597 27028 12631
rect 26976 12588 27028 12597
rect 8172 12486 8224 12538
rect 8236 12486 8288 12538
rect 8300 12486 8352 12538
rect 8364 12486 8416 12538
rect 8428 12486 8480 12538
rect 15946 12486 15998 12538
rect 16010 12486 16062 12538
rect 16074 12486 16126 12538
rect 16138 12486 16190 12538
rect 16202 12486 16254 12538
rect 23720 12486 23772 12538
rect 23784 12486 23836 12538
rect 23848 12486 23900 12538
rect 23912 12486 23964 12538
rect 23976 12486 24028 12538
rect 31494 12486 31546 12538
rect 31558 12486 31610 12538
rect 31622 12486 31674 12538
rect 31686 12486 31738 12538
rect 31750 12486 31802 12538
rect 3056 12384 3108 12436
rect 3608 12316 3660 12368
rect 4068 12384 4120 12436
rect 5356 12384 5408 12436
rect 4712 12316 4764 12368
rect 6092 12384 6144 12436
rect 3332 12180 3384 12232
rect 13084 12384 13136 12436
rect 14740 12384 14792 12436
rect 16396 12384 16448 12436
rect 16856 12384 16908 12436
rect 17776 12384 17828 12436
rect 18328 12384 18380 12436
rect 20536 12384 20588 12436
rect 22652 12427 22704 12436
rect 22652 12393 22661 12427
rect 22661 12393 22695 12427
rect 22695 12393 22704 12427
rect 22652 12384 22704 12393
rect 26424 12427 26476 12436
rect 26424 12393 26433 12427
rect 26433 12393 26467 12427
rect 26467 12393 26476 12427
rect 26424 12384 26476 12393
rect 7196 12248 7248 12300
rect 7288 12291 7340 12300
rect 7288 12257 7297 12291
rect 7297 12257 7331 12291
rect 7331 12257 7340 12291
rect 7288 12248 7340 12257
rect 8024 12248 8076 12300
rect 12716 12316 12768 12368
rect 6368 12180 6420 12232
rect 6552 12180 6604 12232
rect 10416 12248 10468 12300
rect 13728 12248 13780 12300
rect 14648 12248 14700 12300
rect 15200 12248 15252 12300
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 17224 12248 17276 12300
rect 2780 12112 2832 12164
rect 17316 12112 17368 12164
rect 17868 12248 17920 12300
rect 17960 12291 18012 12300
rect 17960 12257 17969 12291
rect 17969 12257 18003 12291
rect 18003 12257 18012 12291
rect 17960 12248 18012 12257
rect 18328 12291 18380 12300
rect 18328 12257 18337 12291
rect 18337 12257 18371 12291
rect 18371 12257 18380 12291
rect 18328 12248 18380 12257
rect 22560 12316 22612 12368
rect 25596 12316 25648 12368
rect 26884 12316 26936 12368
rect 21548 12291 21600 12300
rect 21548 12257 21582 12291
rect 21582 12257 21600 12291
rect 21548 12248 21600 12257
rect 22008 12248 22060 12300
rect 24308 12291 24360 12300
rect 24308 12257 24317 12291
rect 24317 12257 24351 12291
rect 24351 12257 24360 12291
rect 24308 12248 24360 12257
rect 28816 12384 28868 12436
rect 30012 12316 30064 12368
rect 17592 12180 17644 12232
rect 18052 12180 18104 12232
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 27160 12180 27212 12232
rect 26792 12112 26844 12164
rect 28264 12180 28316 12232
rect 6000 12044 6052 12096
rect 6736 12044 6788 12096
rect 8944 12044 8996 12096
rect 9404 12044 9456 12096
rect 11152 12044 11204 12096
rect 16856 12044 16908 12096
rect 21640 12044 21692 12096
rect 21916 12044 21968 12096
rect 23480 12044 23532 12096
rect 24676 12044 24728 12096
rect 4285 11942 4337 11994
rect 4349 11942 4401 11994
rect 4413 11942 4465 11994
rect 4477 11942 4529 11994
rect 4541 11942 4593 11994
rect 12059 11942 12111 11994
rect 12123 11942 12175 11994
rect 12187 11942 12239 11994
rect 12251 11942 12303 11994
rect 12315 11942 12367 11994
rect 19833 11942 19885 11994
rect 19897 11942 19949 11994
rect 19961 11942 20013 11994
rect 20025 11942 20077 11994
rect 20089 11942 20141 11994
rect 27607 11942 27659 11994
rect 27671 11942 27723 11994
rect 27735 11942 27787 11994
rect 27799 11942 27851 11994
rect 27863 11942 27915 11994
rect 4712 11840 4764 11892
rect 6368 11840 6420 11892
rect 10416 11883 10468 11892
rect 10416 11849 10425 11883
rect 10425 11849 10459 11883
rect 10459 11849 10468 11883
rect 10416 11840 10468 11849
rect 14648 11840 14700 11892
rect 15016 11840 15068 11892
rect 4620 11636 4672 11688
rect 5172 11636 5224 11688
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 7196 11704 7248 11756
rect 5724 11568 5776 11620
rect 7288 11568 7340 11620
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 6736 11543 6788 11552
rect 6736 11509 6763 11543
rect 6763 11509 6788 11543
rect 8024 11704 8076 11756
rect 8668 11772 8720 11824
rect 13636 11772 13688 11824
rect 15200 11772 15252 11824
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 9404 11704 9456 11756
rect 6736 11500 6788 11509
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 7564 11500 7616 11509
rect 10508 11500 10560 11552
rect 13360 11636 13412 11688
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 15476 11704 15528 11756
rect 15016 11636 15068 11688
rect 17776 11840 17828 11892
rect 18696 11840 18748 11892
rect 20628 11840 20680 11892
rect 13728 11611 13780 11620
rect 13728 11577 13737 11611
rect 13737 11577 13771 11611
rect 13771 11577 13780 11611
rect 13728 11568 13780 11577
rect 11060 11500 11112 11552
rect 13176 11500 13228 11552
rect 13452 11500 13504 11552
rect 16396 11636 16448 11688
rect 15844 11568 15896 11620
rect 17040 11611 17092 11620
rect 17040 11577 17049 11611
rect 17049 11577 17083 11611
rect 17083 11577 17092 11611
rect 17040 11568 17092 11577
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 17316 11500 17368 11552
rect 18696 11500 18748 11552
rect 19064 11636 19116 11688
rect 22836 11883 22888 11892
rect 22836 11849 22845 11883
rect 22845 11849 22879 11883
rect 22879 11849 22888 11883
rect 22836 11840 22888 11849
rect 23572 11840 23624 11892
rect 24584 11840 24636 11892
rect 25596 11840 25648 11892
rect 24676 11772 24728 11824
rect 22928 11704 22980 11756
rect 23480 11704 23532 11756
rect 21548 11636 21600 11688
rect 24676 11679 24728 11688
rect 24676 11645 24685 11679
rect 24685 11645 24719 11679
rect 24719 11645 24728 11679
rect 24676 11636 24728 11645
rect 24952 11679 25004 11688
rect 24952 11645 24961 11679
rect 24961 11645 24995 11679
rect 24995 11645 25004 11679
rect 24952 11636 25004 11645
rect 25688 11772 25740 11824
rect 20812 11611 20864 11620
rect 20812 11577 20821 11611
rect 20821 11577 20855 11611
rect 20855 11577 20864 11611
rect 20812 11568 20864 11577
rect 20628 11500 20680 11552
rect 21732 11611 21784 11620
rect 21732 11577 21766 11611
rect 21766 11577 21784 11611
rect 21732 11568 21784 11577
rect 21824 11568 21876 11620
rect 28356 11840 28408 11892
rect 28724 11840 28776 11892
rect 30012 11840 30064 11892
rect 26792 11704 26844 11756
rect 28448 11704 28500 11756
rect 30104 11704 30156 11756
rect 20996 11543 21048 11552
rect 20996 11509 21005 11543
rect 21005 11509 21039 11543
rect 21039 11509 21048 11543
rect 20996 11500 21048 11509
rect 21088 11543 21140 11552
rect 21088 11509 21097 11543
rect 21097 11509 21131 11543
rect 21131 11509 21140 11543
rect 21088 11500 21140 11509
rect 22744 11500 22796 11552
rect 28540 11568 28592 11620
rect 28264 11500 28316 11552
rect 8172 11398 8224 11450
rect 8236 11398 8288 11450
rect 8300 11398 8352 11450
rect 8364 11398 8416 11450
rect 8428 11398 8480 11450
rect 15946 11398 15998 11450
rect 16010 11398 16062 11450
rect 16074 11398 16126 11450
rect 16138 11398 16190 11450
rect 16202 11398 16254 11450
rect 23720 11398 23772 11450
rect 23784 11398 23836 11450
rect 23848 11398 23900 11450
rect 23912 11398 23964 11450
rect 23976 11398 24028 11450
rect 31494 11398 31546 11450
rect 31558 11398 31610 11450
rect 31622 11398 31674 11450
rect 31686 11398 31738 11450
rect 31750 11398 31802 11450
rect 3424 11296 3476 11348
rect 6276 11296 6328 11348
rect 7564 11296 7616 11348
rect 8576 11296 8628 11348
rect 10416 11296 10468 11348
rect 13820 11339 13872 11348
rect 5816 11228 5868 11280
rect 7104 11228 7156 11280
rect 8668 11228 8720 11280
rect 12440 11228 12492 11280
rect 13820 11305 13829 11339
rect 13829 11305 13863 11339
rect 13863 11305 13872 11339
rect 13820 11296 13872 11305
rect 15752 11296 15804 11348
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 3700 11092 3752 11144
rect 5724 11092 5776 11144
rect 6460 11092 6512 11144
rect 6552 11092 6604 11144
rect 8944 11160 8996 11212
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 13636 11271 13688 11280
rect 13636 11237 13645 11271
rect 13645 11237 13679 11271
rect 13679 11237 13688 11271
rect 13636 11228 13688 11237
rect 13728 11228 13780 11280
rect 14832 11228 14884 11280
rect 11060 11092 11112 11144
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 7196 11024 7248 11076
rect 13728 11092 13780 11144
rect 15660 11160 15712 11212
rect 16856 11296 16908 11348
rect 17040 11296 17092 11348
rect 17684 11296 17736 11348
rect 21088 11296 21140 11348
rect 21548 11339 21600 11348
rect 21548 11305 21557 11339
rect 21557 11305 21591 11339
rect 21591 11305 21600 11339
rect 21548 11296 21600 11305
rect 21732 11296 21784 11348
rect 17960 11228 18012 11280
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 20628 11160 20680 11212
rect 21916 11203 21968 11212
rect 21916 11169 21925 11203
rect 21925 11169 21959 11203
rect 21959 11169 21968 11203
rect 21916 11160 21968 11169
rect 22744 11160 22796 11212
rect 21548 11092 21600 11144
rect 23480 11160 23532 11212
rect 22928 11135 22980 11144
rect 22928 11101 22937 11135
rect 22937 11101 22971 11135
rect 22971 11101 22980 11135
rect 22928 11092 22980 11101
rect 24768 11296 24820 11348
rect 28080 11296 28132 11348
rect 28448 11296 28500 11348
rect 28540 11339 28592 11348
rect 28540 11305 28549 11339
rect 28549 11305 28583 11339
rect 28583 11305 28592 11339
rect 28540 11296 28592 11305
rect 24676 11228 24728 11280
rect 27436 11228 27488 11280
rect 25412 11203 25464 11212
rect 25412 11169 25421 11203
rect 25421 11169 25455 11203
rect 25455 11169 25464 11203
rect 25412 11160 25464 11169
rect 28724 11160 28776 11212
rect 7748 10956 7800 11008
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 13176 10956 13228 10965
rect 13452 10999 13504 11008
rect 13452 10965 13461 10999
rect 13461 10965 13495 10999
rect 13495 10965 13504 10999
rect 13452 10956 13504 10965
rect 14004 10956 14056 11008
rect 14096 10956 14148 11008
rect 19432 10956 19484 11008
rect 20812 10956 20864 11008
rect 21732 10956 21784 11008
rect 4285 10854 4337 10906
rect 4349 10854 4401 10906
rect 4413 10854 4465 10906
rect 4477 10854 4529 10906
rect 4541 10854 4593 10906
rect 12059 10854 12111 10906
rect 12123 10854 12175 10906
rect 12187 10854 12239 10906
rect 12251 10854 12303 10906
rect 12315 10854 12367 10906
rect 19833 10854 19885 10906
rect 19897 10854 19949 10906
rect 19961 10854 20013 10906
rect 20025 10854 20077 10906
rect 20089 10854 20141 10906
rect 27607 10854 27659 10906
rect 27671 10854 27723 10906
rect 27735 10854 27787 10906
rect 27799 10854 27851 10906
rect 27863 10854 27915 10906
rect 7104 10752 7156 10804
rect 7472 10752 7524 10804
rect 11428 10752 11480 10804
rect 12440 10752 12492 10804
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 20628 10752 20680 10804
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 25412 10752 25464 10804
rect 27436 10795 27488 10804
rect 27436 10761 27445 10795
rect 27445 10761 27479 10795
rect 27479 10761 27488 10795
rect 27436 10752 27488 10761
rect 6460 10659 6512 10668
rect 6460 10625 6469 10659
rect 6469 10625 6503 10659
rect 6503 10625 6512 10659
rect 6460 10616 6512 10625
rect 7748 10616 7800 10668
rect 8668 10616 8720 10668
rect 11980 10616 12032 10668
rect 5724 10548 5776 10600
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10692 10548 10744 10600
rect 11060 10548 11112 10600
rect 8576 10412 8628 10464
rect 10416 10480 10468 10532
rect 13452 10548 13504 10600
rect 13176 10480 13228 10532
rect 16396 10659 16448 10668
rect 16396 10625 16405 10659
rect 16405 10625 16439 10659
rect 16439 10625 16448 10659
rect 16396 10616 16448 10625
rect 14004 10548 14056 10600
rect 19432 10616 19484 10668
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 24308 10616 24360 10668
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 13820 10523 13872 10532
rect 13820 10489 13829 10523
rect 13829 10489 13863 10523
rect 13863 10489 13872 10523
rect 13820 10480 13872 10489
rect 16672 10523 16724 10532
rect 16672 10489 16681 10523
rect 16681 10489 16715 10523
rect 16715 10489 16724 10523
rect 16672 10480 16724 10489
rect 18696 10480 18748 10532
rect 15200 10412 15252 10464
rect 17684 10412 17736 10464
rect 18052 10412 18104 10464
rect 21548 10548 21600 10600
rect 19800 10480 19852 10532
rect 20352 10412 20404 10464
rect 25688 10548 25740 10600
rect 23020 10480 23072 10532
rect 24216 10523 24268 10532
rect 24216 10489 24225 10523
rect 24225 10489 24259 10523
rect 24259 10489 24268 10523
rect 24216 10480 24268 10489
rect 8172 10310 8224 10362
rect 8236 10310 8288 10362
rect 8300 10310 8352 10362
rect 8364 10310 8416 10362
rect 8428 10310 8480 10362
rect 15946 10310 15998 10362
rect 16010 10310 16062 10362
rect 16074 10310 16126 10362
rect 16138 10310 16190 10362
rect 16202 10310 16254 10362
rect 23720 10310 23772 10362
rect 23784 10310 23836 10362
rect 23848 10310 23900 10362
rect 23912 10310 23964 10362
rect 23976 10310 24028 10362
rect 31494 10310 31546 10362
rect 31558 10310 31610 10362
rect 31622 10310 31674 10362
rect 31686 10310 31738 10362
rect 31750 10310 31802 10362
rect 8576 10208 8628 10260
rect 10416 10208 10468 10260
rect 11152 10208 11204 10260
rect 10508 10072 10560 10124
rect 13728 10208 13780 10260
rect 15292 10208 15344 10260
rect 16672 10208 16724 10260
rect 19800 10251 19852 10260
rect 19800 10217 19809 10251
rect 19809 10217 19843 10251
rect 19843 10217 19852 10251
rect 19800 10208 19852 10217
rect 21180 10208 21232 10260
rect 12532 10140 12584 10192
rect 13452 10140 13504 10192
rect 15200 10072 15252 10124
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 13912 10047 13964 10056
rect 13912 10013 13921 10047
rect 13921 10013 13955 10047
rect 13955 10013 13964 10047
rect 13912 10004 13964 10013
rect 16856 10140 16908 10192
rect 17684 10072 17736 10124
rect 18696 10072 18748 10124
rect 22008 10208 22060 10260
rect 23020 10208 23072 10260
rect 24216 10208 24268 10260
rect 21732 10140 21784 10192
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 22008 10072 22060 10124
rect 21916 10004 21968 10056
rect 25412 9936 25464 9988
rect 21640 9868 21692 9920
rect 4285 9766 4337 9818
rect 4349 9766 4401 9818
rect 4413 9766 4465 9818
rect 4477 9766 4529 9818
rect 4541 9766 4593 9818
rect 12059 9766 12111 9818
rect 12123 9766 12175 9818
rect 12187 9766 12239 9818
rect 12251 9766 12303 9818
rect 12315 9766 12367 9818
rect 19833 9766 19885 9818
rect 19897 9766 19949 9818
rect 19961 9766 20013 9818
rect 20025 9766 20077 9818
rect 20089 9766 20141 9818
rect 27607 9766 27659 9818
rect 27671 9766 27723 9818
rect 27735 9766 27787 9818
rect 27799 9766 27851 9818
rect 27863 9766 27915 9818
rect 11520 9664 11572 9716
rect 13912 9664 13964 9716
rect 12532 9596 12584 9648
rect 11980 9528 12032 9580
rect 13452 9528 13504 9580
rect 13636 9460 13688 9512
rect 8172 9222 8224 9274
rect 8236 9222 8288 9274
rect 8300 9222 8352 9274
rect 8364 9222 8416 9274
rect 8428 9222 8480 9274
rect 15946 9222 15998 9274
rect 16010 9222 16062 9274
rect 16074 9222 16126 9274
rect 16138 9222 16190 9274
rect 16202 9222 16254 9274
rect 23720 9222 23772 9274
rect 23784 9222 23836 9274
rect 23848 9222 23900 9274
rect 23912 9222 23964 9274
rect 23976 9222 24028 9274
rect 31494 9222 31546 9274
rect 31558 9222 31610 9274
rect 31622 9222 31674 9274
rect 31686 9222 31738 9274
rect 31750 9222 31802 9274
rect 4285 8678 4337 8730
rect 4349 8678 4401 8730
rect 4413 8678 4465 8730
rect 4477 8678 4529 8730
rect 4541 8678 4593 8730
rect 12059 8678 12111 8730
rect 12123 8678 12175 8730
rect 12187 8678 12239 8730
rect 12251 8678 12303 8730
rect 12315 8678 12367 8730
rect 19833 8678 19885 8730
rect 19897 8678 19949 8730
rect 19961 8678 20013 8730
rect 20025 8678 20077 8730
rect 20089 8678 20141 8730
rect 27607 8678 27659 8730
rect 27671 8678 27723 8730
rect 27735 8678 27787 8730
rect 27799 8678 27851 8730
rect 27863 8678 27915 8730
rect 8172 8134 8224 8186
rect 8236 8134 8288 8186
rect 8300 8134 8352 8186
rect 8364 8134 8416 8186
rect 8428 8134 8480 8186
rect 15946 8134 15998 8186
rect 16010 8134 16062 8186
rect 16074 8134 16126 8186
rect 16138 8134 16190 8186
rect 16202 8134 16254 8186
rect 23720 8134 23772 8186
rect 23784 8134 23836 8186
rect 23848 8134 23900 8186
rect 23912 8134 23964 8186
rect 23976 8134 24028 8186
rect 31494 8134 31546 8186
rect 31558 8134 31610 8186
rect 31622 8134 31674 8186
rect 31686 8134 31738 8186
rect 31750 8134 31802 8186
rect 4285 7590 4337 7642
rect 4349 7590 4401 7642
rect 4413 7590 4465 7642
rect 4477 7590 4529 7642
rect 4541 7590 4593 7642
rect 12059 7590 12111 7642
rect 12123 7590 12175 7642
rect 12187 7590 12239 7642
rect 12251 7590 12303 7642
rect 12315 7590 12367 7642
rect 19833 7590 19885 7642
rect 19897 7590 19949 7642
rect 19961 7590 20013 7642
rect 20025 7590 20077 7642
rect 20089 7590 20141 7642
rect 27607 7590 27659 7642
rect 27671 7590 27723 7642
rect 27735 7590 27787 7642
rect 27799 7590 27851 7642
rect 27863 7590 27915 7642
rect 8172 7046 8224 7098
rect 8236 7046 8288 7098
rect 8300 7046 8352 7098
rect 8364 7046 8416 7098
rect 8428 7046 8480 7098
rect 15946 7046 15998 7098
rect 16010 7046 16062 7098
rect 16074 7046 16126 7098
rect 16138 7046 16190 7098
rect 16202 7046 16254 7098
rect 23720 7046 23772 7098
rect 23784 7046 23836 7098
rect 23848 7046 23900 7098
rect 23912 7046 23964 7098
rect 23976 7046 24028 7098
rect 31494 7046 31546 7098
rect 31558 7046 31610 7098
rect 31622 7046 31674 7098
rect 31686 7046 31738 7098
rect 31750 7046 31802 7098
rect 4285 6502 4337 6554
rect 4349 6502 4401 6554
rect 4413 6502 4465 6554
rect 4477 6502 4529 6554
rect 4541 6502 4593 6554
rect 12059 6502 12111 6554
rect 12123 6502 12175 6554
rect 12187 6502 12239 6554
rect 12251 6502 12303 6554
rect 12315 6502 12367 6554
rect 19833 6502 19885 6554
rect 19897 6502 19949 6554
rect 19961 6502 20013 6554
rect 20025 6502 20077 6554
rect 20089 6502 20141 6554
rect 27607 6502 27659 6554
rect 27671 6502 27723 6554
rect 27735 6502 27787 6554
rect 27799 6502 27851 6554
rect 27863 6502 27915 6554
rect 8172 5958 8224 6010
rect 8236 5958 8288 6010
rect 8300 5958 8352 6010
rect 8364 5958 8416 6010
rect 8428 5958 8480 6010
rect 15946 5958 15998 6010
rect 16010 5958 16062 6010
rect 16074 5958 16126 6010
rect 16138 5958 16190 6010
rect 16202 5958 16254 6010
rect 23720 5958 23772 6010
rect 23784 5958 23836 6010
rect 23848 5958 23900 6010
rect 23912 5958 23964 6010
rect 23976 5958 24028 6010
rect 31494 5958 31546 6010
rect 31558 5958 31610 6010
rect 31622 5958 31674 6010
rect 31686 5958 31738 6010
rect 31750 5958 31802 6010
rect 4285 5414 4337 5466
rect 4349 5414 4401 5466
rect 4413 5414 4465 5466
rect 4477 5414 4529 5466
rect 4541 5414 4593 5466
rect 12059 5414 12111 5466
rect 12123 5414 12175 5466
rect 12187 5414 12239 5466
rect 12251 5414 12303 5466
rect 12315 5414 12367 5466
rect 19833 5414 19885 5466
rect 19897 5414 19949 5466
rect 19961 5414 20013 5466
rect 20025 5414 20077 5466
rect 20089 5414 20141 5466
rect 27607 5414 27659 5466
rect 27671 5414 27723 5466
rect 27735 5414 27787 5466
rect 27799 5414 27851 5466
rect 27863 5414 27915 5466
rect 8172 4870 8224 4922
rect 8236 4870 8288 4922
rect 8300 4870 8352 4922
rect 8364 4870 8416 4922
rect 8428 4870 8480 4922
rect 15946 4870 15998 4922
rect 16010 4870 16062 4922
rect 16074 4870 16126 4922
rect 16138 4870 16190 4922
rect 16202 4870 16254 4922
rect 23720 4870 23772 4922
rect 23784 4870 23836 4922
rect 23848 4870 23900 4922
rect 23912 4870 23964 4922
rect 23976 4870 24028 4922
rect 31494 4870 31546 4922
rect 31558 4870 31610 4922
rect 31622 4870 31674 4922
rect 31686 4870 31738 4922
rect 31750 4870 31802 4922
rect 4285 4326 4337 4378
rect 4349 4326 4401 4378
rect 4413 4326 4465 4378
rect 4477 4326 4529 4378
rect 4541 4326 4593 4378
rect 12059 4326 12111 4378
rect 12123 4326 12175 4378
rect 12187 4326 12239 4378
rect 12251 4326 12303 4378
rect 12315 4326 12367 4378
rect 19833 4326 19885 4378
rect 19897 4326 19949 4378
rect 19961 4326 20013 4378
rect 20025 4326 20077 4378
rect 20089 4326 20141 4378
rect 27607 4326 27659 4378
rect 27671 4326 27723 4378
rect 27735 4326 27787 4378
rect 27799 4326 27851 4378
rect 27863 4326 27915 4378
rect 8172 3782 8224 3834
rect 8236 3782 8288 3834
rect 8300 3782 8352 3834
rect 8364 3782 8416 3834
rect 8428 3782 8480 3834
rect 15946 3782 15998 3834
rect 16010 3782 16062 3834
rect 16074 3782 16126 3834
rect 16138 3782 16190 3834
rect 16202 3782 16254 3834
rect 23720 3782 23772 3834
rect 23784 3782 23836 3834
rect 23848 3782 23900 3834
rect 23912 3782 23964 3834
rect 23976 3782 24028 3834
rect 31494 3782 31546 3834
rect 31558 3782 31610 3834
rect 31622 3782 31674 3834
rect 31686 3782 31738 3834
rect 31750 3782 31802 3834
rect 4285 3238 4337 3290
rect 4349 3238 4401 3290
rect 4413 3238 4465 3290
rect 4477 3238 4529 3290
rect 4541 3238 4593 3290
rect 12059 3238 12111 3290
rect 12123 3238 12175 3290
rect 12187 3238 12239 3290
rect 12251 3238 12303 3290
rect 12315 3238 12367 3290
rect 19833 3238 19885 3290
rect 19897 3238 19949 3290
rect 19961 3238 20013 3290
rect 20025 3238 20077 3290
rect 20089 3238 20141 3290
rect 27607 3238 27659 3290
rect 27671 3238 27723 3290
rect 27735 3238 27787 3290
rect 27799 3238 27851 3290
rect 27863 3238 27915 3290
rect 8172 2694 8224 2746
rect 8236 2694 8288 2746
rect 8300 2694 8352 2746
rect 8364 2694 8416 2746
rect 8428 2694 8480 2746
rect 15946 2694 15998 2746
rect 16010 2694 16062 2746
rect 16074 2694 16126 2746
rect 16138 2694 16190 2746
rect 16202 2694 16254 2746
rect 23720 2694 23772 2746
rect 23784 2694 23836 2746
rect 23848 2694 23900 2746
rect 23912 2694 23964 2746
rect 23976 2694 24028 2746
rect 31494 2694 31546 2746
rect 31558 2694 31610 2746
rect 31622 2694 31674 2746
rect 31686 2694 31738 2746
rect 31750 2694 31802 2746
rect 4285 2150 4337 2202
rect 4349 2150 4401 2202
rect 4413 2150 4465 2202
rect 4477 2150 4529 2202
rect 4541 2150 4593 2202
rect 12059 2150 12111 2202
rect 12123 2150 12175 2202
rect 12187 2150 12239 2202
rect 12251 2150 12303 2202
rect 12315 2150 12367 2202
rect 19833 2150 19885 2202
rect 19897 2150 19949 2202
rect 19961 2150 20013 2202
rect 20025 2150 20077 2202
rect 20089 2150 20141 2202
rect 27607 2150 27659 2202
rect 27671 2150 27723 2202
rect 27735 2150 27787 2202
rect 27799 2150 27851 2202
rect 27863 2150 27915 2202
rect 8172 1606 8224 1658
rect 8236 1606 8288 1658
rect 8300 1606 8352 1658
rect 8364 1606 8416 1658
rect 8428 1606 8480 1658
rect 15946 1606 15998 1658
rect 16010 1606 16062 1658
rect 16074 1606 16126 1658
rect 16138 1606 16190 1658
rect 16202 1606 16254 1658
rect 23720 1606 23772 1658
rect 23784 1606 23836 1658
rect 23848 1606 23900 1658
rect 23912 1606 23964 1658
rect 23976 1606 24028 1658
rect 31494 1606 31546 1658
rect 31558 1606 31610 1658
rect 31622 1606 31674 1658
rect 31686 1606 31738 1658
rect 31750 1606 31802 1658
rect 4285 1062 4337 1114
rect 4349 1062 4401 1114
rect 4413 1062 4465 1114
rect 4477 1062 4529 1114
rect 4541 1062 4593 1114
rect 12059 1062 12111 1114
rect 12123 1062 12175 1114
rect 12187 1062 12239 1114
rect 12251 1062 12303 1114
rect 12315 1062 12367 1114
rect 19833 1062 19885 1114
rect 19897 1062 19949 1114
rect 19961 1062 20013 1114
rect 20025 1062 20077 1114
rect 20089 1062 20141 1114
rect 27607 1062 27659 1114
rect 27671 1062 27723 1114
rect 27735 1062 27787 1114
rect 27799 1062 27851 1114
rect 27863 1062 27915 1114
rect 8172 518 8224 570
rect 8236 518 8288 570
rect 8300 518 8352 570
rect 8364 518 8416 570
rect 8428 518 8480 570
rect 15946 518 15998 570
rect 16010 518 16062 570
rect 16074 518 16126 570
rect 16138 518 16190 570
rect 16202 518 16254 570
rect 23720 518 23772 570
rect 23784 518 23836 570
rect 23848 518 23900 570
rect 23912 518 23964 570
rect 23976 518 24028 570
rect 31494 518 31546 570
rect 31558 518 31610 570
rect 31622 518 31674 570
rect 31686 518 31738 570
rect 31750 518 31802 570
<< metal2 >>
rect 4526 21992 4582 22001
rect 8206 21992 8262 22001
rect 4582 21950 4660 21978
rect 4526 21927 4582 21936
rect 846 21856 902 21865
rect 846 21791 902 21800
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 2318 21856 2374 21865
rect 2318 21791 2374 21800
rect 3238 21856 3294 21865
rect 3238 21791 3294 21800
rect 3790 21856 3846 21865
rect 3790 21791 3846 21800
rect 860 21690 888 21791
rect 1596 21690 1624 21791
rect 2332 21690 2360 21791
rect 3252 21690 3280 21791
rect 3804 21690 3832 21791
rect 4285 21788 4593 21797
rect 4285 21786 4291 21788
rect 4347 21786 4371 21788
rect 4427 21786 4451 21788
rect 4507 21786 4531 21788
rect 4587 21786 4593 21788
rect 4347 21734 4349 21786
rect 4529 21734 4531 21786
rect 4285 21732 4291 21734
rect 4347 21732 4371 21734
rect 4427 21732 4451 21734
rect 4507 21732 4531 21734
rect 4587 21732 4593 21734
rect 4285 21723 4593 21732
rect 4632 21690 4660 21950
rect 8206 21927 8262 21936
rect 28998 21992 29054 22001
rect 28998 21927 29054 21936
rect 5262 21856 5318 21865
rect 5262 21791 5318 21800
rect 5998 21856 6054 21865
rect 5998 21791 6054 21800
rect 6734 21856 6790 21865
rect 6734 21791 6790 21800
rect 7470 21856 7526 21865
rect 7470 21791 7526 21800
rect 5276 21690 5304 21791
rect 6012 21690 6040 21791
rect 6748 21690 6776 21791
rect 7484 21690 7512 21791
rect 8220 21690 8248 21927
rect 16304 21888 16356 21894
rect 8758 21856 8814 21865
rect 8758 21791 8814 21800
rect 9678 21856 9734 21865
rect 9678 21791 9734 21800
rect 10414 21856 10470 21865
rect 10414 21791 10470 21800
rect 11150 21856 11206 21865
rect 16304 21830 16356 21836
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 25870 21856 25926 21865
rect 11150 21791 11206 21800
rect 8772 21690 8800 21791
rect 9692 21690 9720 21791
rect 10428 21690 10456 21791
rect 11164 21690 11192 21791
rect 12059 21788 12367 21797
rect 12059 21786 12065 21788
rect 12121 21786 12145 21788
rect 12201 21786 12225 21788
rect 12281 21786 12305 21788
rect 12361 21786 12367 21788
rect 12121 21734 12123 21786
rect 12303 21734 12305 21786
rect 12059 21732 12065 21734
rect 12121 21732 12145 21734
rect 12201 21732 12225 21734
rect 12281 21732 12305 21734
rect 12361 21732 12367 21734
rect 12059 21723 12367 21732
rect 16316 21690 16344 21830
rect 19833 21788 20141 21797
rect 19833 21786 19839 21788
rect 19895 21786 19919 21788
rect 19975 21786 19999 21788
rect 20055 21786 20079 21788
rect 20135 21786 20141 21788
rect 19895 21734 19897 21786
rect 20077 21734 20079 21786
rect 19833 21732 19839 21734
rect 19895 21732 19919 21734
rect 19975 21732 19999 21734
rect 20055 21732 20079 21734
rect 20135 21732 20141 21734
rect 19833 21723 20141 21732
rect 23952 21690 23980 21830
rect 25870 21791 25926 21800
rect 26790 21856 26846 21865
rect 26790 21791 26846 21800
rect 28538 21856 28594 21865
rect 848 21684 900 21690
rect 848 21626 900 21632
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8760 21684 8812 21690
rect 8760 21626 8812 21632
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 14648 21616 14700 21622
rect 11886 21584 11942 21593
rect 11886 21519 11942 21528
rect 13358 21584 13414 21593
rect 14648 21558 14700 21564
rect 13358 21519 13414 21528
rect 14372 21548 14424 21554
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 4285 20700 4593 20709
rect 4285 20698 4291 20700
rect 4347 20698 4371 20700
rect 4427 20698 4451 20700
rect 4507 20698 4531 20700
rect 4587 20698 4593 20700
rect 4347 20646 4349 20698
rect 4529 20646 4531 20698
rect 4285 20644 4291 20646
rect 4347 20644 4371 20646
rect 4427 20644 4451 20646
rect 4507 20644 4531 20646
rect 4587 20644 4593 20646
rect 4285 20635 4593 20644
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5092 19922 5120 20334
rect 6460 20324 6512 20330
rect 6460 20266 6512 20272
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 2976 19514 3004 19858
rect 3344 19514 3372 19858
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3608 19440 3660 19446
rect 3608 19382 3660 19388
rect 2412 18828 2464 18834
rect 3620 18816 3648 19382
rect 3712 19310 3740 19654
rect 4172 19310 4200 19654
rect 4285 19612 4593 19621
rect 4285 19610 4291 19612
rect 4347 19610 4371 19612
rect 4427 19610 4451 19612
rect 4507 19610 4531 19612
rect 4587 19610 4593 19612
rect 4347 19558 4349 19610
rect 4529 19558 4531 19610
rect 4285 19556 4291 19558
rect 4347 19556 4371 19558
rect 4427 19556 4451 19558
rect 4507 19556 4531 19558
rect 4587 19556 4593 19558
rect 4285 19547 4593 19556
rect 4632 19514 4660 19654
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4344 19168 4396 19174
rect 4080 19128 4344 19156
rect 4080 18834 4108 19128
rect 4344 19110 4396 19116
rect 3976 18828 4028 18834
rect 3620 18788 3976 18816
rect 2412 18770 2464 18776
rect 3976 18770 4028 18776
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 1216 17536 1268 17542
rect 1216 17478 1268 17484
rect 1228 17134 1256 17478
rect 1216 17128 1268 17134
rect 1216 17070 1268 17076
rect 1228 16574 1256 17070
rect 1492 17060 1544 17066
rect 1492 17002 1544 17008
rect 2228 17060 2280 17066
rect 2228 17002 2280 17008
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1504 16794 1532 17002
rect 2240 16794 2268 17002
rect 1492 16788 1544 16794
rect 1492 16730 1544 16736
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2424 16658 2452 18770
rect 4080 18630 4108 18770
rect 4632 18766 4660 19450
rect 4724 18834 4752 19722
rect 5184 19310 5212 20198
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4816 18766 4844 19246
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4804 18760 4856 18766
rect 5000 18737 5028 19246
rect 5276 19242 5304 19654
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5080 18760 5132 18766
rect 4804 18702 4856 18708
rect 4986 18728 5042 18737
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4080 18222 4108 18566
rect 4285 18524 4593 18533
rect 4285 18522 4291 18524
rect 4347 18522 4371 18524
rect 4427 18522 4451 18524
rect 4507 18522 4531 18524
rect 4587 18522 4593 18524
rect 4347 18470 4349 18522
rect 4529 18470 4531 18522
rect 4285 18468 4291 18470
rect 4347 18468 4371 18470
rect 4427 18468 4451 18470
rect 4507 18468 4531 18470
rect 4587 18468 4593 18470
rect 4285 18459 4593 18468
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4264 17882 4292 18362
rect 4436 18284 4488 18290
rect 4632 18272 4660 18702
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4488 18244 4660 18272
rect 4436 18226 4488 18232
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4356 17746 4384 18158
rect 4724 18086 4752 18566
rect 4816 18086 4844 18702
rect 5080 18702 5132 18708
rect 4986 18663 5042 18672
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4908 18222 4936 18566
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4724 17762 4752 18022
rect 4540 17746 4752 17762
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4528 17740 4752 17746
rect 4580 17734 4752 17740
rect 4528 17682 4580 17688
rect 4285 17436 4593 17445
rect 4285 17434 4291 17436
rect 4347 17434 4371 17436
rect 4427 17434 4451 17436
rect 4507 17434 4531 17436
rect 4587 17434 4593 17436
rect 4347 17382 4349 17434
rect 4529 17382 4531 17434
rect 4285 17380 4291 17382
rect 4347 17380 4371 17382
rect 4427 17380 4451 17382
rect 4507 17380 4531 17382
rect 4587 17380 4593 17382
rect 4285 17371 4593 17380
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3344 16658 3372 17070
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 1136 16546 1256 16574
rect 1308 16584 1360 16590
rect 1136 16114 1164 16546
rect 1308 16526 1360 16532
rect 1124 16108 1176 16114
rect 1124 16050 1176 16056
rect 1136 15586 1164 16050
rect 1216 16040 1268 16046
rect 1216 15982 1268 15988
rect 1228 15706 1256 15982
rect 1320 15910 1348 16526
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2608 15978 2636 16390
rect 2596 15972 2648 15978
rect 2596 15914 2648 15920
rect 1308 15904 1360 15910
rect 1308 15846 1360 15852
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 1320 15706 1348 15846
rect 2424 15706 2452 15846
rect 1216 15700 1268 15706
rect 1216 15642 1268 15648
rect 1308 15700 1360 15706
rect 1308 15642 1360 15648
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3700 15700 3752 15706
rect 3804 15688 3832 16594
rect 4285 16348 4593 16357
rect 4285 16346 4291 16348
rect 4347 16346 4371 16348
rect 4427 16346 4451 16348
rect 4507 16346 4531 16348
rect 4587 16346 4593 16348
rect 4347 16294 4349 16346
rect 4529 16294 4531 16346
rect 4285 16292 4291 16294
rect 4347 16292 4371 16294
rect 4427 16292 4451 16294
rect 4507 16292 4531 16294
rect 4587 16292 4593 16294
rect 4285 16283 4593 16292
rect 3752 15660 3832 15688
rect 3700 15642 3752 15648
rect 1136 15558 1348 15586
rect 1320 14550 1348 15558
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1308 14544 1360 14550
rect 1308 14486 1360 14492
rect 1032 14272 1084 14278
rect 1032 14214 1084 14220
rect 1044 13870 1072 14214
rect 1320 14006 1348 14486
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 14074 1440 14350
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1308 14000 1360 14006
rect 1308 13942 1360 13948
rect 1032 13864 1084 13870
rect 1032 13806 1084 13812
rect 1320 13462 1348 13942
rect 1688 13938 1716 15302
rect 2056 14278 2084 15370
rect 2976 14958 3004 15438
rect 3068 14958 3096 15642
rect 4724 15570 4752 17734
rect 4816 16726 4844 18022
rect 4908 17882 4936 18158
rect 5000 17882 5028 18663
rect 5092 18154 5120 18702
rect 5184 18154 5212 18770
rect 5276 18698 5304 19178
rect 5368 18873 5396 19858
rect 5460 19786 5488 20198
rect 6196 20058 6224 20198
rect 6472 20058 6500 20266
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5460 18970 5488 19722
rect 5644 19514 5672 19790
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5920 19446 5948 19926
rect 6656 19922 6684 21422
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8172 21244 8480 21253
rect 8172 21242 8178 21244
rect 8234 21242 8258 21244
rect 8314 21242 8338 21244
rect 8394 21242 8418 21244
rect 8474 21242 8480 21244
rect 8234 21190 8236 21242
rect 8416 21190 8418 21242
rect 8172 21188 8178 21190
rect 8234 21188 8258 21190
rect 8314 21188 8338 21190
rect 8394 21188 8418 21190
rect 8474 21188 8480 21190
rect 8172 21179 8480 21188
rect 8772 20942 8800 21286
rect 11440 21146 11468 21354
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 8852 21004 8904 21010
rect 8852 20946 8904 20952
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 8772 20466 8800 20878
rect 8864 20602 8892 20946
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 9876 20398 9904 20946
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10244 20398 10272 20742
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 7196 20324 7248 20330
rect 7196 20266 7248 20272
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6092 19712 6144 19718
rect 6092 19654 6144 19660
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5920 19334 5948 19382
rect 5920 19306 6040 19334
rect 6104 19310 6132 19654
rect 5630 19000 5686 19009
rect 5448 18964 5500 18970
rect 5630 18935 5686 18944
rect 5448 18906 5500 18912
rect 5644 18902 5672 18935
rect 5632 18896 5684 18902
rect 5354 18864 5410 18873
rect 5632 18838 5684 18844
rect 6012 18834 6040 19306
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6380 19292 6408 19858
rect 6460 19304 6512 19310
rect 6380 19264 6460 19292
rect 5354 18799 5356 18808
rect 5408 18799 5410 18808
rect 6000 18828 6052 18834
rect 5356 18770 5408 18776
rect 6000 18770 6052 18776
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 5092 17746 5120 18090
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5000 17134 5028 17682
rect 5080 17196 5132 17202
rect 5184 17184 5212 17818
rect 5276 17746 5304 18022
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5460 17610 5488 18158
rect 5920 17746 5948 18226
rect 5908 17740 5960 17746
rect 6012 17728 6040 18770
rect 6092 18284 6144 18290
rect 6196 18272 6224 18770
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 6380 18748 6408 19264
rect 6460 19246 6512 19252
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 19009 6500 19110
rect 6458 19000 6514 19009
rect 6458 18935 6514 18944
rect 6550 18864 6606 18873
rect 6550 18799 6552 18808
rect 6604 18799 6606 18808
rect 6552 18770 6604 18776
rect 6460 18760 6512 18766
rect 6380 18720 6460 18748
rect 6144 18244 6224 18272
rect 6092 18226 6144 18232
rect 6288 18086 6316 18702
rect 6380 18630 6408 18720
rect 6460 18702 6512 18708
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6092 17740 6144 17746
rect 6012 17700 6092 17728
rect 5908 17682 5960 17688
rect 6092 17682 6144 17688
rect 6472 17678 6500 18158
rect 6460 17672 6512 17678
rect 6656 17626 6684 19858
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6748 18698 6776 19246
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18873 6868 19110
rect 6826 18864 6882 18873
rect 6826 18799 6882 18808
rect 6826 18728 6882 18737
rect 6736 18692 6788 18698
rect 6826 18663 6828 18672
rect 6736 18634 6788 18640
rect 6880 18663 6882 18672
rect 6828 18634 6880 18640
rect 6932 18290 6960 19246
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7116 18970 7144 19110
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7104 18760 7156 18766
rect 7208 18748 7236 20266
rect 8172 20156 8480 20165
rect 8172 20154 8178 20156
rect 8234 20154 8258 20156
rect 8314 20154 8338 20156
rect 8394 20154 8418 20156
rect 8474 20154 8480 20156
rect 8234 20102 8236 20154
rect 8416 20102 8418 20154
rect 8172 20100 8178 20102
rect 8234 20100 8258 20102
rect 8314 20100 8338 20102
rect 8394 20100 8418 20102
rect 8474 20100 8480 20102
rect 8172 20091 8480 20100
rect 8864 19922 8892 20334
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 9048 19922 9076 20198
rect 9220 19984 9272 19990
rect 9218 19952 9220 19961
rect 9272 19952 9274 19961
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 9036 19916 9088 19922
rect 9416 19922 9444 20334
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 20058 9812 20198
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9218 19887 9274 19896
rect 9404 19916 9456 19922
rect 9036 19858 9088 19864
rect 9404 19858 9456 19864
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7156 18720 7236 18748
rect 7104 18702 7156 18708
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6460 17614 6512 17620
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 6564 17598 6684 17626
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 5132 17156 5212 17184
rect 5080 17138 5132 17144
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 3896 15434 3924 15506
rect 3884 15428 3936 15434
rect 3884 15370 3936 15376
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2884 14278 2912 14758
rect 3068 14618 3096 14758
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 3252 13530 3280 14282
rect 3344 14006 3372 14894
rect 3436 14482 3464 15302
rect 4285 15260 4593 15269
rect 4285 15258 4291 15260
rect 4347 15258 4371 15260
rect 4427 15258 4451 15260
rect 4507 15258 4531 15260
rect 4587 15258 4593 15260
rect 4347 15206 4349 15258
rect 4529 15206 4531 15258
rect 4285 15204 4291 15206
rect 4347 15204 4371 15206
rect 4427 15204 4451 15206
rect 4507 15204 4531 15206
rect 4587 15204 4593 15206
rect 4285 15195 4593 15204
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 3620 14618 3648 14826
rect 4356 14618 4384 14826
rect 4816 14618 4844 16662
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 5000 15026 5028 15982
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 5092 15434 5120 15914
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5080 15428 5132 15434
rect 5080 15370 5132 15376
rect 5092 15162 5120 15370
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4172 14006 4200 14350
rect 4285 14172 4593 14181
rect 4285 14170 4291 14172
rect 4347 14170 4371 14172
rect 4427 14170 4451 14172
rect 4507 14170 4531 14172
rect 4587 14170 4593 14172
rect 4347 14118 4349 14170
rect 4529 14118 4531 14170
rect 4285 14116 4291 14118
rect 4347 14116 4371 14118
rect 4427 14116 4451 14118
rect 4507 14116 4531 14118
rect 4587 14116 4593 14118
rect 4285 14107 4593 14116
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 1308 13456 1360 13462
rect 1308 13398 1360 13404
rect 3344 13326 3372 13942
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13462 3832 13670
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 1412 12986 1440 13262
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 2884 12782 2912 13126
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2872 12640 2924 12646
rect 2792 12600 2872 12628
rect 2792 12170 2820 12600
rect 2872 12582 2924 12588
rect 3068 12442 3096 12650
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3344 12238 3372 13262
rect 4172 12986 4200 13806
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4285 13084 4593 13093
rect 4285 13082 4291 13084
rect 4347 13082 4371 13084
rect 4427 13082 4451 13084
rect 4507 13082 4531 13084
rect 4587 13082 4593 13084
rect 4347 13030 4349 13082
rect 4529 13030 4531 13082
rect 4285 13028 4291 13030
rect 4347 13028 4371 13030
rect 4427 13028 4451 13030
rect 4507 13028 4531 13030
rect 4587 13028 4593 13030
rect 4285 13019 4593 13028
rect 4724 12986 4752 13398
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4816 12782 4844 14554
rect 5460 14482 5488 14962
rect 5552 14958 5580 15302
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5460 13938 5488 14418
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5184 13530 5212 13806
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5276 12986 5304 13806
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 3608 12776 3660 12782
rect 4804 12776 4856 12782
rect 3608 12718 3660 12724
rect 4632 12736 4804 12764
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11150 2820 12106
rect 3344 11150 3372 12174
rect 3436 11354 3464 12650
rect 3620 12434 3648 12718
rect 4068 12436 4120 12442
rect 3620 12406 4068 12434
rect 3620 12374 3648 12406
rect 4068 12378 4120 12384
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 4285 11996 4593 12005
rect 4285 11994 4291 11996
rect 4347 11994 4371 11996
rect 4427 11994 4451 11996
rect 4507 11994 4531 11996
rect 4587 11994 4593 11996
rect 4347 11942 4349 11994
rect 4529 11942 4531 11994
rect 4285 11940 4291 11942
rect 4347 11940 4371 11942
rect 4427 11940 4451 11942
rect 4507 11940 4531 11942
rect 4587 11940 4593 11942
rect 4285 11931 4593 11940
rect 4632 11694 4660 12736
rect 4804 12718 4856 12724
rect 5172 12776 5224 12782
rect 5552 12730 5580 13330
rect 5644 12986 5672 13330
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5172 12718 5224 12724
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4724 11898 4752 12310
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 5184 11694 5212 12718
rect 5460 12702 5580 12730
rect 5736 12714 5764 15506
rect 6472 15348 6500 17478
rect 6564 16114 6592 17598
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6656 17202 6684 17478
rect 6748 17338 6776 17614
rect 6932 17610 6960 18226
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7024 17746 7052 18022
rect 7208 17814 7236 18720
rect 7484 18086 7512 19314
rect 8588 19310 8616 19654
rect 8680 19514 8708 19790
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8864 19310 8892 19858
rect 8942 19816 8998 19825
rect 8942 19751 8998 19760
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 8576 19304 8628 19310
rect 8760 19304 8812 19310
rect 8576 19246 8628 19252
rect 8758 19272 8760 19281
rect 8852 19304 8904 19310
rect 8812 19272 8814 19281
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7576 17864 7604 18158
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7300 17836 7604 17864
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7196 17672 7248 17678
rect 7300 17660 7328 17836
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7248 17632 7328 17660
rect 7196 17614 7248 17620
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6840 17218 6868 17478
rect 7116 17218 7144 17546
rect 6644 17196 6696 17202
rect 6840 17190 7144 17218
rect 6644 17138 6696 17144
rect 7116 17134 7144 17190
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7024 16794 7052 17070
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 15502 6592 16050
rect 7116 16046 7144 16934
rect 7392 16658 7420 17682
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7484 15706 7512 16526
rect 7576 16522 7604 17836
rect 7760 17814 7788 18022
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7668 17066 7696 17138
rect 7760 17134 7788 17478
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7668 16658 7696 16730
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 16250 7788 16390
rect 7852 16250 7880 16526
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6472 15320 6592 15348
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 13394 5948 13738
rect 6104 13530 6132 14418
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 6472 13326 6500 13806
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12986 5856 13126
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5724 12708 5776 12714
rect 5356 12436 5408 12442
rect 5460 12434 5488 12702
rect 5724 12650 5776 12656
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6104 12442 6132 12582
rect 5408 12406 5488 12434
rect 6092 12436 6144 12442
rect 5356 12378 5408 12384
rect 6092 12378 6144 12384
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11694 6040 12038
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 5736 11150 5764 11562
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11286 5856 11494
rect 6288 11354 6316 13194
rect 6472 12850 6500 13262
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6380 12238 6408 12650
rect 6564 12238 6592 15320
rect 7392 15026 7420 15506
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7564 14952 7616 14958
rect 6826 14920 6882 14929
rect 7564 14894 7616 14900
rect 6826 14855 6882 14864
rect 6840 14822 6868 14855
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 14618 7512 14758
rect 7576 14618 7604 14894
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7668 14482 7696 15438
rect 7852 15094 7880 15506
rect 7944 15162 7972 18226
rect 8036 18086 8064 19246
rect 8852 19246 8904 19252
rect 8758 19207 8814 19216
rect 8956 19174 8984 19751
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8172 19068 8480 19077
rect 8172 19066 8178 19068
rect 8234 19066 8258 19068
rect 8314 19066 8338 19068
rect 8394 19066 8418 19068
rect 8474 19066 8480 19068
rect 8234 19014 8236 19066
rect 8416 19014 8418 19066
rect 8172 19012 8178 19014
rect 8234 19012 8258 19014
rect 8314 19012 8338 19014
rect 8394 19012 8418 19014
rect 8474 19012 8480 19014
rect 8172 19003 8480 19012
rect 9048 18902 9076 19858
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19514 9352 19790
rect 9876 19786 9904 20334
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9692 19446 9720 19722
rect 9784 19514 9812 19722
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9772 19304 9824 19310
rect 9864 19304 9916 19310
rect 9772 19246 9824 19252
rect 9862 19272 9864 19281
rect 9916 19272 9918 19281
rect 9324 19145 9352 19246
rect 9310 19136 9366 19145
rect 9310 19071 9366 19080
rect 9218 19000 9274 19009
rect 9218 18935 9274 18944
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 8482 18728 8538 18737
rect 9232 18698 9260 18935
rect 8482 18663 8484 18672
rect 8536 18663 8538 18672
rect 9220 18692 9272 18698
rect 8484 18634 8536 18640
rect 9220 18634 9272 18640
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 8172 17980 8480 17989
rect 8172 17978 8178 17980
rect 8234 17978 8258 17980
rect 8314 17978 8338 17980
rect 8394 17978 8418 17980
rect 8474 17978 8480 17980
rect 8234 17926 8236 17978
rect 8416 17926 8418 17978
rect 8172 17924 8178 17926
rect 8234 17924 8258 17926
rect 8314 17924 8338 17926
rect 8394 17924 8418 17926
rect 8474 17924 8480 17926
rect 8172 17915 8480 17924
rect 8172 16892 8480 16901
rect 8172 16890 8178 16892
rect 8234 16890 8258 16892
rect 8314 16890 8338 16892
rect 8394 16890 8418 16892
rect 8474 16890 8480 16892
rect 8234 16838 8236 16890
rect 8416 16838 8418 16890
rect 8172 16836 8178 16838
rect 8234 16836 8258 16838
rect 8314 16836 8338 16838
rect 8394 16836 8418 16838
rect 8474 16836 8480 16838
rect 8172 16827 8480 16836
rect 9048 16046 9076 18566
rect 9324 18426 9352 19071
rect 9416 18970 9444 19246
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9416 18426 9444 18770
rect 9508 18698 9536 19178
rect 9600 19009 9628 19246
rect 9586 19000 9642 19009
rect 9586 18935 9642 18944
rect 9692 18834 9720 19246
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9784 18426 9812 19246
rect 9862 19207 9918 19216
rect 9864 19168 9916 19174
rect 9968 19145 9996 19926
rect 10060 19378 10088 19994
rect 10416 19916 10468 19922
rect 10468 19876 10548 19904
rect 10416 19858 10468 19864
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 9864 19110 9916 19116
rect 9954 19136 10010 19145
rect 9876 18952 9904 19110
rect 10010 19094 10088 19122
rect 9954 19071 10010 19080
rect 9876 18924 9996 18952
rect 9864 18850 9916 18856
rect 9864 18792 9916 18798
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9876 18358 9904 18792
rect 9968 18766 9996 18924
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 10060 18630 10088 19094
rect 10520 18952 10548 19876
rect 10428 18924 10548 18952
rect 10324 18828 10376 18834
rect 10244 18788 10324 18816
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10244 18426 10272 18788
rect 10324 18770 10376 18776
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10336 18358 10364 18566
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9600 17762 9628 18090
rect 9784 17882 9812 18090
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9600 17746 9720 17762
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9588 17740 9720 17746
rect 9640 17734 9720 17740
rect 9588 17682 9640 17688
rect 9416 17542 9444 17682
rect 9586 17640 9642 17649
rect 9586 17575 9642 17584
rect 9692 17626 9720 17734
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9692 17598 9904 17626
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9600 17338 9628 17575
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9692 16250 9720 17598
rect 9876 17542 9904 17598
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9784 17338 9812 17478
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9968 17270 9996 17682
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9968 16794 9996 17206
rect 10060 17134 10088 18158
rect 10152 17882 10180 18226
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10428 17814 10456 18924
rect 10612 18834 10640 19994
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10244 17542 10272 17750
rect 10428 17542 10456 17750
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10520 17338 10548 18362
rect 10796 18290 10824 19654
rect 10888 19242 10916 20742
rect 10980 19990 11008 20946
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 11072 19514 11100 20946
rect 11532 20602 11560 21422
rect 11900 21010 11928 21519
rect 13372 21146 13400 21519
rect 14372 21490 14424 21496
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12059 20700 12367 20709
rect 12059 20698 12065 20700
rect 12121 20698 12145 20700
rect 12201 20698 12225 20700
rect 12281 20698 12305 20700
rect 12361 20698 12367 20700
rect 12121 20646 12123 20698
rect 12303 20646 12305 20698
rect 12059 20644 12065 20646
rect 12121 20644 12145 20646
rect 12201 20644 12225 20646
rect 12281 20644 12305 20646
rect 12361 20644 12367 20646
rect 12059 20635 12367 20644
rect 12820 20602 12848 20742
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 11440 19514 11468 20334
rect 11532 19718 11560 20538
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11256 19394 11284 19450
rect 11072 19378 11284 19394
rect 11060 19372 11284 19378
rect 11112 19366 11284 19372
rect 11060 19314 11112 19320
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10980 18970 11008 19178
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 18358 10916 18566
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10612 17746 10640 18226
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10704 17882 10732 18158
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10704 17338 10732 17546
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 10428 17134 10456 17206
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 8116 16040 8168 16046
rect 8036 15988 8116 15994
rect 8036 15982 8168 15988
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8036 15966 8156 15982
rect 8036 15570 8064 15966
rect 8172 15804 8480 15813
rect 8172 15802 8178 15804
rect 8234 15802 8258 15804
rect 8314 15802 8338 15804
rect 8394 15802 8418 15804
rect 8474 15802 8480 15804
rect 8234 15750 8236 15802
rect 8416 15750 8418 15802
rect 8172 15748 8178 15750
rect 8234 15748 8258 15750
rect 8314 15748 8338 15750
rect 8394 15748 8418 15750
rect 8474 15748 8480 15750
rect 8172 15739 8480 15748
rect 8680 15570 8708 15982
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7840 14952 7892 14958
rect 7944 14940 7972 15098
rect 9324 14958 9352 15506
rect 9692 15162 9720 16186
rect 10336 16046 10364 16594
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10244 15502 10272 15982
rect 10428 15570 10456 17070
rect 10520 16658 10548 17138
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 10612 16794 10640 17002
rect 10704 16794 10732 17274
rect 10796 17116 10824 18226
rect 10968 18148 11020 18154
rect 11072 18136 11100 18770
rect 11150 18728 11206 18737
rect 11150 18663 11152 18672
rect 11204 18663 11206 18672
rect 11152 18634 11204 18640
rect 11020 18108 11100 18136
rect 10968 18090 11020 18096
rect 11072 17882 11100 18108
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10876 17128 10928 17134
rect 10796 17088 10876 17116
rect 10876 17070 10928 17076
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10796 16522 10824 16662
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10784 15972 10836 15978
rect 10968 15972 11020 15978
rect 10836 15932 10968 15960
rect 10784 15914 10836 15920
rect 10968 15914 11020 15920
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 7892 14912 7972 14940
rect 8668 14952 8720 14958
rect 7840 14894 7892 14900
rect 8668 14894 8720 14900
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7194 14376 7250 14385
rect 7194 14311 7196 14320
rect 7248 14311 7250 14320
rect 7196 14282 7248 14288
rect 7760 14074 7788 14894
rect 8172 14716 8480 14725
rect 8172 14714 8178 14716
rect 8234 14714 8258 14716
rect 8314 14714 8338 14716
rect 8394 14714 8418 14716
rect 8474 14714 8480 14716
rect 8234 14662 8236 14714
rect 8416 14662 8418 14714
rect 8172 14660 8178 14662
rect 8234 14660 8258 14662
rect 8314 14660 8338 14662
rect 8394 14660 8418 14662
rect 8474 14660 8480 14662
rect 8172 14651 8480 14660
rect 8680 14550 8708 14894
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 9232 14346 9260 14758
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 8172 13628 8480 13637
rect 8172 13626 8178 13628
rect 8234 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8480 13628
rect 8234 13574 8236 13626
rect 8416 13574 8418 13626
rect 8172 13572 8178 13574
rect 8234 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8480 13574
rect 8172 13563 8480 13572
rect 9324 13190 9352 14894
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9416 14278 9444 14418
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9508 14074 9536 14758
rect 10244 14618 10272 14826
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10520 14498 10548 15098
rect 10980 14958 11008 15438
rect 10968 14952 11020 14958
rect 11020 14900 11192 14906
rect 10968 14894 11192 14900
rect 10980 14878 11192 14894
rect 10520 14482 11008 14498
rect 10508 14476 11008 14482
rect 10560 14470 11008 14476
rect 10508 14418 10560 14424
rect 10980 14414 11008 14470
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 9784 14074 9812 14350
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10244 14074 10272 14214
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10336 13870 10364 14214
rect 10428 14074 10456 14282
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10704 13734 10732 13942
rect 10796 13734 10824 14282
rect 11072 14074 11100 14282
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11164 13852 11192 14878
rect 11256 14482 11284 19366
rect 11532 19310 11560 19654
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11520 18148 11572 18154
rect 11520 18090 11572 18096
rect 11334 17776 11390 17785
rect 11532 17746 11560 18090
rect 11334 17711 11336 17720
rect 11388 17711 11390 17720
rect 11520 17740 11572 17746
rect 11336 17682 11388 17688
rect 11520 17682 11572 17688
rect 11336 14544 11388 14550
rect 11520 14544 11572 14550
rect 11388 14504 11520 14532
rect 11336 14486 11388 14492
rect 11520 14486 11572 14492
rect 11624 14482 11652 20198
rect 11716 18834 11744 20334
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12059 19612 12367 19621
rect 12059 19610 12065 19612
rect 12121 19610 12145 19612
rect 12201 19610 12225 19612
rect 12281 19610 12305 19612
rect 12361 19610 12367 19612
rect 12121 19558 12123 19610
rect 12303 19558 12305 19610
rect 12059 19556 12065 19558
rect 12121 19556 12145 19558
rect 12201 19556 12225 19558
rect 12281 19556 12305 19558
rect 12361 19556 12367 19558
rect 12059 19547 12367 19556
rect 12728 19514 12756 19654
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12059 18524 12367 18533
rect 12059 18522 12065 18524
rect 12121 18522 12145 18524
rect 12201 18522 12225 18524
rect 12281 18522 12305 18524
rect 12361 18522 12367 18524
rect 12121 18470 12123 18522
rect 12303 18470 12305 18522
rect 12059 18468 12065 18470
rect 12121 18468 12145 18470
rect 12201 18468 12225 18470
rect 12281 18468 12305 18470
rect 12361 18468 12367 18470
rect 12059 18459 12367 18468
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17649 11744 17682
rect 12452 17678 12480 18294
rect 12820 17882 12848 18770
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12912 17762 12940 20742
rect 13556 20534 13584 20878
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 19922 13492 20198
rect 13544 19984 13596 19990
rect 13542 19952 13544 19961
rect 13596 19952 13598 19961
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13268 19916 13320 19922
rect 13452 19916 13504 19922
rect 13268 19858 13320 19864
rect 13372 19876 13452 19904
rect 13188 19786 13216 19858
rect 13280 19825 13308 19858
rect 13266 19816 13322 19825
rect 13176 19780 13228 19786
rect 13266 19751 13322 19760
rect 13176 19722 13228 19728
rect 13188 18986 13216 19722
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 13004 18958 13216 18986
rect 13004 18766 13032 18958
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13176 18828 13228 18834
rect 13280 18816 13308 19382
rect 13372 18902 13400 19876
rect 13542 19887 13598 19896
rect 13452 19858 13504 19864
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13556 18834 13584 19110
rect 13228 18788 13308 18816
rect 13452 18828 13504 18834
rect 13176 18770 13228 18776
rect 13452 18770 13504 18776
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13096 18426 13124 18770
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13188 18306 13216 18770
rect 13464 18630 13492 18770
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 12820 17734 12940 17762
rect 13096 18278 13216 18306
rect 12440 17672 12492 17678
rect 11702 17640 11758 17649
rect 12440 17614 12492 17620
rect 11702 17575 11758 17584
rect 12059 17436 12367 17445
rect 12059 17434 12065 17436
rect 12121 17434 12145 17436
rect 12201 17434 12225 17436
rect 12281 17434 12305 17436
rect 12361 17434 12367 17436
rect 12121 17382 12123 17434
rect 12303 17382 12305 17434
rect 12059 17380 12065 17382
rect 12121 17380 12145 17382
rect 12201 17380 12225 17382
rect 12281 17380 12305 17382
rect 12361 17380 12367 17382
rect 12059 17371 12367 17380
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11520 14408 11572 14414
rect 11518 14376 11520 14385
rect 11572 14376 11574 14385
rect 11518 14311 11574 14320
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 14074 11376 14214
rect 11624 14074 11652 14418
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11336 13864 11388 13870
rect 11164 13824 11336 13852
rect 11336 13806 11388 13812
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10704 13394 10732 13670
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 8312 12850 8340 13126
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 11348 12782 11376 13806
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6380 11898 6408 12174
rect 6748 12102 6776 12582
rect 7208 12306 7236 12650
rect 7300 12306 7328 12650
rect 8172 12540 8480 12549
rect 8172 12538 8178 12540
rect 8234 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8480 12540
rect 8234 12486 8236 12538
rect 8416 12486 8418 12538
rect 8172 12484 8178 12486
rect 8234 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8480 12486
rect 8172 12475 8480 12484
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6748 11558 6776 12038
rect 7208 11762 7236 12242
rect 7300 11778 7328 12242
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7300 11750 7512 11778
rect 8036 11762 8064 12242
rect 9416 12238 9444 12650
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 6564 11150 6592 11494
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 3332 11144 3384 11150
rect 3700 11144 3752 11150
rect 3384 11092 3700 11098
rect 3332 11086 3752 11092
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 3344 11070 3740 11086
rect 4285 10908 4593 10917
rect 4285 10906 4291 10908
rect 4347 10906 4371 10908
rect 4427 10906 4451 10908
rect 4507 10906 4531 10908
rect 4587 10906 4593 10908
rect 4347 10854 4349 10906
rect 4529 10854 4531 10906
rect 4285 10852 4291 10854
rect 4347 10852 4371 10854
rect 4427 10852 4451 10854
rect 4507 10852 4531 10854
rect 4587 10852 4593 10854
rect 4285 10843 4593 10852
rect 5736 10606 5764 11086
rect 6472 10674 6500 11086
rect 7116 10810 7144 11222
rect 7208 11082 7236 11698
rect 7300 11626 7328 11750
rect 7484 11694 7512 11750
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7484 10810 7512 11630
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11354 7604 11494
rect 8172 11452 8480 11461
rect 8172 11450 8178 11452
rect 8234 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8480 11452
rect 8234 11398 8236 11450
rect 8416 11398 8418 11450
rect 8172 11396 8178 11398
rect 8234 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8480 11398
rect 8172 11387 8480 11396
rect 8588 11354 8616 11630
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8680 11286 8708 11766
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7760 10674 7788 10950
rect 8680 10674 8708 11222
rect 8956 11218 8984 12038
rect 9416 11762 9444 12038
rect 10428 11898 10456 12242
rect 10980 12238 11008 12650
rect 11624 12646 11652 13330
rect 11992 12918 12020 17138
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12059 16348 12367 16357
rect 12059 16346 12065 16348
rect 12121 16346 12145 16348
rect 12201 16346 12225 16348
rect 12281 16346 12305 16348
rect 12361 16346 12367 16348
rect 12121 16294 12123 16346
rect 12303 16294 12305 16346
rect 12059 16292 12065 16294
rect 12121 16292 12145 16294
rect 12201 16292 12225 16294
rect 12281 16292 12305 16294
rect 12361 16292 12367 16294
rect 12059 16283 12367 16292
rect 12544 16114 12572 17002
rect 12532 16108 12584 16114
rect 12584 16068 12756 16096
rect 12532 16050 12584 16056
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12059 15260 12367 15269
rect 12059 15258 12065 15260
rect 12121 15258 12145 15260
rect 12201 15258 12225 15260
rect 12281 15258 12305 15260
rect 12361 15258 12367 15260
rect 12121 15206 12123 15258
rect 12303 15206 12305 15258
rect 12059 15204 12065 15206
rect 12121 15204 12145 15206
rect 12201 15204 12225 15206
rect 12281 15204 12305 15206
rect 12361 15204 12367 15206
rect 12059 15195 12367 15204
rect 12452 14958 12480 15302
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12544 14482 12572 15914
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12059 14172 12367 14181
rect 12059 14170 12065 14172
rect 12121 14170 12145 14172
rect 12201 14170 12225 14172
rect 12281 14170 12305 14172
rect 12361 14170 12367 14172
rect 12121 14118 12123 14170
rect 12303 14118 12305 14170
rect 12059 14116 12065 14118
rect 12121 14116 12145 14118
rect 12201 14116 12225 14118
rect 12281 14116 12305 14118
rect 12361 14116 12367 14118
rect 12059 14107 12367 14116
rect 12452 13258 12480 14418
rect 12544 14278 12572 14418
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12636 13394 12664 15506
rect 12728 15348 12756 16068
rect 12820 15502 12848 17734
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12728 15320 12848 15348
rect 12820 14482 12848 15320
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12728 14074 12756 14418
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12059 13084 12367 13093
rect 12059 13082 12065 13084
rect 12121 13082 12145 13084
rect 12201 13082 12225 13084
rect 12281 13082 12305 13084
rect 12361 13082 12367 13084
rect 12121 13030 12123 13082
rect 12303 13030 12305 13082
rect 12059 13028 12065 13030
rect 12121 13028 12145 13030
rect 12201 13028 12225 13030
rect 12281 13028 12305 13030
rect 12361 13028 12367 13030
rect 12059 13019 12367 13028
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 12728 12782 12756 13262
rect 12912 12986 12940 17614
rect 13096 16658 13124 18278
rect 13372 17882 13400 18566
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13188 17134 13216 17682
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13280 16658 13308 17682
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17338 13492 17478
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13556 16794 13584 17614
rect 13648 17082 13676 20334
rect 13726 19952 13782 19961
rect 13726 19887 13728 19896
rect 13780 19887 13782 19896
rect 13728 19858 13780 19864
rect 13832 19786 13860 21354
rect 14384 21350 14412 21490
rect 14660 21350 14688 21558
rect 16316 21486 16344 21626
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 25412 21616 25464 21622
rect 25412 21558 25464 21564
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 14384 21146 14412 21286
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 14094 20496 14150 20505
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 17746 13768 19654
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13832 18970 13860 19178
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13924 18834 13952 20470
rect 14094 20431 14096 20440
rect 14148 20431 14150 20440
rect 14096 20402 14148 20408
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14016 19514 14044 19790
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14200 18986 14228 20946
rect 14556 20936 14608 20942
rect 14660 20924 14688 21286
rect 14608 20896 14780 20924
rect 14556 20878 14608 20884
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14646 20768 14702 20777
rect 14568 20466 14596 20742
rect 14646 20703 14702 20712
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14280 19848 14332 19854
rect 14278 19816 14280 19825
rect 14332 19816 14334 19825
rect 14278 19751 14334 19760
rect 14200 18958 14320 18986
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 17338 13860 17478
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13728 17264 13780 17270
rect 13780 17212 13860 17218
rect 13728 17206 13860 17212
rect 13740 17190 13860 17206
rect 13648 17054 13768 17082
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13648 16726 13676 16934
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13004 13190 13032 16526
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 12728 12374 12756 12718
rect 13096 12442 13124 15914
rect 13188 15570 13216 16458
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 15570 13308 16390
rect 13450 16144 13506 16153
rect 13450 16079 13506 16088
rect 13464 15570 13492 16079
rect 13740 16046 13768 17054
rect 13832 16590 13860 17190
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 14016 16096 14044 16730
rect 14200 16250 14228 18770
rect 14292 17082 14320 18958
rect 14568 18902 14596 20402
rect 14660 18970 14688 20703
rect 14752 19242 14780 20896
rect 15028 20398 15056 21286
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15290 20496 15346 20505
rect 15290 20431 15346 20440
rect 15304 20398 15332 20431
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15120 20058 15148 20334
rect 15488 20058 15516 20538
rect 15764 20466 15792 21082
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 14830 19952 14886 19961
rect 15106 19952 15162 19961
rect 14886 19910 15056 19938
rect 14830 19887 14886 19896
rect 15028 19258 15056 19910
rect 15106 19887 15108 19896
rect 15160 19887 15162 19896
rect 15108 19858 15160 19864
rect 15764 19378 15792 20402
rect 15856 19718 15884 21286
rect 15946 21244 16254 21253
rect 15946 21242 15952 21244
rect 16008 21242 16032 21244
rect 16088 21242 16112 21244
rect 16168 21242 16192 21244
rect 16248 21242 16254 21244
rect 16008 21190 16010 21242
rect 16190 21190 16192 21242
rect 15946 21188 15952 21190
rect 16008 21188 16032 21190
rect 16088 21188 16112 21190
rect 16168 21188 16192 21190
rect 16248 21188 16254 21190
rect 15946 21179 16254 21188
rect 16684 21146 16712 21490
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 17130 21312 17186 21321
rect 17130 21247 17186 21256
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 15946 20156 16254 20165
rect 15946 20154 15952 20156
rect 16008 20154 16032 20156
rect 16088 20154 16112 20156
rect 16168 20154 16192 20156
rect 16248 20154 16254 20156
rect 16008 20102 16010 20154
rect 16190 20102 16192 20154
rect 15946 20100 15952 20102
rect 16008 20100 16032 20102
rect 16088 20100 16112 20102
rect 16168 20100 16192 20102
rect 16248 20100 16254 20102
rect 15946 20091 16254 20100
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 14740 19236 14792 19242
rect 15028 19230 15148 19258
rect 14740 19178 14792 19184
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14568 18154 14596 18838
rect 14752 18766 14780 19178
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17338 14412 17478
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14568 17202 14596 18090
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14292 17054 14412 17082
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 13924 16068 14044 16096
rect 14096 16108 14148 16114
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13648 15638 13676 15982
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15722 13860 15846
rect 13740 15694 13860 15722
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13740 15570 13768 15694
rect 13924 15570 13952 16068
rect 14096 16050 14148 16056
rect 14108 15994 14136 16050
rect 14016 15966 14136 15994
rect 14188 15972 14240 15978
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 13188 15094 13216 15370
rect 13832 15162 13860 15506
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13924 15008 13952 15506
rect 14016 15502 14044 15966
rect 14188 15914 14240 15920
rect 14200 15706 14228 15914
rect 14292 15706 14320 16526
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13832 14980 13952 15008
rect 13544 14952 13596 14958
rect 13636 14952 13688 14958
rect 13544 14894 13596 14900
rect 13634 14920 13636 14929
rect 13688 14920 13690 14929
rect 13556 14618 13584 14894
rect 13634 14855 13690 14864
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13740 14482 13768 14758
rect 13832 14482 13860 14980
rect 14108 14958 14136 15506
rect 14200 15162 14228 15506
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8956 10606 8984 11154
rect 9416 10606 9444 11698
rect 10428 11354 10456 11834
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 10520 10554 10548 11494
rect 11072 11150 11100 11494
rect 11164 11218 11192 12038
rect 12059 11996 12367 12005
rect 12059 11994 12065 11996
rect 12121 11994 12145 11996
rect 12201 11994 12225 11996
rect 12281 11994 12305 11996
rect 12361 11994 12367 11996
rect 12121 11942 12123 11994
rect 12303 11942 12305 11994
rect 12059 11940 12065 11942
rect 12121 11940 12145 11942
rect 12201 11940 12225 11942
rect 12281 11940 12305 11942
rect 12361 11940 12367 11942
rect 12059 11931 12367 11940
rect 13188 11558 13216 12650
rect 13372 11694 13400 13330
rect 13924 12986 13952 14826
rect 14108 14482 14136 14894
rect 14200 14618 14228 14894
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14384 14550 14412 17054
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14476 15706 14504 16118
rect 14568 16046 14596 17138
rect 14660 16114 14688 18634
rect 14752 18290 14780 18702
rect 15028 18630 15056 19110
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14738 17912 14794 17921
rect 14936 17882 14964 18022
rect 14738 17847 14794 17856
rect 14924 17876 14976 17882
rect 14752 17338 14780 17847
rect 14924 17818 14976 17824
rect 15028 17678 15056 18566
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14844 17338 14872 17614
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 16182 14780 16526
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 15028 15570 15056 17614
rect 15120 17610 15148 19230
rect 15566 19136 15622 19145
rect 15566 19071 15622 19080
rect 15200 18896 15252 18902
rect 15198 18864 15200 18873
rect 15252 18864 15254 18873
rect 15198 18799 15254 18808
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15120 16658 15148 17546
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15580 16114 15608 19071
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17134 15700 17478
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15764 16250 15792 16594
rect 15856 16590 15884 19654
rect 15948 19378 15976 19654
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15946 19068 16254 19077
rect 15946 19066 15952 19068
rect 16008 19066 16032 19068
rect 16088 19066 16112 19068
rect 16168 19066 16192 19068
rect 16248 19066 16254 19068
rect 16008 19014 16010 19066
rect 16190 19014 16192 19066
rect 15946 19012 15952 19014
rect 16008 19012 16032 19014
rect 16088 19012 16112 19014
rect 16168 19012 16192 19014
rect 16248 19012 16254 19014
rect 15946 19003 16254 19012
rect 16316 18426 16344 20946
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 20398 16620 20742
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16868 20058 16896 20946
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16500 19514 16528 19858
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16500 19417 16528 19450
rect 16486 19408 16542 19417
rect 16486 19343 16542 19352
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16684 18358 16712 19994
rect 16960 19990 16988 20742
rect 17144 20466 17172 21247
rect 17960 21072 18012 21078
rect 17960 21014 18012 21020
rect 17972 20602 18000 21014
rect 18248 20942 18276 21422
rect 19064 21412 19116 21418
rect 19064 21354 19116 21360
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17316 20392 17368 20398
rect 17314 20360 17316 20369
rect 17368 20360 17370 20369
rect 17314 20295 17370 20304
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 15946 17980 16254 17989
rect 15946 17978 15952 17980
rect 16008 17978 16032 17980
rect 16088 17978 16112 17980
rect 16168 17978 16192 17980
rect 16248 17978 16254 17980
rect 16008 17926 16010 17978
rect 16190 17926 16192 17978
rect 15946 17924 15952 17926
rect 16008 17924 16032 17926
rect 16088 17924 16112 17926
rect 16168 17924 16192 17926
rect 16248 17924 16254 17926
rect 15946 17915 16254 17924
rect 16578 17912 16634 17921
rect 16578 17847 16634 17856
rect 17040 17876 17092 17882
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 15946 16892 16254 16901
rect 15946 16890 15952 16892
rect 16008 16890 16032 16892
rect 16088 16890 16112 16892
rect 16168 16890 16192 16892
rect 16248 16890 16254 16892
rect 16008 16838 16010 16890
rect 16190 16838 16192 16890
rect 15946 16836 15952 16838
rect 16008 16836 16032 16838
rect 16088 16836 16112 16838
rect 16168 16836 16192 16838
rect 16248 16836 16254 16838
rect 15946 16827 16254 16836
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15856 16130 15884 16526
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15764 16102 15884 16130
rect 15108 16040 15160 16046
rect 15106 16008 15108 16017
rect 15292 16040 15344 16046
rect 15160 16008 15162 16017
rect 15292 15982 15344 15988
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15106 15943 15162 15952
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15212 15162 15240 15370
rect 15304 15162 15332 15982
rect 15488 15706 15516 15982
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15396 15026 15424 15302
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 15108 14952 15160 14958
rect 15488 14906 15516 15506
rect 15108 14894 15160 14900
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14016 13530 14044 14418
rect 14200 14074 14228 14418
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14660 13870 14688 14282
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14660 13462 14688 13806
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14752 12442 14780 14826
rect 14844 14414 14872 14894
rect 15120 14618 15148 14894
rect 15212 14878 15516 14906
rect 15212 14822 15240 14878
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10606 11100 11086
rect 10692 10600 10744 10606
rect 10520 10548 10692 10554
rect 10520 10542 10744 10548
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10520 10526 10732 10542
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8172 10364 8480 10373
rect 8172 10362 8178 10364
rect 8234 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8480 10364
rect 8234 10310 8236 10362
rect 8416 10310 8418 10362
rect 8172 10308 8178 10310
rect 8234 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8480 10310
rect 8172 10299 8480 10308
rect 8588 10266 8616 10406
rect 10428 10266 10456 10474
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10520 10130 10548 10526
rect 11164 10266 11192 11154
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10810 11468 11086
rect 12059 10908 12367 10917
rect 12059 10906 12065 10908
rect 12121 10906 12145 10908
rect 12201 10906 12225 10908
rect 12281 10906 12305 10908
rect 12361 10906 12367 10908
rect 12121 10854 12123 10906
rect 12303 10854 12305 10906
rect 12059 10852 12065 10854
rect 12121 10852 12145 10854
rect 12201 10852 12225 10854
rect 12281 10852 12305 10854
rect 12361 10852 12367 10854
rect 12059 10843 12367 10852
rect 12452 10810 12480 11222
rect 13464 11014 13492 11494
rect 13648 11286 13676 11766
rect 13740 11626 13768 12242
rect 14660 11898 14688 12242
rect 15028 11898 15056 13330
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15028 11694 15056 11834
rect 15212 11830 15240 12242
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 11286 13768 11562
rect 13832 11354 13860 11630
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 4285 9820 4593 9829
rect 4285 9818 4291 9820
rect 4347 9818 4371 9820
rect 4427 9818 4451 9820
rect 4507 9818 4531 9820
rect 4587 9818 4593 9820
rect 4347 9766 4349 9818
rect 4529 9766 4531 9818
rect 4285 9764 4291 9766
rect 4347 9764 4371 9766
rect 4427 9764 4451 9766
rect 4507 9764 4531 9766
rect 4587 9764 4593 9766
rect 4285 9755 4593 9764
rect 11532 9722 11560 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11992 9586 12020 10610
rect 13188 10538 13216 10950
rect 13464 10606 13492 10950
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13464 10198 13492 10542
rect 13648 10470 13676 11222
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 12059 9820 12367 9829
rect 12059 9818 12065 9820
rect 12121 9818 12145 9820
rect 12201 9818 12225 9820
rect 12281 9818 12305 9820
rect 12361 9818 12367 9820
rect 12121 9766 12123 9818
rect 12303 9766 12305 9818
rect 12059 9764 12065 9766
rect 12121 9764 12145 9766
rect 12201 9764 12225 9766
rect 12281 9764 12305 9766
rect 12361 9764 12367 9766
rect 12059 9755 12367 9764
rect 12544 9654 12572 10134
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 13464 9586 13492 10134
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13648 9518 13676 10406
rect 13740 10266 13768 11086
rect 13832 10538 13860 11290
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14016 10606 14044 10950
rect 14108 10810 14136 10950
rect 14844 10810 14872 11222
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 15212 10554 15240 11766
rect 15488 11762 15516 14282
rect 15580 13530 15608 15846
rect 15764 15502 15792 16102
rect 16316 16046 16344 16934
rect 16408 16590 16436 17070
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 15946 15804 16254 15813
rect 15946 15802 15952 15804
rect 16008 15802 16032 15804
rect 16088 15802 16112 15804
rect 16168 15802 16192 15804
rect 16248 15802 16254 15804
rect 16008 15750 16010 15802
rect 16190 15750 16192 15802
rect 15946 15748 15952 15750
rect 16008 15748 16032 15750
rect 16088 15748 16112 15750
rect 16168 15748 16192 15750
rect 16248 15748 16254 15750
rect 15946 15739 16254 15748
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15672 11218 15700 14826
rect 15764 14346 15792 15438
rect 16316 14958 16344 15438
rect 16304 14952 16356 14958
rect 15856 14890 15976 14906
rect 16304 14894 16356 14900
rect 15856 14884 15988 14890
rect 15856 14878 15936 14884
rect 15856 14550 15884 14878
rect 15936 14826 15988 14832
rect 15946 14716 16254 14725
rect 15946 14714 15952 14716
rect 16008 14714 16032 14716
rect 16088 14714 16112 14716
rect 16168 14714 16192 14716
rect 16248 14714 16254 14716
rect 16008 14662 16010 14714
rect 16190 14662 16192 14714
rect 15946 14660 15952 14662
rect 16008 14660 16032 14662
rect 16088 14660 16112 14662
rect 16168 14660 16192 14662
rect 16248 14660 16254 14662
rect 15946 14651 16254 14660
rect 15844 14544 15896 14550
rect 16316 14498 16344 14894
rect 15844 14486 15896 14492
rect 16224 14482 16344 14498
rect 16212 14476 16344 14482
rect 16264 14470 16344 14476
rect 16212 14418 16264 14424
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15946 13628 16254 13637
rect 15946 13626 15952 13628
rect 16008 13626 16032 13628
rect 16088 13626 16112 13628
rect 16168 13626 16192 13628
rect 16248 13626 16254 13628
rect 16008 13574 16010 13626
rect 16190 13574 16192 13626
rect 15946 13572 15952 13574
rect 16008 13572 16032 13574
rect 16088 13572 16112 13574
rect 16168 13572 16192 13574
rect 16248 13572 16254 13574
rect 15946 13563 16254 13572
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 11626 15884 12718
rect 15946 12540 16254 12549
rect 15946 12538 15952 12540
rect 16008 12538 16032 12540
rect 16088 12538 16112 12540
rect 16168 12538 16192 12540
rect 16248 12538 16254 12540
rect 16008 12486 16010 12538
rect 16190 12486 16192 12538
rect 15946 12484 15952 12486
rect 16008 12484 16032 12486
rect 16088 12484 16112 12486
rect 16168 12484 16192 12486
rect 16248 12484 16254 12486
rect 15946 12475 16254 12484
rect 16408 12442 16436 15982
rect 16500 15162 16528 17206
rect 16592 17202 16620 17847
rect 17040 17818 17092 17824
rect 17052 17746 17080 17818
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 17144 17134 17172 19110
rect 17328 18154 17356 20295
rect 17972 20233 18000 20402
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17958 20224 18014 20233
rect 17958 20159 18014 20168
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17512 19854 17540 19994
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17328 17202 17356 18090
rect 17512 17882 17540 19790
rect 17604 19514 17632 19790
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17696 19310 17724 19926
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17604 17814 17632 18566
rect 17696 18426 17724 19246
rect 17788 18970 17816 19314
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 17972 18970 18000 19178
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 18064 17218 18092 20334
rect 18156 19174 18184 20742
rect 18248 20058 18276 20878
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18236 19372 18288 19378
rect 18340 19360 18368 20946
rect 18708 20262 18736 21286
rect 19076 21146 19104 21354
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 20444 21072 20496 21078
rect 20496 21020 20760 21026
rect 20444 21014 20760 21020
rect 19248 21004 19300 21010
rect 20456 20998 20760 21014
rect 19248 20946 19300 20952
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18984 20330 19012 20538
rect 19064 20392 19116 20398
rect 19116 20352 19196 20380
rect 19064 20334 19116 20340
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 18696 20256 18748 20262
rect 19168 20233 19196 20352
rect 18696 20198 18748 20204
rect 19154 20224 19210 20233
rect 19154 20159 19210 20168
rect 19260 19922 19288 20946
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 19833 20700 20141 20709
rect 19833 20698 19839 20700
rect 19895 20698 19919 20700
rect 19975 20698 19999 20700
rect 20055 20698 20079 20700
rect 20135 20698 20141 20700
rect 19895 20646 19897 20698
rect 20077 20646 20079 20698
rect 19833 20644 19839 20646
rect 19895 20644 19919 20646
rect 19975 20644 19999 20646
rect 20055 20644 20079 20646
rect 20135 20644 20141 20646
rect 19833 20635 20141 20644
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 20168 20392 20220 20398
rect 20258 20360 20314 20369
rect 20220 20340 20258 20346
rect 20168 20334 20258 20340
rect 19352 20058 19380 20334
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19064 19440 19116 19446
rect 19064 19382 19116 19388
rect 18288 19332 18368 19360
rect 18236 19314 18288 19320
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18248 18834 18276 19314
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18340 18970 18368 19178
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18524 18834 18552 19246
rect 19076 19156 19104 19382
rect 19168 19310 19196 19858
rect 19260 19514 19288 19858
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19156 19168 19208 19174
rect 19076 19128 19156 19156
rect 19156 19110 19208 19116
rect 19168 18834 19196 19110
rect 19536 18873 19564 20334
rect 20180 20318 20258 20334
rect 20258 20295 20314 20304
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 19996 20097 20024 20198
rect 19982 20088 20038 20097
rect 19982 20023 20038 20032
rect 20088 19961 20116 20198
rect 20074 19952 20130 19961
rect 20074 19887 20130 19896
rect 20076 19712 20128 19718
rect 20128 19672 20208 19700
rect 20076 19654 20128 19660
rect 19833 19612 20141 19621
rect 19833 19610 19839 19612
rect 19895 19610 19919 19612
rect 19975 19610 19999 19612
rect 20055 19610 20079 19612
rect 20135 19610 20141 19612
rect 19895 19558 19897 19610
rect 20077 19558 20079 19610
rect 19833 19556 19839 19558
rect 19895 19556 19919 19558
rect 19975 19556 19999 19558
rect 20055 19556 20079 19558
rect 20135 19556 20141 19558
rect 19833 19547 20141 19556
rect 20180 19514 20208 19672
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 19708 19304 19760 19310
rect 19628 19264 19708 19292
rect 19522 18864 19578 18873
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 19432 18828 19484 18834
rect 19522 18799 19578 18808
rect 19432 18770 19484 18776
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18236 18352 18288 18358
rect 18236 18294 18288 18300
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 17316 17196 17368 17202
rect 17684 17196 17736 17202
rect 17316 17138 17368 17144
rect 17604 17156 17684 17184
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 16046 16620 16390
rect 16776 16250 16804 16662
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17052 15502 17080 15982
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 17052 14958 17080 15438
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17144 14074 17172 15846
rect 17328 14890 17356 17138
rect 17604 16590 17632 17156
rect 17684 17138 17736 17144
rect 17972 17190 18092 17218
rect 17972 17082 18000 17190
rect 17880 17054 18000 17082
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17880 16810 17908 17054
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17696 16794 17908 16810
rect 17684 16788 17908 16794
rect 17736 16782 17908 16788
rect 17684 16730 17736 16736
rect 17972 16658 18000 16934
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 18064 16250 18092 17070
rect 18156 16969 18184 17274
rect 18248 17270 18276 18294
rect 18696 18148 18748 18154
rect 18696 18090 18748 18096
rect 18708 17882 18736 18090
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18524 17542 18552 17614
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18340 17377 18368 17478
rect 18326 17368 18382 17377
rect 18326 17303 18382 17312
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18142 16960 18198 16969
rect 18142 16895 18198 16904
rect 18142 16688 18198 16697
rect 18248 16658 18276 17206
rect 18524 17134 18552 17478
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18142 16623 18144 16632
rect 18196 16623 18198 16632
rect 18236 16652 18288 16658
rect 18144 16594 18196 16600
rect 18236 16594 18288 16600
rect 18616 16590 18644 17818
rect 18892 17746 18920 18566
rect 18984 18426 19012 18770
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18972 18080 19024 18086
rect 19076 18034 19104 18566
rect 19024 18028 19104 18034
rect 18972 18022 19104 18028
rect 18984 18006 19104 18022
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18970 17096 19026 17105
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18786 16960 18842 16969
rect 18604 16584 18656 16590
rect 18510 16552 18566 16561
rect 18604 16526 18656 16532
rect 18510 16487 18566 16496
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18248 16114 18276 16390
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18340 16046 18368 16186
rect 17500 16040 17552 16046
rect 17498 16008 17500 16017
rect 18144 16040 18196 16046
rect 17552 16008 17554 16017
rect 18144 15982 18196 15988
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 17498 15943 17554 15952
rect 17512 14958 17540 15943
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15026 17632 15846
rect 18156 15570 18184 15982
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 17788 15162 17816 15506
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17420 14618 17448 14826
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17604 13870 17632 14350
rect 18340 14074 18368 15846
rect 18432 14958 18460 15846
rect 18524 15706 18552 16487
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18708 14958 18736 16934
rect 18786 16895 18842 16904
rect 18800 16726 18828 16895
rect 18892 16794 18920 17070
rect 18970 17031 18972 17040
rect 19024 17031 19026 17040
rect 18972 17002 19024 17008
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18432 14278 18460 14894
rect 18800 14414 18828 15438
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17604 13394 17632 13806
rect 18432 13802 18460 14214
rect 17684 13796 17736 13802
rect 17684 13738 17736 13744
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17696 12918 17724 13738
rect 18892 13530 18920 14894
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16868 12442 16896 12650
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16856 12436 16908 12442
rect 17696 12434 17724 12854
rect 17972 12646 18000 13398
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 16856 12378 16908 12384
rect 17604 12406 17724 12434
rect 17776 12436 17828 12442
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11354 15792 11494
rect 15946 11452 16254 11461
rect 15946 11450 15952 11452
rect 16008 11450 16032 11452
rect 16088 11450 16112 11452
rect 16168 11450 16192 11452
rect 16248 11450 16254 11452
rect 16008 11398 16010 11450
rect 16190 11398 16192 11450
rect 15946 11396 15952 11398
rect 16008 11396 16032 11398
rect 16088 11396 16112 11398
rect 16168 11396 16192 11398
rect 16248 11396 16254 11398
rect 15946 11387 16254 11396
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 16408 10674 16436 11630
rect 16868 11354 16896 12038
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 17052 11354 17080 11562
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 13820 10532 13872 10538
rect 15212 10526 15332 10554
rect 13820 10474 13872 10480
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 15212 10130 15240 10406
rect 15304 10266 15332 10526
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 15946 10364 16254 10373
rect 15946 10362 15952 10364
rect 16008 10362 16032 10364
rect 16088 10362 16112 10364
rect 16168 10362 16192 10364
rect 16248 10362 16254 10364
rect 16008 10310 16010 10362
rect 16190 10310 16192 10362
rect 15946 10308 15952 10310
rect 16008 10308 16032 10310
rect 16088 10308 16112 10310
rect 16168 10308 16192 10310
rect 16248 10308 16254 10310
rect 15946 10299 16254 10308
rect 16684 10266 16712 10474
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16868 10198 16896 11290
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 17236 10062 17264 12242
rect 17604 12238 17632 12406
rect 17776 12378 17828 12384
rect 17788 12322 17816 12378
rect 17696 12294 17816 12322
rect 17880 12306 17908 12582
rect 17972 12306 18000 12582
rect 18340 12442 18368 12718
rect 18984 12714 19012 15506
rect 19076 13462 19104 18006
rect 19168 14482 19196 18770
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19260 18426 19288 18702
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19338 18320 19394 18329
rect 19338 18255 19340 18264
rect 19392 18255 19394 18264
rect 19340 18226 19392 18232
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19260 17746 19288 18158
rect 19444 18086 19472 18770
rect 19522 18728 19578 18737
rect 19522 18663 19524 18672
rect 19576 18663 19578 18672
rect 19524 18634 19576 18640
rect 19522 18184 19578 18193
rect 19522 18119 19578 18128
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19246 17368 19302 17377
rect 19246 17303 19302 17312
rect 19260 17134 19288 17303
rect 19444 17134 19472 18022
rect 19536 17610 19564 18119
rect 19628 17746 19656 19264
rect 19708 19246 19760 19252
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19904 19174 19932 19246
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 20088 18902 20116 19450
rect 20272 19310 20300 20198
rect 20364 19904 20392 20878
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 20398 20576 20742
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20640 20262 20668 20538
rect 20732 20398 20760 20998
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20824 20602 20852 20878
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20456 20058 20484 20198
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20444 19916 20496 19922
rect 20364 19876 20444 19904
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20260 19304 20312 19310
rect 20364 19281 20392 19876
rect 20444 19858 20496 19864
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20260 19246 20312 19252
rect 20350 19272 20406 19281
rect 20180 19174 20208 19246
rect 20168 19168 20220 19174
rect 20272 19156 20300 19246
rect 20456 19224 20484 19722
rect 20350 19207 20406 19216
rect 20444 19196 20484 19224
rect 20444 19156 20472 19196
rect 20272 19128 20392 19156
rect 20444 19128 20484 19156
rect 20168 19110 20220 19116
rect 20076 18896 20128 18902
rect 20076 18838 20128 18844
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19812 18612 19840 18770
rect 19904 18630 19932 18770
rect 19720 18584 19840 18612
rect 19892 18624 19944 18630
rect 19720 18426 19748 18584
rect 19892 18566 19944 18572
rect 19833 18524 20141 18533
rect 19833 18522 19839 18524
rect 19895 18522 19919 18524
rect 19975 18522 19999 18524
rect 20055 18522 20079 18524
rect 20135 18522 20141 18524
rect 19895 18470 19897 18522
rect 20077 18470 20079 18522
rect 19833 18468 19839 18470
rect 19895 18468 19919 18470
rect 19975 18468 19999 18470
rect 20055 18468 20079 18470
rect 20135 18468 20141 18470
rect 19833 18459 20141 18468
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19720 17882 19748 18158
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19524 17604 19576 17610
rect 19524 17546 19576 17552
rect 19833 17436 20141 17445
rect 19833 17434 19839 17436
rect 19895 17434 19919 17436
rect 19975 17434 19999 17436
rect 20055 17434 20079 17436
rect 20135 17434 20141 17436
rect 19895 17382 19897 17434
rect 20077 17382 20079 17434
rect 19833 17380 19839 17382
rect 19895 17380 19919 17382
rect 19975 17380 19999 17382
rect 20055 17380 20079 17382
rect 20135 17380 20141 17382
rect 19833 17371 20141 17380
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16726 19380 16934
rect 19536 16794 19564 17274
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19833 16348 20141 16357
rect 19833 16346 19839 16348
rect 19895 16346 19919 16348
rect 19975 16346 19999 16348
rect 20055 16346 20079 16348
rect 20135 16346 20141 16348
rect 19895 16294 19897 16346
rect 20077 16294 20079 16346
rect 19833 16292 19839 16294
rect 19895 16292 19919 16294
rect 19975 16292 19999 16294
rect 20055 16292 20079 16294
rect 20135 16292 20141 16294
rect 19833 16283 20141 16292
rect 20076 16040 20128 16046
rect 20074 16008 20076 16017
rect 20128 16008 20130 16017
rect 20074 15943 20130 15952
rect 19833 15260 20141 15269
rect 19833 15258 19839 15260
rect 19895 15258 19919 15260
rect 19975 15258 19999 15260
rect 20055 15258 20079 15260
rect 20135 15258 20141 15260
rect 19895 15206 19897 15258
rect 20077 15206 20079 15258
rect 19833 15204 19839 15206
rect 19895 15204 19919 15206
rect 19975 15204 19999 15206
rect 20055 15204 20079 15206
rect 20135 15204 20141 15206
rect 19833 15195 20141 15204
rect 20180 14958 20208 19110
rect 20260 18352 20312 18358
rect 20258 18320 20260 18329
rect 20312 18320 20314 18329
rect 20258 18255 20314 18264
rect 20260 18216 20312 18222
rect 20364 18204 20392 19128
rect 20312 18176 20392 18204
rect 20260 18158 20312 18164
rect 20272 17746 20300 18158
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20456 17610 20484 19128
rect 20548 18873 20576 19926
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19258 20668 19654
rect 20824 19446 20852 19790
rect 20916 19514 20944 19858
rect 21008 19854 21036 21422
rect 21468 21146 21496 21422
rect 22192 21412 22244 21418
rect 22192 21354 22244 21360
rect 22204 21146 22232 21354
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 21088 20392 21140 20398
rect 21086 20360 21088 20369
rect 21140 20360 21142 20369
rect 21086 20295 21142 20304
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21008 19514 21036 19790
rect 21192 19786 21220 21082
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21468 20466 21496 20742
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21824 20392 21876 20398
rect 21824 20334 21876 20340
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20904 19304 20956 19310
rect 20640 19230 20852 19258
rect 20904 19246 20956 19252
rect 20994 19272 21050 19281
rect 20534 18864 20590 18873
rect 20824 18816 20852 19230
rect 20534 18799 20590 18808
rect 20548 18222 20576 18799
rect 20732 18788 20852 18816
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20272 17270 20300 17546
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19720 13530 19748 14826
rect 20272 14226 20300 16050
rect 20364 15026 20392 17070
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 15978 20484 16390
rect 20548 16250 20576 18158
rect 20732 17746 20760 18788
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20824 18358 20852 18634
rect 20916 18630 20944 19246
rect 20994 19207 21050 19216
rect 21008 18834 21036 19207
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20916 18222 20944 18566
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20824 16250 20852 18158
rect 21008 17134 21036 18566
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21100 17134 21128 17478
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 21008 16590 21036 16662
rect 21652 16658 21680 16934
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20916 15706 20944 15914
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20364 14822 20392 14962
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20732 14618 20760 15302
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20628 14272 20680 14278
rect 20272 14198 20576 14226
rect 20628 14214 20680 14220
rect 19833 14172 20141 14181
rect 19833 14170 19839 14172
rect 19895 14170 19919 14172
rect 19975 14170 19999 14172
rect 20055 14170 20079 14172
rect 20135 14170 20141 14172
rect 19895 14118 19897 14170
rect 20077 14118 20079 14170
rect 19833 14116 19839 14118
rect 19895 14116 19919 14118
rect 19975 14116 19999 14118
rect 20055 14116 20079 14118
rect 20135 14116 20141 14118
rect 19833 14107 20141 14116
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18432 12322 18460 12582
rect 18340 12306 18460 12322
rect 17868 12300 17920 12306
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17328 11558 17356 12106
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17696 11354 17724 12294
rect 17868 12242 17920 12248
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18328 12300 18460 12306
rect 18380 12294 18460 12300
rect 18328 12242 18380 12248
rect 17880 12186 17908 12242
rect 17788 12158 17908 12186
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 17788 11898 17816 12158
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17788 11234 17816 11834
rect 17960 11280 18012 11286
rect 17788 11228 17960 11234
rect 17788 11222 18012 11228
rect 17788 11206 18000 11222
rect 18064 11218 18092 12174
rect 18708 11898 18736 12174
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 19076 11694 19104 13398
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12986 19472 13262
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 19833 13084 20141 13093
rect 19833 13082 19839 13084
rect 19895 13082 19919 13084
rect 19975 13082 19999 13084
rect 20055 13082 20079 13084
rect 20135 13082 20141 13084
rect 19895 13030 19897 13082
rect 20077 13030 20079 13082
rect 19833 13028 19839 13030
rect 19895 13028 19919 13030
rect 19975 13028 19999 13030
rect 20055 13028 20079 13030
rect 20135 13028 20141 13030
rect 19833 13019 20141 13028
rect 20180 12986 20208 13126
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20364 12714 20392 13194
rect 20352 12708 20404 12714
rect 20352 12650 20404 12656
rect 19833 11996 20141 12005
rect 19833 11994 19839 11996
rect 19895 11994 19919 11996
rect 19975 11994 19999 11996
rect 20055 11994 20079 11996
rect 20135 11994 20141 11996
rect 19895 11942 19897 11994
rect 20077 11942 20079 11994
rect 19833 11940 19839 11942
rect 19895 11940 19919 11942
rect 19975 11940 19999 11942
rect 20055 11940 20079 11942
rect 20135 11940 20141 11942
rect 19833 11931 20141 11940
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18064 10470 18092 11154
rect 18708 10538 18736 11494
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19444 10674 19472 10950
rect 19833 10908 20141 10917
rect 19833 10906 19839 10908
rect 19895 10906 19919 10908
rect 19975 10906 19999 10908
rect 20055 10906 20079 10908
rect 20135 10906 20141 10908
rect 19895 10854 19897 10906
rect 20077 10854 20079 10906
rect 19833 10852 19839 10854
rect 19895 10852 19919 10854
rect 19975 10852 19999 10854
rect 20055 10852 20079 10854
rect 20135 10852 20141 10854
rect 19833 10843 20141 10852
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 19800 10532 19852 10538
rect 19800 10474 19852 10480
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17696 10130 17724 10406
rect 18708 10130 18736 10474
rect 19812 10266 19840 10474
rect 20364 10470 20392 12650
rect 20548 12442 20576 14198
rect 20640 14074 20668 14214
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 21008 13870 21036 16526
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 14482 21312 15846
rect 21376 15570 21404 16118
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21468 15706 21496 15982
rect 21560 15910 21588 16594
rect 21836 16114 21864 20334
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22112 19514 22140 19858
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 22112 17066 22140 18158
rect 22296 17134 22324 19110
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22100 17060 22152 17066
rect 22100 17002 22152 17008
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 22008 15972 22060 15978
rect 22112 15960 22140 16526
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22060 15932 22140 15960
rect 22008 15914 22060 15920
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 22112 15638 22140 15932
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 22204 15366 22232 16390
rect 22388 16250 22416 20334
rect 22480 16998 22508 20334
rect 22664 20210 22692 21286
rect 22756 20398 22784 21286
rect 23032 21010 23060 21558
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 23720 21244 24028 21253
rect 23720 21242 23726 21244
rect 23782 21242 23806 21244
rect 23862 21242 23886 21244
rect 23942 21242 23966 21244
rect 24022 21242 24028 21244
rect 23782 21190 23784 21242
rect 23964 21190 23966 21242
rect 23720 21188 23726 21190
rect 23782 21188 23806 21190
rect 23862 21188 23886 21190
rect 23942 21188 23966 21190
rect 24022 21188 24028 21190
rect 23720 21179 24028 21188
rect 24596 21146 24624 21286
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 23020 21004 23072 21010
rect 23020 20946 23072 20952
rect 24688 20874 24716 21286
rect 24872 21146 24900 21354
rect 25240 21146 25268 21422
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 25228 21140 25280 21146
rect 25228 21082 25280 21088
rect 25424 21010 25452 21558
rect 25884 21486 25912 21791
rect 26804 21486 26832 21791
rect 27607 21788 27915 21797
rect 28538 21791 28594 21800
rect 27607 21786 27613 21788
rect 27669 21786 27693 21788
rect 27749 21786 27773 21788
rect 27829 21786 27853 21788
rect 27909 21786 27915 21788
rect 27669 21734 27671 21786
rect 27851 21734 27853 21786
rect 27607 21732 27613 21734
rect 27669 21732 27693 21734
rect 27749 21732 27773 21734
rect 27829 21732 27853 21734
rect 27909 21732 27915 21734
rect 27607 21723 27915 21732
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 26884 21548 26936 21554
rect 26884 21490 26936 21496
rect 25872 21480 25924 21486
rect 25872 21422 25924 21428
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 25516 21146 25544 21286
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25412 21004 25464 21010
rect 25412 20946 25464 20952
rect 25516 20874 25544 21082
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 25504 20868 25556 20874
rect 25504 20810 25556 20816
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 23112 20392 23164 20398
rect 23112 20334 23164 20340
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22848 20233 22876 20266
rect 22834 20224 22890 20233
rect 22664 20182 22784 20210
rect 22756 19854 22784 20182
rect 22834 20159 22890 20168
rect 22940 20058 22968 20334
rect 22928 20052 22980 20058
rect 22928 19994 22980 20000
rect 23124 19990 23152 20334
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22652 18760 22704 18766
rect 22756 18748 22784 19790
rect 23020 19236 23072 19242
rect 23020 19178 23072 19184
rect 23032 18970 23060 19178
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 22704 18720 22784 18748
rect 22652 18702 22704 18708
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22572 18222 22600 18634
rect 22652 18352 22704 18358
rect 22650 18320 22652 18329
rect 22704 18320 22706 18329
rect 22650 18255 22706 18264
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22756 18170 22784 18720
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 23032 18222 23060 18634
rect 23216 18290 23244 18634
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23020 18216 23072 18222
rect 22664 17542 22692 18158
rect 22756 18142 22968 18170
rect 23020 18158 23072 18164
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22480 16794 22508 16934
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22572 16726 22600 17070
rect 22848 16726 22876 17818
rect 22940 17746 22968 18142
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23216 17814 23244 18022
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22836 16720 22888 16726
rect 22836 16662 22888 16668
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22480 16250 22508 16594
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22468 16040 22520 16046
rect 22374 16008 22430 16017
rect 22284 15972 22336 15978
rect 22468 15982 22520 15988
rect 22374 15943 22430 15952
rect 22284 15914 22336 15920
rect 22296 15706 22324 15914
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22388 15638 22416 15943
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22100 14884 22152 14890
rect 22100 14826 22152 14832
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 21744 14618 21772 14758
rect 22020 14618 22048 14758
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21744 14074 21772 14214
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 22112 13938 22140 14826
rect 22204 14482 22232 14894
rect 22296 14618 22324 15506
rect 22480 15366 22508 15982
rect 22572 15570 22600 16390
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 14958 22508 15302
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22284 14612 22336 14618
rect 22664 14600 22692 16186
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22284 14554 22336 14560
rect 22572 14572 22692 14600
rect 22572 14482 22600 14572
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22100 13932 22152 13938
rect 22020 13892 22100 13920
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20640 11898 20668 13806
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12782 21404 13126
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 22020 12306 22048 13892
rect 22100 13874 22152 13880
rect 22572 13802 22600 14418
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22112 13326 22140 13738
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22112 12986 22140 13262
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22572 12374 22600 12582
rect 22664 12442 22692 14418
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 21560 11694 21588 12242
rect 21640 12096 21692 12102
rect 21916 12096 21968 12102
rect 21692 12044 21864 12050
rect 21640 12038 21864 12044
rect 21916 12038 21968 12044
rect 21652 12022 21864 12038
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21836 11626 21864 12022
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 11218 20668 11494
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20640 10810 20668 11154
rect 20824 11014 20852 11562
rect 20996 11552 21048 11558
rect 20994 11520 20996 11529
rect 21088 11552 21140 11558
rect 21048 11520 21050 11529
rect 21744 11529 21772 11562
rect 21088 11494 21140 11500
rect 21730 11520 21786 11529
rect 20994 11455 21050 11464
rect 21100 11354 21128 11494
rect 21730 11455 21786 11464
rect 21744 11354 21772 11455
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21548 11348 21600 11354
rect 21732 11348 21784 11354
rect 21548 11290 21600 11296
rect 21652 11308 21732 11336
rect 21560 11150 21588 11290
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 21192 10266 21220 10610
rect 21560 10606 21588 11086
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 13924 9722 13952 9998
rect 21652 9926 21680 11308
rect 21732 11290 21784 11296
rect 21928 11218 21956 12038
rect 22756 11558 22784 12582
rect 22848 11898 22876 15982
rect 22940 14958 22968 16934
rect 23124 16794 23152 16934
rect 23216 16794 23244 17274
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23308 16658 23336 19858
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23296 16652 23348 16658
rect 23296 16594 23348 16600
rect 23216 16561 23244 16594
rect 23202 16552 23258 16561
rect 23202 16487 23258 16496
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23032 15366 23060 15982
rect 23400 15978 23428 20266
rect 23720 20156 24028 20165
rect 23720 20154 23726 20156
rect 23782 20154 23806 20156
rect 23862 20154 23886 20156
rect 23942 20154 23966 20156
rect 24022 20154 24028 20156
rect 23782 20102 23784 20154
rect 23964 20102 23966 20154
rect 23720 20100 23726 20102
rect 23782 20100 23806 20102
rect 23862 20100 23886 20102
rect 23942 20100 23966 20102
rect 24022 20100 24028 20102
rect 23720 20091 24028 20100
rect 24412 20058 24440 20742
rect 24492 20528 24544 20534
rect 24490 20496 24492 20505
rect 24676 20528 24728 20534
rect 24544 20496 24546 20505
rect 24676 20470 24728 20476
rect 24490 20431 24546 20440
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 24400 20052 24452 20058
rect 24400 19994 24452 20000
rect 24308 19916 24360 19922
rect 24308 19858 24360 19864
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 23676 19514 23704 19654
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23754 19408 23810 19417
rect 23754 19343 23810 19352
rect 23768 19310 23796 19343
rect 24136 19310 24164 19654
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 23720 19068 24028 19077
rect 23720 19066 23726 19068
rect 23782 19066 23806 19068
rect 23862 19066 23886 19068
rect 23942 19066 23966 19068
rect 24022 19066 24028 19068
rect 23782 19014 23784 19066
rect 23964 19014 23966 19066
rect 23720 19012 23726 19014
rect 23782 19012 23806 19014
rect 23862 19012 23886 19014
rect 23942 19012 23966 19014
rect 24022 19012 24028 19014
rect 23720 19003 24028 19012
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23492 16153 23520 18906
rect 23572 18760 23624 18766
rect 23570 18728 23572 18737
rect 23624 18728 23626 18737
rect 23570 18663 23626 18672
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23570 18320 23626 18329
rect 23860 18290 23888 18634
rect 23570 18255 23626 18264
rect 23848 18284 23900 18290
rect 23584 18222 23612 18255
rect 23848 18226 23900 18232
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23584 17542 23612 18022
rect 23720 17980 24028 17989
rect 23720 17978 23726 17980
rect 23782 17978 23806 17980
rect 23862 17978 23886 17980
rect 23942 17978 23966 17980
rect 24022 17978 24028 17980
rect 23782 17926 23784 17978
rect 23964 17926 23966 17978
rect 23720 17924 23726 17926
rect 23782 17924 23806 17926
rect 23862 17924 23886 17926
rect 23942 17924 23966 17926
rect 24022 17924 24028 17926
rect 23720 17915 24028 17924
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23584 16658 23612 17478
rect 23720 16892 24028 16901
rect 23720 16890 23726 16892
rect 23782 16890 23806 16892
rect 23862 16890 23886 16892
rect 23942 16890 23966 16892
rect 24022 16890 24028 16892
rect 23782 16838 23784 16890
rect 23964 16838 23966 16890
rect 23720 16836 23726 16838
rect 23782 16836 23806 16838
rect 23862 16836 23886 16838
rect 23942 16836 23966 16838
rect 24022 16836 24028 16838
rect 23720 16827 24028 16836
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 24228 16454 24256 19654
rect 24320 19242 24348 19858
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24308 19236 24360 19242
rect 24308 19178 24360 19184
rect 24320 18154 24348 19178
rect 24400 18896 24452 18902
rect 24400 18838 24452 18844
rect 24412 18222 24440 18838
rect 24504 18630 24532 19246
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24400 18216 24452 18222
rect 24504 18193 24532 18566
rect 24400 18158 24452 18164
rect 24490 18184 24546 18193
rect 24308 18148 24360 18154
rect 24308 18090 24360 18096
rect 24412 17626 24440 18158
rect 24490 18119 24546 18128
rect 24412 17598 24532 17626
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 23860 16182 23888 16390
rect 24412 16250 24440 17478
rect 24504 17338 24532 17598
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 23848 16176 23900 16182
rect 23478 16144 23534 16153
rect 23848 16118 23900 16124
rect 24030 16144 24086 16153
rect 23478 16079 23534 16088
rect 24596 16130 24624 20266
rect 24688 19514 24716 20470
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24780 20058 24808 20198
rect 24872 20058 24900 20334
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 25688 20052 25740 20058
rect 25688 19994 25740 20000
rect 24780 19514 24808 19994
rect 24858 19952 24914 19961
rect 24858 19887 24860 19896
rect 24912 19887 24914 19896
rect 24860 19858 24912 19864
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 24964 18970 24992 19246
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24688 18154 24716 18702
rect 24964 18358 24992 18906
rect 25056 18902 25084 19246
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25044 18896 25096 18902
rect 25044 18838 25096 18844
rect 25056 18698 25084 18838
rect 25044 18692 25096 18698
rect 25044 18634 25096 18640
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24964 18222 24992 18294
rect 24952 18216 25004 18222
rect 24872 18176 24952 18204
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24872 17814 24900 18176
rect 24952 18158 25004 18164
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24860 17808 24912 17814
rect 24780 17756 24860 17762
rect 24780 17750 24912 17756
rect 24780 17734 24900 17750
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24688 16658 24716 17206
rect 24780 17066 24808 17734
rect 24964 17678 24992 18022
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24768 17060 24820 17066
rect 24768 17002 24820 17008
rect 24872 16794 24900 17546
rect 24964 16998 24992 17614
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 25240 16658 25268 19110
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25320 16992 25372 16998
rect 25320 16934 25372 16940
rect 25332 16658 25360 16934
rect 25424 16658 25452 18566
rect 25700 16658 25728 19994
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25792 18630 25820 19110
rect 25872 18828 25924 18834
rect 25872 18770 25924 18776
rect 25884 18630 25912 18770
rect 25780 18624 25832 18630
rect 25780 18566 25832 18572
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25884 17814 25912 18566
rect 25872 17808 25924 17814
rect 25872 17750 25924 17756
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 24030 16079 24086 16088
rect 24412 16102 24624 16130
rect 24044 16046 24072 16079
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23020 15360 23072 15366
rect 23020 15302 23072 15308
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23308 14346 23336 14758
rect 23400 14414 23428 15914
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 23720 15804 24028 15813
rect 23720 15802 23726 15804
rect 23782 15802 23806 15804
rect 23862 15802 23886 15804
rect 23942 15802 23966 15804
rect 24022 15802 24028 15804
rect 23782 15750 23784 15802
rect 23964 15750 23966 15802
rect 23720 15748 23726 15750
rect 23782 15748 23806 15750
rect 23862 15748 23886 15750
rect 23942 15748 23966 15750
rect 24022 15748 24028 15750
rect 23720 15739 24028 15748
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23480 14884 23532 14890
rect 23480 14826 23532 14832
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23308 13326 23336 14282
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22940 12646 22968 12922
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 23032 12434 23060 13126
rect 23492 12782 23520 14826
rect 23584 14074 23612 15506
rect 23720 14716 24028 14725
rect 23720 14714 23726 14716
rect 23782 14714 23806 14716
rect 23862 14714 23886 14716
rect 23942 14714 23966 14716
rect 24022 14714 24028 14716
rect 23782 14662 23784 14714
rect 23964 14662 23966 14714
rect 23720 14660 23726 14662
rect 23782 14660 23806 14662
rect 23862 14660 23886 14662
rect 23942 14660 23966 14662
rect 24022 14660 24028 14662
rect 23720 14651 24028 14660
rect 24136 14618 24164 15846
rect 24412 15434 24440 16102
rect 24688 15502 24716 16594
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24400 15428 24452 15434
rect 24400 15370 24452 15376
rect 24492 15360 24544 15366
rect 24492 15302 24544 15308
rect 24504 14958 24532 15302
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 24044 13870 24072 14418
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24320 13870 24348 14214
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 23720 13628 24028 13637
rect 23720 13626 23726 13628
rect 23782 13626 23806 13628
rect 23862 13626 23886 13628
rect 23942 13626 23966 13628
rect 24022 13626 24028 13628
rect 23782 13574 23784 13626
rect 23964 13574 23966 13626
rect 23720 13572 23726 13574
rect 23782 13572 23806 13574
rect 23862 13572 23886 13574
rect 23942 13572 23966 13574
rect 24022 13572 24028 13574
rect 23720 13563 24028 13572
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23676 12782 23704 13126
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 22940 12406 23060 12434
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22940 11762 22968 12406
rect 23492 12186 23520 12718
rect 23720 12540 24028 12549
rect 23720 12538 23726 12540
rect 23782 12538 23806 12540
rect 23862 12538 23886 12540
rect 23942 12538 23966 12540
rect 24022 12538 24028 12540
rect 23782 12486 23784 12538
rect 23964 12486 23966 12538
rect 23720 12484 23726 12486
rect 23782 12484 23806 12486
rect 23862 12484 23886 12486
rect 23942 12484 23966 12486
rect 24022 12484 24028 12486
rect 23720 12475 24028 12484
rect 24320 12306 24348 13806
rect 24400 13728 24452 13734
rect 24400 13670 24452 13676
rect 24412 13326 24440 13670
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24412 12986 24440 13262
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24688 12646 24716 13126
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 23492 12158 23612 12186
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23492 11762 23520 12038
rect 23584 11898 23612 12158
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 22756 11218 22784 11494
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21744 10198 21772 10950
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21928 10062 21956 11154
rect 22940 11150 22968 11698
rect 23720 11452 24028 11461
rect 23720 11450 23726 11452
rect 23782 11450 23806 11452
rect 23862 11450 23886 11452
rect 23942 11450 23966 11452
rect 24022 11450 24028 11452
rect 23782 11398 23784 11450
rect 23964 11398 23966 11450
rect 23720 11396 23726 11398
rect 23782 11396 23806 11398
rect 23862 11396 23886 11398
rect 23942 11396 23966 11398
rect 24022 11396 24028 11398
rect 23720 11387 24028 11396
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 23492 10810 23520 11154
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 24320 10674 24348 12242
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 11898 24624 12174
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24688 11830 24716 12038
rect 24676 11824 24728 11830
rect 24676 11766 24728 11772
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24688 11286 24716 11630
rect 24780 11354 24808 16594
rect 25516 16250 25544 16594
rect 25700 16561 25728 16594
rect 25686 16552 25742 16561
rect 25686 16487 25742 16496
rect 25780 16516 25832 16522
rect 25780 16458 25832 16464
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25792 15638 25820 16458
rect 25872 15904 25924 15910
rect 25872 15846 25924 15852
rect 25884 15638 25912 15846
rect 25976 15638 26004 20742
rect 26068 19922 26096 21286
rect 26160 20058 26188 21286
rect 26424 20868 26476 20874
rect 26608 20868 26660 20874
rect 26476 20828 26608 20856
rect 26424 20810 26476 20816
rect 26608 20810 26660 20816
rect 26436 20398 26464 20810
rect 26896 20398 26924 21490
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26884 20392 26936 20398
rect 26884 20334 26936 20340
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 26068 19378 26096 19858
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 26068 18834 26096 19314
rect 26160 18970 26188 19994
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 26056 18828 26108 18834
rect 26056 18770 26108 18776
rect 26056 18692 26108 18698
rect 26056 18634 26108 18640
rect 26068 17882 26096 18634
rect 26160 18222 26188 18906
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 26160 17542 26188 18158
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 25228 15632 25280 15638
rect 25228 15574 25280 15580
rect 25780 15632 25832 15638
rect 25780 15574 25832 15580
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 25240 15162 25268 15574
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 25884 14958 25912 15574
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24872 12986 24900 14554
rect 25884 14414 25912 14894
rect 26056 14884 26108 14890
rect 26056 14826 26108 14832
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 25976 14414 26004 14554
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 26068 14074 26096 14826
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24964 13394 24992 13670
rect 25056 13394 25084 14010
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25240 13530 25268 13874
rect 25596 13796 25648 13802
rect 25596 13738 25648 13744
rect 25608 13530 25636 13738
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 25148 12646 25176 13466
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25332 12866 25360 13330
rect 26068 13326 26096 14010
rect 26252 13870 26280 20198
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26712 19310 26740 19654
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 27080 19242 27108 20946
rect 27172 20505 27200 21626
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 27252 21412 27304 21418
rect 27252 21354 27304 21360
rect 27264 21010 27292 21354
rect 27252 21004 27304 21010
rect 27252 20946 27304 20952
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 27158 20496 27214 20505
rect 27158 20431 27214 20440
rect 27264 20330 27292 20742
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27172 20058 27200 20198
rect 27160 20052 27212 20058
rect 27160 19994 27212 20000
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 27068 19236 27120 19242
rect 27068 19178 27120 19184
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 26976 19168 27028 19174
rect 26976 19110 27028 19116
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 27264 19122 27292 19450
rect 27356 19310 27384 21558
rect 28552 21486 28580 21791
rect 29012 21486 29040 21927
rect 29368 21888 29420 21894
rect 29368 21830 29420 21836
rect 30010 21856 30066 21865
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 29000 21480 29052 21486
rect 29000 21422 29052 21428
rect 28080 21412 28132 21418
rect 28080 21354 28132 21360
rect 28092 21298 28120 21354
rect 28264 21344 28316 21350
rect 28092 21270 28212 21298
rect 28264 21286 28316 21292
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27988 21004 28040 21010
rect 27988 20946 28040 20952
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 27448 20466 27476 20878
rect 27540 20602 27568 20946
rect 27607 20700 27915 20709
rect 27607 20698 27613 20700
rect 27669 20698 27693 20700
rect 27749 20698 27773 20700
rect 27829 20698 27853 20700
rect 27909 20698 27915 20700
rect 27669 20646 27671 20698
rect 27851 20646 27853 20698
rect 27607 20644 27613 20646
rect 27669 20644 27693 20646
rect 27749 20644 27773 20646
rect 27829 20644 27853 20646
rect 27909 20644 27915 20646
rect 27607 20635 27915 20644
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27526 20496 27582 20505
rect 27436 20460 27488 20466
rect 27582 20454 27660 20482
rect 27526 20431 27582 20440
rect 27436 20402 27488 20408
rect 27632 20398 27660 20454
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27632 20058 27660 20334
rect 28000 20262 28028 20946
rect 28092 20398 28120 20946
rect 28080 20392 28132 20398
rect 28080 20334 28132 20340
rect 27988 20256 28040 20262
rect 27988 20198 28040 20204
rect 27620 20052 27672 20058
rect 27620 19994 27672 20000
rect 27607 19612 27915 19621
rect 27607 19610 27613 19612
rect 27669 19610 27693 19612
rect 27749 19610 27773 19612
rect 27829 19610 27853 19612
rect 27909 19610 27915 19612
rect 27669 19558 27671 19610
rect 27851 19558 27853 19610
rect 27607 19556 27613 19558
rect 27669 19556 27693 19558
rect 27749 19556 27773 19558
rect 27829 19556 27853 19558
rect 27909 19556 27915 19558
rect 27607 19547 27915 19556
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27436 19168 27488 19174
rect 26896 18970 26924 19110
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 26896 18426 26924 18906
rect 26988 18902 27016 19110
rect 26976 18896 27028 18902
rect 26976 18838 27028 18844
rect 26884 18420 26936 18426
rect 26884 18362 26936 18368
rect 27172 18222 27200 19110
rect 27264 19094 27384 19122
rect 27436 19110 27488 19116
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 27264 18426 27292 18566
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27356 18358 27384 19094
rect 27448 18970 27476 19110
rect 27436 18964 27488 18970
rect 27436 18906 27488 18912
rect 27448 18834 27476 18906
rect 27436 18828 27488 18834
rect 27436 18770 27488 18776
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27448 18426 27476 18634
rect 27607 18524 27915 18533
rect 27607 18522 27613 18524
rect 27669 18522 27693 18524
rect 27749 18522 27773 18524
rect 27829 18522 27853 18524
rect 27909 18522 27915 18524
rect 27669 18470 27671 18522
rect 27851 18470 27853 18522
rect 27607 18468 27613 18470
rect 27669 18468 27693 18470
rect 27749 18468 27773 18470
rect 27829 18468 27853 18470
rect 27909 18468 27915 18470
rect 27607 18459 27915 18468
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27344 18352 27396 18358
rect 27344 18294 27396 18300
rect 26424 18216 26476 18222
rect 26424 18158 26476 18164
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 26330 17776 26386 17785
rect 26330 17711 26386 17720
rect 26344 17542 26372 17711
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 17134 26372 17478
rect 26436 17134 26464 18158
rect 26804 17882 26832 18158
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 26620 17338 26648 17614
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26700 17264 26752 17270
rect 26700 17206 26752 17212
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26344 16153 26372 16186
rect 26712 16182 26740 17206
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26896 16794 26924 16934
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27448 16590 27476 16730
rect 27436 16584 27488 16590
rect 27436 16526 27488 16532
rect 27252 16516 27304 16522
rect 27252 16458 27304 16464
rect 26700 16176 26752 16182
rect 26330 16144 26386 16153
rect 26700 16118 26752 16124
rect 26330 16079 26386 16088
rect 27160 15972 27212 15978
rect 27160 15914 27212 15920
rect 27172 15706 27200 15914
rect 27160 15700 27212 15706
rect 27160 15642 27212 15648
rect 27264 15570 27292 16458
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 27540 15162 27568 17614
rect 28000 17610 28028 18770
rect 27988 17604 28040 17610
rect 27988 17546 28040 17552
rect 27607 17436 27915 17445
rect 27607 17434 27613 17436
rect 27669 17434 27693 17436
rect 27749 17434 27773 17436
rect 27829 17434 27853 17436
rect 27909 17434 27915 17436
rect 27669 17382 27671 17434
rect 27851 17382 27853 17434
rect 27607 17380 27613 17382
rect 27669 17380 27693 17382
rect 27749 17380 27773 17382
rect 27829 17380 27853 17382
rect 27909 17380 27915 17382
rect 27607 17371 27915 17380
rect 28092 17218 28120 20334
rect 28184 17542 28212 21270
rect 28276 19922 28304 21286
rect 29380 21146 29408 21830
rect 30010 21791 30066 21800
rect 29550 21720 29606 21729
rect 29550 21655 29606 21664
rect 29564 21486 29592 21655
rect 30024 21486 30052 21791
rect 29552 21480 29604 21486
rect 29552 21422 29604 21428
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29748 21146 29776 21286
rect 31494 21244 31802 21253
rect 31494 21242 31500 21244
rect 31556 21242 31580 21244
rect 31636 21242 31660 21244
rect 31716 21242 31740 21244
rect 31796 21242 31802 21244
rect 31556 21190 31558 21242
rect 31738 21190 31740 21242
rect 31494 21188 31500 21190
rect 31556 21188 31580 21190
rect 31636 21188 31660 21190
rect 31716 21188 31740 21190
rect 31796 21188 31802 21190
rect 31494 21179 31802 21188
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29736 21140 29788 21146
rect 29736 21082 29788 21088
rect 29276 20936 29328 20942
rect 29276 20878 29328 20884
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 28644 20369 28672 20402
rect 29288 20398 29316 20878
rect 29276 20392 29328 20398
rect 28630 20360 28686 20369
rect 28356 20324 28408 20330
rect 29276 20334 29328 20340
rect 28630 20295 28686 20304
rect 28816 20324 28868 20330
rect 28356 20266 28408 20272
rect 28816 20266 28868 20272
rect 28368 20058 28396 20266
rect 28828 20058 28856 20266
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28264 19916 28316 19922
rect 28264 19858 28316 19864
rect 28356 19916 28408 19922
rect 28356 19858 28408 19864
rect 29092 19916 29144 19922
rect 29092 19858 29144 19864
rect 28368 18698 28396 19858
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 29012 19394 29040 19450
rect 29104 19446 29132 19858
rect 29288 19718 29316 20334
rect 29380 19990 29408 21082
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 30024 20602 30052 20946
rect 30012 20596 30064 20602
rect 30012 20538 30064 20544
rect 29920 20324 29972 20330
rect 29920 20266 29972 20272
rect 29932 20058 29960 20266
rect 31494 20156 31802 20165
rect 31494 20154 31500 20156
rect 31556 20154 31580 20156
rect 31636 20154 31660 20156
rect 31716 20154 31740 20156
rect 31796 20154 31802 20156
rect 31556 20102 31558 20154
rect 31738 20102 31740 20154
rect 31494 20100 31500 20102
rect 31556 20100 31580 20102
rect 31636 20100 31660 20102
rect 31716 20100 31740 20102
rect 31796 20100 31802 20102
rect 31494 20091 31802 20100
rect 29920 20052 29972 20058
rect 29920 19994 29972 20000
rect 29368 19984 29420 19990
rect 29368 19926 29420 19932
rect 29644 19984 29696 19990
rect 29644 19926 29696 19932
rect 29368 19780 29420 19786
rect 29368 19722 29420 19728
rect 29276 19712 29328 19718
rect 29276 19654 29328 19660
rect 28920 19366 29040 19394
rect 29092 19440 29144 19446
rect 29092 19382 29144 19388
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28552 18222 28580 19246
rect 28920 18834 28948 19366
rect 29090 19272 29146 19281
rect 29000 19236 29052 19242
rect 29090 19207 29146 19216
rect 29000 19178 29052 19184
rect 29012 18970 29040 19178
rect 29104 19174 29132 19207
rect 29092 19168 29144 19174
rect 29092 19110 29144 19116
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 28908 18828 28960 18834
rect 28908 18770 28960 18776
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 28736 18426 28764 18770
rect 29012 18698 29040 18770
rect 28816 18692 28868 18698
rect 28816 18634 28868 18640
rect 29000 18692 29052 18698
rect 29000 18634 29052 18640
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28828 17678 28856 18634
rect 29104 18306 29132 19110
rect 29288 18850 29316 19654
rect 29380 19378 29408 19722
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29460 19346 29512 19352
rect 29460 19288 29512 19294
rect 29368 19236 29420 19242
rect 29368 19178 29420 19184
rect 29380 18970 29408 19178
rect 29472 19174 29500 19288
rect 29552 19282 29604 19288
rect 29550 19272 29552 19281
rect 29604 19272 29606 19281
rect 29550 19207 29606 19216
rect 29460 19168 29512 19174
rect 29460 19110 29512 19116
rect 29552 19168 29604 19174
rect 29552 19110 29604 19116
rect 29368 18964 29420 18970
rect 29368 18906 29420 18912
rect 29288 18834 29500 18850
rect 29184 18828 29236 18834
rect 29184 18770 29236 18776
rect 29288 18828 29512 18834
rect 29288 18822 29460 18828
rect 29196 18358 29224 18770
rect 28920 18278 29132 18306
rect 29184 18352 29236 18358
rect 29184 18294 29236 18300
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 27816 17202 28120 17218
rect 27804 17196 28120 17202
rect 27856 17190 28120 17196
rect 27804 17138 27856 17144
rect 27816 16658 27844 17138
rect 28920 17134 28948 18278
rect 29104 18154 29132 18278
rect 29288 18204 29316 18822
rect 29460 18770 29512 18776
rect 29564 18714 29592 19110
rect 29472 18686 29592 18714
rect 29472 18426 29500 18686
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18426 29592 18566
rect 29460 18420 29512 18426
rect 29460 18362 29512 18368
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29368 18216 29420 18222
rect 29288 18176 29368 18204
rect 29000 18148 29052 18154
rect 29000 18090 29052 18096
rect 29092 18148 29144 18154
rect 29092 18090 29144 18096
rect 29012 17882 29040 18090
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29288 17746 29316 18176
rect 29368 18158 29420 18164
rect 29472 17882 29500 18226
rect 29460 17876 29512 17882
rect 29460 17818 29512 17824
rect 29000 17740 29052 17746
rect 29000 17682 29052 17688
rect 29092 17740 29144 17746
rect 29092 17682 29144 17688
rect 29276 17740 29328 17746
rect 29276 17682 29328 17688
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 28908 17128 28960 17134
rect 28908 17070 28960 17076
rect 27988 17060 28040 17066
rect 27988 17002 28040 17008
rect 28080 17060 28132 17066
rect 28080 17002 28132 17008
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27607 16348 27915 16357
rect 27607 16346 27613 16348
rect 27669 16346 27693 16348
rect 27749 16346 27773 16348
rect 27829 16346 27853 16348
rect 27909 16346 27915 16348
rect 27669 16294 27671 16346
rect 27851 16294 27853 16346
rect 27607 16292 27613 16294
rect 27669 16292 27693 16294
rect 27749 16292 27773 16294
rect 27829 16292 27853 16294
rect 27909 16292 27915 16294
rect 27607 16283 27915 16292
rect 28000 15570 28028 17002
rect 28092 16794 28120 17002
rect 28080 16788 28132 16794
rect 28080 16730 28132 16736
rect 28920 16658 28948 17070
rect 29012 16998 29040 17682
rect 29104 17134 29132 17682
rect 29288 17218 29316 17682
rect 29460 17604 29512 17610
rect 29460 17546 29512 17552
rect 29196 17190 29316 17218
rect 29472 17218 29500 17546
rect 29564 17338 29592 17682
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 29472 17190 29592 17218
rect 29092 17128 29144 17134
rect 29092 17070 29144 17076
rect 29000 16992 29052 16998
rect 29000 16934 29052 16940
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 29012 16522 29040 16934
rect 29104 16794 29132 17070
rect 29196 17066 29224 17190
rect 29184 17060 29236 17066
rect 29184 17002 29236 17008
rect 29276 17060 29328 17066
rect 29276 17002 29328 17008
rect 29288 16794 29316 17002
rect 29092 16788 29144 16794
rect 29092 16730 29144 16736
rect 29276 16788 29328 16794
rect 29276 16730 29328 16736
rect 29564 16658 29592 17190
rect 29552 16652 29604 16658
rect 29552 16594 29604 16600
rect 29000 16516 29052 16522
rect 29000 16458 29052 16464
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 27988 15564 28040 15570
rect 27988 15506 28040 15512
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 27607 15260 27915 15269
rect 27607 15258 27613 15260
rect 27669 15258 27693 15260
rect 27749 15258 27773 15260
rect 27829 15258 27853 15260
rect 27909 15258 27915 15260
rect 27669 15206 27671 15258
rect 27851 15206 27853 15258
rect 27607 15204 27613 15206
rect 27669 15204 27693 15206
rect 27749 15204 27773 15206
rect 27829 15204 27853 15206
rect 27909 15204 27915 15206
rect 27607 15195 27915 15204
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25240 12838 25360 12866
rect 25976 12850 26004 13194
rect 25964 12844 26016 12850
rect 25240 12782 25268 12838
rect 25964 12786 26016 12792
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24964 11694 24992 12582
rect 25976 12434 26004 12786
rect 26252 12782 26280 13806
rect 26620 13530 26648 14418
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 26804 14074 26832 14214
rect 27607 14172 27915 14181
rect 27607 14170 27613 14172
rect 27669 14170 27693 14172
rect 27749 14170 27773 14172
rect 27829 14170 27853 14172
rect 27909 14170 27915 14172
rect 27669 14118 27671 14170
rect 27851 14118 27853 14170
rect 27607 14116 27613 14118
rect 27669 14116 27693 14118
rect 27749 14116 27773 14118
rect 27829 14116 27853 14118
rect 27909 14116 27915 14118
rect 27607 14107 27915 14116
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 28000 13462 28028 14214
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 28092 13462 28120 14010
rect 27988 13456 28040 13462
rect 27988 13398 28040 13404
rect 28080 13456 28132 13462
rect 28080 13398 28132 13404
rect 27607 13084 27915 13093
rect 27607 13082 27613 13084
rect 27669 13082 27693 13084
rect 27749 13082 27773 13084
rect 27829 13082 27853 13084
rect 27909 13082 27915 13084
rect 27669 13030 27671 13082
rect 27851 13030 27853 13082
rect 27607 13028 27613 13030
rect 27669 13028 27693 13030
rect 27749 13028 27773 13030
rect 27829 13028 27853 13030
rect 27909 13028 27915 13030
rect 27607 13019 27915 13028
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26240 12776 26292 12782
rect 26240 12718 26292 12724
rect 26436 12442 26464 12922
rect 27160 12912 27212 12918
rect 27160 12854 27212 12860
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 25700 12406 26004 12434
rect 26424 12436 26476 12442
rect 25596 12368 25648 12374
rect 25596 12310 25648 12316
rect 25608 11898 25636 12310
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25700 11830 25728 12406
rect 26424 12378 26476 12384
rect 26804 12170 26832 12582
rect 26988 12434 27016 12582
rect 26896 12406 27016 12434
rect 26896 12374 26924 12406
rect 26884 12368 26936 12374
rect 26884 12310 26936 12316
rect 27172 12238 27200 12854
rect 28092 12850 28120 13398
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 26792 12164 26844 12170
rect 26792 12106 26844 12112
rect 25688 11824 25740 11830
rect 25688 11766 25740 11772
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 25412 11212 25464 11218
rect 25412 11154 25464 11160
rect 25424 10810 25452 11154
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 23020 10532 23072 10538
rect 23020 10474 23072 10480
rect 24216 10532 24268 10538
rect 24216 10474 24268 10480
rect 23032 10266 23060 10474
rect 23720 10364 24028 10373
rect 23720 10362 23726 10364
rect 23782 10362 23806 10364
rect 23862 10362 23886 10364
rect 23942 10362 23966 10364
rect 24022 10362 24028 10364
rect 23782 10310 23784 10362
rect 23964 10310 23966 10362
rect 23720 10308 23726 10310
rect 23782 10308 23806 10310
rect 23862 10308 23886 10310
rect 23942 10308 23966 10310
rect 24022 10308 24028 10310
rect 23720 10299 24028 10308
rect 24228 10266 24256 10474
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 22020 10130 22048 10202
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 25424 9994 25452 10746
rect 25700 10606 25728 11766
rect 26804 11762 26832 12106
rect 27607 11996 27915 12005
rect 27607 11994 27613 11996
rect 27669 11994 27693 11996
rect 27749 11994 27773 11996
rect 27829 11994 27853 11996
rect 27909 11994 27915 11996
rect 27669 11942 27671 11994
rect 27851 11942 27853 11994
rect 27607 11940 27613 11942
rect 27669 11940 27693 11942
rect 27749 11940 27773 11942
rect 27829 11940 27853 11942
rect 27909 11940 27915 11942
rect 27607 11931 27915 11940
rect 26792 11756 26844 11762
rect 26792 11698 26844 11704
rect 28092 11354 28120 12786
rect 28276 12238 28304 13126
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 28276 11558 28304 12174
rect 28368 11898 28396 15506
rect 28644 15366 28672 16118
rect 29012 16114 29040 16458
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29656 15978 29684 19926
rect 29920 19168 29972 19174
rect 29920 19110 29972 19116
rect 30472 19168 30524 19174
rect 30472 19110 30524 19116
rect 29932 17814 29960 19110
rect 30484 18970 30512 19110
rect 31494 19068 31802 19077
rect 31494 19066 31500 19068
rect 31556 19066 31580 19068
rect 31636 19066 31660 19068
rect 31716 19066 31740 19068
rect 31796 19066 31802 19068
rect 31556 19014 31558 19066
rect 31738 19014 31740 19066
rect 31494 19012 31500 19014
rect 31556 19012 31580 19014
rect 31636 19012 31660 19014
rect 31716 19012 31740 19014
rect 31796 19012 31802 19014
rect 31494 19003 31802 19012
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 31494 17980 31802 17989
rect 31494 17978 31500 17980
rect 31556 17978 31580 17980
rect 31636 17978 31660 17980
rect 31716 17978 31740 17980
rect 31796 17978 31802 17980
rect 31556 17926 31558 17978
rect 31738 17926 31740 17978
rect 31494 17924 31500 17926
rect 31556 17924 31580 17926
rect 31636 17924 31660 17926
rect 31716 17924 31740 17926
rect 31796 17924 31802 17926
rect 31494 17915 31802 17924
rect 29920 17808 29972 17814
rect 29920 17750 29972 17756
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 30380 17196 30432 17202
rect 30380 17138 30432 17144
rect 29828 16992 29880 16998
rect 29828 16934 29880 16940
rect 29920 16992 29972 16998
rect 29920 16934 29972 16940
rect 29840 16658 29868 16934
rect 29932 16794 29960 16934
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 29828 16652 29880 16658
rect 29828 16594 29880 16600
rect 29644 15972 29696 15978
rect 29644 15914 29696 15920
rect 30392 15706 30420 17138
rect 31036 17105 31064 17478
rect 31022 17096 31078 17105
rect 31022 17031 31078 17040
rect 31494 16892 31802 16901
rect 31494 16890 31500 16892
rect 31556 16890 31580 16892
rect 31636 16890 31660 16892
rect 31716 16890 31740 16892
rect 31796 16890 31802 16892
rect 31556 16838 31558 16890
rect 31738 16838 31740 16890
rect 31494 16836 31500 16838
rect 31556 16836 31580 16838
rect 31636 16836 31660 16838
rect 31716 16836 31740 16838
rect 31796 16836 31802 16838
rect 31494 16827 31802 16836
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 31312 16697 31340 16730
rect 31298 16688 31354 16697
rect 31298 16623 31354 16632
rect 31494 15804 31802 15813
rect 31494 15802 31500 15804
rect 31556 15802 31580 15804
rect 31636 15802 31660 15804
rect 31716 15802 31740 15804
rect 31796 15802 31802 15804
rect 31556 15750 31558 15802
rect 31738 15750 31740 15802
rect 31494 15748 31500 15750
rect 31556 15748 31580 15750
rect 31636 15748 31660 15750
rect 31716 15748 31740 15750
rect 31796 15748 31802 15750
rect 31494 15739 31802 15748
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 30380 15700 30432 15706
rect 30380 15642 30432 15648
rect 28816 15564 28868 15570
rect 28816 15506 28868 15512
rect 28632 15360 28684 15366
rect 28632 15302 28684 15308
rect 28644 15026 28672 15302
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28644 14482 28672 14962
rect 28724 14884 28776 14890
rect 28724 14826 28776 14832
rect 28736 14482 28764 14826
rect 28828 14550 28856 15506
rect 29104 14550 29132 15642
rect 31494 14716 31802 14725
rect 31494 14714 31500 14716
rect 31556 14714 31580 14716
rect 31636 14714 31660 14716
rect 31716 14714 31740 14716
rect 31796 14714 31802 14716
rect 31556 14662 31558 14714
rect 31738 14662 31740 14714
rect 31494 14660 31500 14662
rect 31556 14660 31580 14662
rect 31636 14660 31660 14662
rect 31716 14660 31740 14662
rect 31796 14660 31802 14662
rect 31494 14651 31802 14660
rect 28816 14544 28868 14550
rect 28816 14486 28868 14492
rect 29092 14544 29144 14550
rect 29092 14486 29144 14492
rect 28632 14476 28684 14482
rect 28632 14418 28684 14424
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28540 13388 28592 13394
rect 28540 13330 28592 13336
rect 28552 12782 28580 13330
rect 28644 12782 28672 14214
rect 28736 14074 28764 14418
rect 28724 14068 28776 14074
rect 28724 14010 28776 14016
rect 28736 13394 28764 14010
rect 28828 13802 28856 14486
rect 29000 14000 29052 14006
rect 29000 13942 29052 13948
rect 28816 13796 28868 13802
rect 28816 13738 28868 13744
rect 28828 13530 28856 13738
rect 29012 13530 29040 13942
rect 29104 13734 29132 14486
rect 29184 14476 29236 14482
rect 29184 14418 29236 14424
rect 29092 13728 29144 13734
rect 29092 13670 29144 13676
rect 28816 13524 28868 13530
rect 28816 13466 28868 13472
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 28724 13388 28776 13394
rect 28724 13330 28776 13336
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28736 12850 28764 13126
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 28632 12776 28684 12782
rect 28632 12718 28684 12724
rect 28552 12434 28580 12718
rect 28828 12442 28856 13466
rect 29000 13388 29052 13394
rect 29104 13376 29132 13670
rect 29196 13394 29224 14418
rect 29460 13796 29512 13802
rect 29460 13738 29512 13744
rect 30196 13796 30248 13802
rect 30196 13738 30248 13744
rect 29472 13530 29500 13738
rect 30208 13530 30236 13738
rect 31494 13628 31802 13637
rect 31494 13626 31500 13628
rect 31556 13626 31580 13628
rect 31636 13626 31660 13628
rect 31716 13626 31740 13628
rect 31796 13626 31802 13628
rect 31556 13574 31558 13626
rect 31738 13574 31740 13626
rect 31494 13572 31500 13574
rect 31556 13572 31580 13574
rect 31636 13572 31660 13574
rect 31716 13572 31740 13574
rect 31796 13572 31802 13574
rect 31494 13563 31802 13572
rect 29460 13524 29512 13530
rect 29460 13466 29512 13472
rect 30196 13524 30248 13530
rect 30196 13466 30248 13472
rect 29052 13348 29132 13376
rect 29184 13388 29236 13394
rect 29000 13330 29052 13336
rect 29184 13330 29236 13336
rect 30104 13388 30156 13394
rect 30104 13330 30156 13336
rect 29196 12986 29224 13330
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 30116 12850 30144 13330
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 28460 12406 28580 12434
rect 28816 12436 28868 12442
rect 28356 11892 28408 11898
rect 28356 11834 28408 11840
rect 28460 11762 28488 12406
rect 28816 12378 28868 12384
rect 30012 12368 30064 12374
rect 30012 12310 30064 12316
rect 30024 11898 30052 12310
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28460 11354 28488 11698
rect 28540 11620 28592 11626
rect 28540 11562 28592 11568
rect 28552 11354 28580 11562
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28540 11348 28592 11354
rect 28540 11290 28592 11296
rect 27436 11280 27488 11286
rect 27436 11222 27488 11228
rect 27448 10810 27476 11222
rect 28736 11218 28764 11834
rect 30116 11762 30144 12786
rect 31494 12540 31802 12549
rect 31494 12538 31500 12540
rect 31556 12538 31580 12540
rect 31636 12538 31660 12540
rect 31716 12538 31740 12540
rect 31796 12538 31802 12540
rect 31556 12486 31558 12538
rect 31738 12486 31740 12538
rect 31494 12484 31500 12486
rect 31556 12484 31580 12486
rect 31636 12484 31660 12486
rect 31716 12484 31740 12486
rect 31796 12484 31802 12486
rect 31494 12475 31802 12484
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 31494 11452 31802 11461
rect 31494 11450 31500 11452
rect 31556 11450 31580 11452
rect 31636 11450 31660 11452
rect 31716 11450 31740 11452
rect 31796 11450 31802 11452
rect 31556 11398 31558 11450
rect 31738 11398 31740 11450
rect 31494 11396 31500 11398
rect 31556 11396 31580 11398
rect 31636 11396 31660 11398
rect 31716 11396 31740 11398
rect 31796 11396 31802 11398
rect 31494 11387 31802 11396
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 27607 10908 27915 10917
rect 27607 10906 27613 10908
rect 27669 10906 27693 10908
rect 27749 10906 27773 10908
rect 27829 10906 27853 10908
rect 27909 10906 27915 10908
rect 27669 10854 27671 10906
rect 27851 10854 27853 10906
rect 27607 10852 27613 10854
rect 27669 10852 27693 10854
rect 27749 10852 27773 10854
rect 27829 10852 27853 10854
rect 27909 10852 27915 10854
rect 27607 10843 27915 10852
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 31494 10364 31802 10373
rect 31494 10362 31500 10364
rect 31556 10362 31580 10364
rect 31636 10362 31660 10364
rect 31716 10362 31740 10364
rect 31796 10362 31802 10364
rect 31556 10310 31558 10362
rect 31738 10310 31740 10362
rect 31494 10308 31500 10310
rect 31556 10308 31580 10310
rect 31636 10308 31660 10310
rect 31716 10308 31740 10310
rect 31796 10308 31802 10310
rect 31494 10299 31802 10308
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 19833 9820 20141 9829
rect 19833 9818 19839 9820
rect 19895 9818 19919 9820
rect 19975 9818 19999 9820
rect 20055 9818 20079 9820
rect 20135 9818 20141 9820
rect 19895 9766 19897 9818
rect 20077 9766 20079 9818
rect 19833 9764 19839 9766
rect 19895 9764 19919 9766
rect 19975 9764 19999 9766
rect 20055 9764 20079 9766
rect 20135 9764 20141 9766
rect 19833 9755 20141 9764
rect 27607 9820 27915 9829
rect 27607 9818 27613 9820
rect 27669 9818 27693 9820
rect 27749 9818 27773 9820
rect 27829 9818 27853 9820
rect 27909 9818 27915 9820
rect 27669 9766 27671 9818
rect 27851 9766 27853 9818
rect 27607 9764 27613 9766
rect 27669 9764 27693 9766
rect 27749 9764 27773 9766
rect 27829 9764 27853 9766
rect 27909 9764 27915 9766
rect 27607 9755 27915 9764
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 8172 9276 8480 9285
rect 8172 9274 8178 9276
rect 8234 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8480 9276
rect 8234 9222 8236 9274
rect 8416 9222 8418 9274
rect 8172 9220 8178 9222
rect 8234 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8480 9222
rect 8172 9211 8480 9220
rect 15946 9276 16254 9285
rect 15946 9274 15952 9276
rect 16008 9274 16032 9276
rect 16088 9274 16112 9276
rect 16168 9274 16192 9276
rect 16248 9274 16254 9276
rect 16008 9222 16010 9274
rect 16190 9222 16192 9274
rect 15946 9220 15952 9222
rect 16008 9220 16032 9222
rect 16088 9220 16112 9222
rect 16168 9220 16192 9222
rect 16248 9220 16254 9222
rect 15946 9211 16254 9220
rect 23720 9276 24028 9285
rect 23720 9274 23726 9276
rect 23782 9274 23806 9276
rect 23862 9274 23886 9276
rect 23942 9274 23966 9276
rect 24022 9274 24028 9276
rect 23782 9222 23784 9274
rect 23964 9222 23966 9274
rect 23720 9220 23726 9222
rect 23782 9220 23806 9222
rect 23862 9220 23886 9222
rect 23942 9220 23966 9222
rect 24022 9220 24028 9222
rect 23720 9211 24028 9220
rect 31494 9276 31802 9285
rect 31494 9274 31500 9276
rect 31556 9274 31580 9276
rect 31636 9274 31660 9276
rect 31716 9274 31740 9276
rect 31796 9274 31802 9276
rect 31556 9222 31558 9274
rect 31738 9222 31740 9274
rect 31494 9220 31500 9222
rect 31556 9220 31580 9222
rect 31636 9220 31660 9222
rect 31716 9220 31740 9222
rect 31796 9220 31802 9222
rect 31494 9211 31802 9220
rect 4285 8732 4593 8741
rect 4285 8730 4291 8732
rect 4347 8730 4371 8732
rect 4427 8730 4451 8732
rect 4507 8730 4531 8732
rect 4587 8730 4593 8732
rect 4347 8678 4349 8730
rect 4529 8678 4531 8730
rect 4285 8676 4291 8678
rect 4347 8676 4371 8678
rect 4427 8676 4451 8678
rect 4507 8676 4531 8678
rect 4587 8676 4593 8678
rect 4285 8667 4593 8676
rect 12059 8732 12367 8741
rect 12059 8730 12065 8732
rect 12121 8730 12145 8732
rect 12201 8730 12225 8732
rect 12281 8730 12305 8732
rect 12361 8730 12367 8732
rect 12121 8678 12123 8730
rect 12303 8678 12305 8730
rect 12059 8676 12065 8678
rect 12121 8676 12145 8678
rect 12201 8676 12225 8678
rect 12281 8676 12305 8678
rect 12361 8676 12367 8678
rect 12059 8667 12367 8676
rect 19833 8732 20141 8741
rect 19833 8730 19839 8732
rect 19895 8730 19919 8732
rect 19975 8730 19999 8732
rect 20055 8730 20079 8732
rect 20135 8730 20141 8732
rect 19895 8678 19897 8730
rect 20077 8678 20079 8730
rect 19833 8676 19839 8678
rect 19895 8676 19919 8678
rect 19975 8676 19999 8678
rect 20055 8676 20079 8678
rect 20135 8676 20141 8678
rect 19833 8667 20141 8676
rect 27607 8732 27915 8741
rect 27607 8730 27613 8732
rect 27669 8730 27693 8732
rect 27749 8730 27773 8732
rect 27829 8730 27853 8732
rect 27909 8730 27915 8732
rect 27669 8678 27671 8730
rect 27851 8678 27853 8730
rect 27607 8676 27613 8678
rect 27669 8676 27693 8678
rect 27749 8676 27773 8678
rect 27829 8676 27853 8678
rect 27909 8676 27915 8678
rect 27607 8667 27915 8676
rect 8172 8188 8480 8197
rect 8172 8186 8178 8188
rect 8234 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8480 8188
rect 8234 8134 8236 8186
rect 8416 8134 8418 8186
rect 8172 8132 8178 8134
rect 8234 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8480 8134
rect 8172 8123 8480 8132
rect 15946 8188 16254 8197
rect 15946 8186 15952 8188
rect 16008 8186 16032 8188
rect 16088 8186 16112 8188
rect 16168 8186 16192 8188
rect 16248 8186 16254 8188
rect 16008 8134 16010 8186
rect 16190 8134 16192 8186
rect 15946 8132 15952 8134
rect 16008 8132 16032 8134
rect 16088 8132 16112 8134
rect 16168 8132 16192 8134
rect 16248 8132 16254 8134
rect 15946 8123 16254 8132
rect 23720 8188 24028 8197
rect 23720 8186 23726 8188
rect 23782 8186 23806 8188
rect 23862 8186 23886 8188
rect 23942 8186 23966 8188
rect 24022 8186 24028 8188
rect 23782 8134 23784 8186
rect 23964 8134 23966 8186
rect 23720 8132 23726 8134
rect 23782 8132 23806 8134
rect 23862 8132 23886 8134
rect 23942 8132 23966 8134
rect 24022 8132 24028 8134
rect 23720 8123 24028 8132
rect 31494 8188 31802 8197
rect 31494 8186 31500 8188
rect 31556 8186 31580 8188
rect 31636 8186 31660 8188
rect 31716 8186 31740 8188
rect 31796 8186 31802 8188
rect 31556 8134 31558 8186
rect 31738 8134 31740 8186
rect 31494 8132 31500 8134
rect 31556 8132 31580 8134
rect 31636 8132 31660 8134
rect 31716 8132 31740 8134
rect 31796 8132 31802 8134
rect 31494 8123 31802 8132
rect 4285 7644 4593 7653
rect 4285 7642 4291 7644
rect 4347 7642 4371 7644
rect 4427 7642 4451 7644
rect 4507 7642 4531 7644
rect 4587 7642 4593 7644
rect 4347 7590 4349 7642
rect 4529 7590 4531 7642
rect 4285 7588 4291 7590
rect 4347 7588 4371 7590
rect 4427 7588 4451 7590
rect 4507 7588 4531 7590
rect 4587 7588 4593 7590
rect 4285 7579 4593 7588
rect 12059 7644 12367 7653
rect 12059 7642 12065 7644
rect 12121 7642 12145 7644
rect 12201 7642 12225 7644
rect 12281 7642 12305 7644
rect 12361 7642 12367 7644
rect 12121 7590 12123 7642
rect 12303 7590 12305 7642
rect 12059 7588 12065 7590
rect 12121 7588 12145 7590
rect 12201 7588 12225 7590
rect 12281 7588 12305 7590
rect 12361 7588 12367 7590
rect 12059 7579 12367 7588
rect 19833 7644 20141 7653
rect 19833 7642 19839 7644
rect 19895 7642 19919 7644
rect 19975 7642 19999 7644
rect 20055 7642 20079 7644
rect 20135 7642 20141 7644
rect 19895 7590 19897 7642
rect 20077 7590 20079 7642
rect 19833 7588 19839 7590
rect 19895 7588 19919 7590
rect 19975 7588 19999 7590
rect 20055 7588 20079 7590
rect 20135 7588 20141 7590
rect 19833 7579 20141 7588
rect 27607 7644 27915 7653
rect 27607 7642 27613 7644
rect 27669 7642 27693 7644
rect 27749 7642 27773 7644
rect 27829 7642 27853 7644
rect 27909 7642 27915 7644
rect 27669 7590 27671 7642
rect 27851 7590 27853 7642
rect 27607 7588 27613 7590
rect 27669 7588 27693 7590
rect 27749 7588 27773 7590
rect 27829 7588 27853 7590
rect 27909 7588 27915 7590
rect 27607 7579 27915 7588
rect 8172 7100 8480 7109
rect 8172 7098 8178 7100
rect 8234 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8480 7100
rect 8234 7046 8236 7098
rect 8416 7046 8418 7098
rect 8172 7044 8178 7046
rect 8234 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8480 7046
rect 8172 7035 8480 7044
rect 15946 7100 16254 7109
rect 15946 7098 15952 7100
rect 16008 7098 16032 7100
rect 16088 7098 16112 7100
rect 16168 7098 16192 7100
rect 16248 7098 16254 7100
rect 16008 7046 16010 7098
rect 16190 7046 16192 7098
rect 15946 7044 15952 7046
rect 16008 7044 16032 7046
rect 16088 7044 16112 7046
rect 16168 7044 16192 7046
rect 16248 7044 16254 7046
rect 15946 7035 16254 7044
rect 23720 7100 24028 7109
rect 23720 7098 23726 7100
rect 23782 7098 23806 7100
rect 23862 7098 23886 7100
rect 23942 7098 23966 7100
rect 24022 7098 24028 7100
rect 23782 7046 23784 7098
rect 23964 7046 23966 7098
rect 23720 7044 23726 7046
rect 23782 7044 23806 7046
rect 23862 7044 23886 7046
rect 23942 7044 23966 7046
rect 24022 7044 24028 7046
rect 23720 7035 24028 7044
rect 31494 7100 31802 7109
rect 31494 7098 31500 7100
rect 31556 7098 31580 7100
rect 31636 7098 31660 7100
rect 31716 7098 31740 7100
rect 31796 7098 31802 7100
rect 31556 7046 31558 7098
rect 31738 7046 31740 7098
rect 31494 7044 31500 7046
rect 31556 7044 31580 7046
rect 31636 7044 31660 7046
rect 31716 7044 31740 7046
rect 31796 7044 31802 7046
rect 31494 7035 31802 7044
rect 4285 6556 4593 6565
rect 4285 6554 4291 6556
rect 4347 6554 4371 6556
rect 4427 6554 4451 6556
rect 4507 6554 4531 6556
rect 4587 6554 4593 6556
rect 4347 6502 4349 6554
rect 4529 6502 4531 6554
rect 4285 6500 4291 6502
rect 4347 6500 4371 6502
rect 4427 6500 4451 6502
rect 4507 6500 4531 6502
rect 4587 6500 4593 6502
rect 4285 6491 4593 6500
rect 12059 6556 12367 6565
rect 12059 6554 12065 6556
rect 12121 6554 12145 6556
rect 12201 6554 12225 6556
rect 12281 6554 12305 6556
rect 12361 6554 12367 6556
rect 12121 6502 12123 6554
rect 12303 6502 12305 6554
rect 12059 6500 12065 6502
rect 12121 6500 12145 6502
rect 12201 6500 12225 6502
rect 12281 6500 12305 6502
rect 12361 6500 12367 6502
rect 12059 6491 12367 6500
rect 19833 6556 20141 6565
rect 19833 6554 19839 6556
rect 19895 6554 19919 6556
rect 19975 6554 19999 6556
rect 20055 6554 20079 6556
rect 20135 6554 20141 6556
rect 19895 6502 19897 6554
rect 20077 6502 20079 6554
rect 19833 6500 19839 6502
rect 19895 6500 19919 6502
rect 19975 6500 19999 6502
rect 20055 6500 20079 6502
rect 20135 6500 20141 6502
rect 19833 6491 20141 6500
rect 27607 6556 27915 6565
rect 27607 6554 27613 6556
rect 27669 6554 27693 6556
rect 27749 6554 27773 6556
rect 27829 6554 27853 6556
rect 27909 6554 27915 6556
rect 27669 6502 27671 6554
rect 27851 6502 27853 6554
rect 27607 6500 27613 6502
rect 27669 6500 27693 6502
rect 27749 6500 27773 6502
rect 27829 6500 27853 6502
rect 27909 6500 27915 6502
rect 27607 6491 27915 6500
rect 8172 6012 8480 6021
rect 8172 6010 8178 6012
rect 8234 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8480 6012
rect 8234 5958 8236 6010
rect 8416 5958 8418 6010
rect 8172 5956 8178 5958
rect 8234 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8480 5958
rect 8172 5947 8480 5956
rect 15946 6012 16254 6021
rect 15946 6010 15952 6012
rect 16008 6010 16032 6012
rect 16088 6010 16112 6012
rect 16168 6010 16192 6012
rect 16248 6010 16254 6012
rect 16008 5958 16010 6010
rect 16190 5958 16192 6010
rect 15946 5956 15952 5958
rect 16008 5956 16032 5958
rect 16088 5956 16112 5958
rect 16168 5956 16192 5958
rect 16248 5956 16254 5958
rect 15946 5947 16254 5956
rect 23720 6012 24028 6021
rect 23720 6010 23726 6012
rect 23782 6010 23806 6012
rect 23862 6010 23886 6012
rect 23942 6010 23966 6012
rect 24022 6010 24028 6012
rect 23782 5958 23784 6010
rect 23964 5958 23966 6010
rect 23720 5956 23726 5958
rect 23782 5956 23806 5958
rect 23862 5956 23886 5958
rect 23942 5956 23966 5958
rect 24022 5956 24028 5958
rect 23720 5947 24028 5956
rect 31494 6012 31802 6021
rect 31494 6010 31500 6012
rect 31556 6010 31580 6012
rect 31636 6010 31660 6012
rect 31716 6010 31740 6012
rect 31796 6010 31802 6012
rect 31556 5958 31558 6010
rect 31738 5958 31740 6010
rect 31494 5956 31500 5958
rect 31556 5956 31580 5958
rect 31636 5956 31660 5958
rect 31716 5956 31740 5958
rect 31796 5956 31802 5958
rect 31494 5947 31802 5956
rect 4285 5468 4593 5477
rect 4285 5466 4291 5468
rect 4347 5466 4371 5468
rect 4427 5466 4451 5468
rect 4507 5466 4531 5468
rect 4587 5466 4593 5468
rect 4347 5414 4349 5466
rect 4529 5414 4531 5466
rect 4285 5412 4291 5414
rect 4347 5412 4371 5414
rect 4427 5412 4451 5414
rect 4507 5412 4531 5414
rect 4587 5412 4593 5414
rect 4285 5403 4593 5412
rect 12059 5468 12367 5477
rect 12059 5466 12065 5468
rect 12121 5466 12145 5468
rect 12201 5466 12225 5468
rect 12281 5466 12305 5468
rect 12361 5466 12367 5468
rect 12121 5414 12123 5466
rect 12303 5414 12305 5466
rect 12059 5412 12065 5414
rect 12121 5412 12145 5414
rect 12201 5412 12225 5414
rect 12281 5412 12305 5414
rect 12361 5412 12367 5414
rect 12059 5403 12367 5412
rect 19833 5468 20141 5477
rect 19833 5466 19839 5468
rect 19895 5466 19919 5468
rect 19975 5466 19999 5468
rect 20055 5466 20079 5468
rect 20135 5466 20141 5468
rect 19895 5414 19897 5466
rect 20077 5414 20079 5466
rect 19833 5412 19839 5414
rect 19895 5412 19919 5414
rect 19975 5412 19999 5414
rect 20055 5412 20079 5414
rect 20135 5412 20141 5414
rect 19833 5403 20141 5412
rect 27607 5468 27915 5477
rect 27607 5466 27613 5468
rect 27669 5466 27693 5468
rect 27749 5466 27773 5468
rect 27829 5466 27853 5468
rect 27909 5466 27915 5468
rect 27669 5414 27671 5466
rect 27851 5414 27853 5466
rect 27607 5412 27613 5414
rect 27669 5412 27693 5414
rect 27749 5412 27773 5414
rect 27829 5412 27853 5414
rect 27909 5412 27915 5414
rect 27607 5403 27915 5412
rect 8172 4924 8480 4933
rect 8172 4922 8178 4924
rect 8234 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8480 4924
rect 8234 4870 8236 4922
rect 8416 4870 8418 4922
rect 8172 4868 8178 4870
rect 8234 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8480 4870
rect 8172 4859 8480 4868
rect 15946 4924 16254 4933
rect 15946 4922 15952 4924
rect 16008 4922 16032 4924
rect 16088 4922 16112 4924
rect 16168 4922 16192 4924
rect 16248 4922 16254 4924
rect 16008 4870 16010 4922
rect 16190 4870 16192 4922
rect 15946 4868 15952 4870
rect 16008 4868 16032 4870
rect 16088 4868 16112 4870
rect 16168 4868 16192 4870
rect 16248 4868 16254 4870
rect 15946 4859 16254 4868
rect 23720 4924 24028 4933
rect 23720 4922 23726 4924
rect 23782 4922 23806 4924
rect 23862 4922 23886 4924
rect 23942 4922 23966 4924
rect 24022 4922 24028 4924
rect 23782 4870 23784 4922
rect 23964 4870 23966 4922
rect 23720 4868 23726 4870
rect 23782 4868 23806 4870
rect 23862 4868 23886 4870
rect 23942 4868 23966 4870
rect 24022 4868 24028 4870
rect 23720 4859 24028 4868
rect 31494 4924 31802 4933
rect 31494 4922 31500 4924
rect 31556 4922 31580 4924
rect 31636 4922 31660 4924
rect 31716 4922 31740 4924
rect 31796 4922 31802 4924
rect 31556 4870 31558 4922
rect 31738 4870 31740 4922
rect 31494 4868 31500 4870
rect 31556 4868 31580 4870
rect 31636 4868 31660 4870
rect 31716 4868 31740 4870
rect 31796 4868 31802 4870
rect 31494 4859 31802 4868
rect 4285 4380 4593 4389
rect 4285 4378 4291 4380
rect 4347 4378 4371 4380
rect 4427 4378 4451 4380
rect 4507 4378 4531 4380
rect 4587 4378 4593 4380
rect 4347 4326 4349 4378
rect 4529 4326 4531 4378
rect 4285 4324 4291 4326
rect 4347 4324 4371 4326
rect 4427 4324 4451 4326
rect 4507 4324 4531 4326
rect 4587 4324 4593 4326
rect 4285 4315 4593 4324
rect 12059 4380 12367 4389
rect 12059 4378 12065 4380
rect 12121 4378 12145 4380
rect 12201 4378 12225 4380
rect 12281 4378 12305 4380
rect 12361 4378 12367 4380
rect 12121 4326 12123 4378
rect 12303 4326 12305 4378
rect 12059 4324 12065 4326
rect 12121 4324 12145 4326
rect 12201 4324 12225 4326
rect 12281 4324 12305 4326
rect 12361 4324 12367 4326
rect 12059 4315 12367 4324
rect 19833 4380 20141 4389
rect 19833 4378 19839 4380
rect 19895 4378 19919 4380
rect 19975 4378 19999 4380
rect 20055 4378 20079 4380
rect 20135 4378 20141 4380
rect 19895 4326 19897 4378
rect 20077 4326 20079 4378
rect 19833 4324 19839 4326
rect 19895 4324 19919 4326
rect 19975 4324 19999 4326
rect 20055 4324 20079 4326
rect 20135 4324 20141 4326
rect 19833 4315 20141 4324
rect 27607 4380 27915 4389
rect 27607 4378 27613 4380
rect 27669 4378 27693 4380
rect 27749 4378 27773 4380
rect 27829 4378 27853 4380
rect 27909 4378 27915 4380
rect 27669 4326 27671 4378
rect 27851 4326 27853 4378
rect 27607 4324 27613 4326
rect 27669 4324 27693 4326
rect 27749 4324 27773 4326
rect 27829 4324 27853 4326
rect 27909 4324 27915 4326
rect 27607 4315 27915 4324
rect 8172 3836 8480 3845
rect 8172 3834 8178 3836
rect 8234 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8480 3836
rect 8234 3782 8236 3834
rect 8416 3782 8418 3834
rect 8172 3780 8178 3782
rect 8234 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8480 3782
rect 8172 3771 8480 3780
rect 15946 3836 16254 3845
rect 15946 3834 15952 3836
rect 16008 3834 16032 3836
rect 16088 3834 16112 3836
rect 16168 3834 16192 3836
rect 16248 3834 16254 3836
rect 16008 3782 16010 3834
rect 16190 3782 16192 3834
rect 15946 3780 15952 3782
rect 16008 3780 16032 3782
rect 16088 3780 16112 3782
rect 16168 3780 16192 3782
rect 16248 3780 16254 3782
rect 15946 3771 16254 3780
rect 23720 3836 24028 3845
rect 23720 3834 23726 3836
rect 23782 3834 23806 3836
rect 23862 3834 23886 3836
rect 23942 3834 23966 3836
rect 24022 3834 24028 3836
rect 23782 3782 23784 3834
rect 23964 3782 23966 3834
rect 23720 3780 23726 3782
rect 23782 3780 23806 3782
rect 23862 3780 23886 3782
rect 23942 3780 23966 3782
rect 24022 3780 24028 3782
rect 23720 3771 24028 3780
rect 31494 3836 31802 3845
rect 31494 3834 31500 3836
rect 31556 3834 31580 3836
rect 31636 3834 31660 3836
rect 31716 3834 31740 3836
rect 31796 3834 31802 3836
rect 31556 3782 31558 3834
rect 31738 3782 31740 3834
rect 31494 3780 31500 3782
rect 31556 3780 31580 3782
rect 31636 3780 31660 3782
rect 31716 3780 31740 3782
rect 31796 3780 31802 3782
rect 31494 3771 31802 3780
rect 4285 3292 4593 3301
rect 4285 3290 4291 3292
rect 4347 3290 4371 3292
rect 4427 3290 4451 3292
rect 4507 3290 4531 3292
rect 4587 3290 4593 3292
rect 4347 3238 4349 3290
rect 4529 3238 4531 3290
rect 4285 3236 4291 3238
rect 4347 3236 4371 3238
rect 4427 3236 4451 3238
rect 4507 3236 4531 3238
rect 4587 3236 4593 3238
rect 4285 3227 4593 3236
rect 12059 3292 12367 3301
rect 12059 3290 12065 3292
rect 12121 3290 12145 3292
rect 12201 3290 12225 3292
rect 12281 3290 12305 3292
rect 12361 3290 12367 3292
rect 12121 3238 12123 3290
rect 12303 3238 12305 3290
rect 12059 3236 12065 3238
rect 12121 3236 12145 3238
rect 12201 3236 12225 3238
rect 12281 3236 12305 3238
rect 12361 3236 12367 3238
rect 12059 3227 12367 3236
rect 19833 3292 20141 3301
rect 19833 3290 19839 3292
rect 19895 3290 19919 3292
rect 19975 3290 19999 3292
rect 20055 3290 20079 3292
rect 20135 3290 20141 3292
rect 19895 3238 19897 3290
rect 20077 3238 20079 3290
rect 19833 3236 19839 3238
rect 19895 3236 19919 3238
rect 19975 3236 19999 3238
rect 20055 3236 20079 3238
rect 20135 3236 20141 3238
rect 19833 3227 20141 3236
rect 27607 3292 27915 3301
rect 27607 3290 27613 3292
rect 27669 3290 27693 3292
rect 27749 3290 27773 3292
rect 27829 3290 27853 3292
rect 27909 3290 27915 3292
rect 27669 3238 27671 3290
rect 27851 3238 27853 3290
rect 27607 3236 27613 3238
rect 27669 3236 27693 3238
rect 27749 3236 27773 3238
rect 27829 3236 27853 3238
rect 27909 3236 27915 3238
rect 27607 3227 27915 3236
rect 8172 2748 8480 2757
rect 8172 2746 8178 2748
rect 8234 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8480 2748
rect 8234 2694 8236 2746
rect 8416 2694 8418 2746
rect 8172 2692 8178 2694
rect 8234 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8480 2694
rect 8172 2683 8480 2692
rect 15946 2748 16254 2757
rect 15946 2746 15952 2748
rect 16008 2746 16032 2748
rect 16088 2746 16112 2748
rect 16168 2746 16192 2748
rect 16248 2746 16254 2748
rect 16008 2694 16010 2746
rect 16190 2694 16192 2746
rect 15946 2692 15952 2694
rect 16008 2692 16032 2694
rect 16088 2692 16112 2694
rect 16168 2692 16192 2694
rect 16248 2692 16254 2694
rect 15946 2683 16254 2692
rect 23720 2748 24028 2757
rect 23720 2746 23726 2748
rect 23782 2746 23806 2748
rect 23862 2746 23886 2748
rect 23942 2746 23966 2748
rect 24022 2746 24028 2748
rect 23782 2694 23784 2746
rect 23964 2694 23966 2746
rect 23720 2692 23726 2694
rect 23782 2692 23806 2694
rect 23862 2692 23886 2694
rect 23942 2692 23966 2694
rect 24022 2692 24028 2694
rect 23720 2683 24028 2692
rect 31494 2748 31802 2757
rect 31494 2746 31500 2748
rect 31556 2746 31580 2748
rect 31636 2746 31660 2748
rect 31716 2746 31740 2748
rect 31796 2746 31802 2748
rect 31556 2694 31558 2746
rect 31738 2694 31740 2746
rect 31494 2692 31500 2694
rect 31556 2692 31580 2694
rect 31636 2692 31660 2694
rect 31716 2692 31740 2694
rect 31796 2692 31802 2694
rect 31494 2683 31802 2692
rect 4285 2204 4593 2213
rect 4285 2202 4291 2204
rect 4347 2202 4371 2204
rect 4427 2202 4451 2204
rect 4507 2202 4531 2204
rect 4587 2202 4593 2204
rect 4347 2150 4349 2202
rect 4529 2150 4531 2202
rect 4285 2148 4291 2150
rect 4347 2148 4371 2150
rect 4427 2148 4451 2150
rect 4507 2148 4531 2150
rect 4587 2148 4593 2150
rect 4285 2139 4593 2148
rect 12059 2204 12367 2213
rect 12059 2202 12065 2204
rect 12121 2202 12145 2204
rect 12201 2202 12225 2204
rect 12281 2202 12305 2204
rect 12361 2202 12367 2204
rect 12121 2150 12123 2202
rect 12303 2150 12305 2202
rect 12059 2148 12065 2150
rect 12121 2148 12145 2150
rect 12201 2148 12225 2150
rect 12281 2148 12305 2150
rect 12361 2148 12367 2150
rect 12059 2139 12367 2148
rect 19833 2204 20141 2213
rect 19833 2202 19839 2204
rect 19895 2202 19919 2204
rect 19975 2202 19999 2204
rect 20055 2202 20079 2204
rect 20135 2202 20141 2204
rect 19895 2150 19897 2202
rect 20077 2150 20079 2202
rect 19833 2148 19839 2150
rect 19895 2148 19919 2150
rect 19975 2148 19999 2150
rect 20055 2148 20079 2150
rect 20135 2148 20141 2150
rect 19833 2139 20141 2148
rect 27607 2204 27915 2213
rect 27607 2202 27613 2204
rect 27669 2202 27693 2204
rect 27749 2202 27773 2204
rect 27829 2202 27853 2204
rect 27909 2202 27915 2204
rect 27669 2150 27671 2202
rect 27851 2150 27853 2202
rect 27607 2148 27613 2150
rect 27669 2148 27693 2150
rect 27749 2148 27773 2150
rect 27829 2148 27853 2150
rect 27909 2148 27915 2150
rect 27607 2139 27915 2148
rect 8172 1660 8480 1669
rect 8172 1658 8178 1660
rect 8234 1658 8258 1660
rect 8314 1658 8338 1660
rect 8394 1658 8418 1660
rect 8474 1658 8480 1660
rect 8234 1606 8236 1658
rect 8416 1606 8418 1658
rect 8172 1604 8178 1606
rect 8234 1604 8258 1606
rect 8314 1604 8338 1606
rect 8394 1604 8418 1606
rect 8474 1604 8480 1606
rect 8172 1595 8480 1604
rect 15946 1660 16254 1669
rect 15946 1658 15952 1660
rect 16008 1658 16032 1660
rect 16088 1658 16112 1660
rect 16168 1658 16192 1660
rect 16248 1658 16254 1660
rect 16008 1606 16010 1658
rect 16190 1606 16192 1658
rect 15946 1604 15952 1606
rect 16008 1604 16032 1606
rect 16088 1604 16112 1606
rect 16168 1604 16192 1606
rect 16248 1604 16254 1606
rect 15946 1595 16254 1604
rect 23720 1660 24028 1669
rect 23720 1658 23726 1660
rect 23782 1658 23806 1660
rect 23862 1658 23886 1660
rect 23942 1658 23966 1660
rect 24022 1658 24028 1660
rect 23782 1606 23784 1658
rect 23964 1606 23966 1658
rect 23720 1604 23726 1606
rect 23782 1604 23806 1606
rect 23862 1604 23886 1606
rect 23942 1604 23966 1606
rect 24022 1604 24028 1606
rect 23720 1595 24028 1604
rect 31494 1660 31802 1669
rect 31494 1658 31500 1660
rect 31556 1658 31580 1660
rect 31636 1658 31660 1660
rect 31716 1658 31740 1660
rect 31796 1658 31802 1660
rect 31556 1606 31558 1658
rect 31738 1606 31740 1658
rect 31494 1604 31500 1606
rect 31556 1604 31580 1606
rect 31636 1604 31660 1606
rect 31716 1604 31740 1606
rect 31796 1604 31802 1606
rect 31494 1595 31802 1604
rect 4285 1116 4593 1125
rect 4285 1114 4291 1116
rect 4347 1114 4371 1116
rect 4427 1114 4451 1116
rect 4507 1114 4531 1116
rect 4587 1114 4593 1116
rect 4347 1062 4349 1114
rect 4529 1062 4531 1114
rect 4285 1060 4291 1062
rect 4347 1060 4371 1062
rect 4427 1060 4451 1062
rect 4507 1060 4531 1062
rect 4587 1060 4593 1062
rect 4285 1051 4593 1060
rect 12059 1116 12367 1125
rect 12059 1114 12065 1116
rect 12121 1114 12145 1116
rect 12201 1114 12225 1116
rect 12281 1114 12305 1116
rect 12361 1114 12367 1116
rect 12121 1062 12123 1114
rect 12303 1062 12305 1114
rect 12059 1060 12065 1062
rect 12121 1060 12145 1062
rect 12201 1060 12225 1062
rect 12281 1060 12305 1062
rect 12361 1060 12367 1062
rect 12059 1051 12367 1060
rect 19833 1116 20141 1125
rect 19833 1114 19839 1116
rect 19895 1114 19919 1116
rect 19975 1114 19999 1116
rect 20055 1114 20079 1116
rect 20135 1114 20141 1116
rect 19895 1062 19897 1114
rect 20077 1062 20079 1114
rect 19833 1060 19839 1062
rect 19895 1060 19919 1062
rect 19975 1060 19999 1062
rect 20055 1060 20079 1062
rect 20135 1060 20141 1062
rect 19833 1051 20141 1060
rect 27607 1116 27915 1125
rect 27607 1114 27613 1116
rect 27669 1114 27693 1116
rect 27749 1114 27773 1116
rect 27829 1114 27853 1116
rect 27909 1114 27915 1116
rect 27669 1062 27671 1114
rect 27851 1062 27853 1114
rect 27607 1060 27613 1062
rect 27669 1060 27693 1062
rect 27749 1060 27773 1062
rect 27829 1060 27853 1062
rect 27909 1060 27915 1062
rect 27607 1051 27915 1060
rect 8172 572 8480 581
rect 8172 570 8178 572
rect 8234 570 8258 572
rect 8314 570 8338 572
rect 8394 570 8418 572
rect 8474 570 8480 572
rect 8234 518 8236 570
rect 8416 518 8418 570
rect 8172 516 8178 518
rect 8234 516 8258 518
rect 8314 516 8338 518
rect 8394 516 8418 518
rect 8474 516 8480 518
rect 8172 507 8480 516
rect 15946 572 16254 581
rect 15946 570 15952 572
rect 16008 570 16032 572
rect 16088 570 16112 572
rect 16168 570 16192 572
rect 16248 570 16254 572
rect 16008 518 16010 570
rect 16190 518 16192 570
rect 15946 516 15952 518
rect 16008 516 16032 518
rect 16088 516 16112 518
rect 16168 516 16192 518
rect 16248 516 16254 518
rect 15946 507 16254 516
rect 23720 572 24028 581
rect 23720 570 23726 572
rect 23782 570 23806 572
rect 23862 570 23886 572
rect 23942 570 23966 572
rect 24022 570 24028 572
rect 23782 518 23784 570
rect 23964 518 23966 570
rect 23720 516 23726 518
rect 23782 516 23806 518
rect 23862 516 23886 518
rect 23942 516 23966 518
rect 24022 516 24028 518
rect 23720 507 24028 516
rect 31494 572 31802 581
rect 31494 570 31500 572
rect 31556 570 31580 572
rect 31636 570 31660 572
rect 31716 570 31740 572
rect 31796 570 31802 572
rect 31556 518 31558 570
rect 31738 518 31740 570
rect 31494 516 31500 518
rect 31556 516 31580 518
rect 31636 516 31660 518
rect 31716 516 31740 518
rect 31796 516 31802 518
rect 31494 507 31802 516
<< via2 >>
rect 4526 21936 4582 21992
rect 846 21800 902 21856
rect 1582 21800 1638 21856
rect 2318 21800 2374 21856
rect 3238 21800 3294 21856
rect 3790 21800 3846 21856
rect 4291 21786 4347 21788
rect 4371 21786 4427 21788
rect 4451 21786 4507 21788
rect 4531 21786 4587 21788
rect 4291 21734 4337 21786
rect 4337 21734 4347 21786
rect 4371 21734 4401 21786
rect 4401 21734 4413 21786
rect 4413 21734 4427 21786
rect 4451 21734 4465 21786
rect 4465 21734 4477 21786
rect 4477 21734 4507 21786
rect 4531 21734 4541 21786
rect 4541 21734 4587 21786
rect 4291 21732 4347 21734
rect 4371 21732 4427 21734
rect 4451 21732 4507 21734
rect 4531 21732 4587 21734
rect 8206 21936 8262 21992
rect 28998 21936 29054 21992
rect 5262 21800 5318 21856
rect 5998 21800 6054 21856
rect 6734 21800 6790 21856
rect 7470 21800 7526 21856
rect 8758 21800 8814 21856
rect 9678 21800 9734 21856
rect 10414 21800 10470 21856
rect 11150 21800 11206 21856
rect 12065 21786 12121 21788
rect 12145 21786 12201 21788
rect 12225 21786 12281 21788
rect 12305 21786 12361 21788
rect 12065 21734 12111 21786
rect 12111 21734 12121 21786
rect 12145 21734 12175 21786
rect 12175 21734 12187 21786
rect 12187 21734 12201 21786
rect 12225 21734 12239 21786
rect 12239 21734 12251 21786
rect 12251 21734 12281 21786
rect 12305 21734 12315 21786
rect 12315 21734 12361 21786
rect 12065 21732 12121 21734
rect 12145 21732 12201 21734
rect 12225 21732 12281 21734
rect 12305 21732 12361 21734
rect 19839 21786 19895 21788
rect 19919 21786 19975 21788
rect 19999 21786 20055 21788
rect 20079 21786 20135 21788
rect 19839 21734 19885 21786
rect 19885 21734 19895 21786
rect 19919 21734 19949 21786
rect 19949 21734 19961 21786
rect 19961 21734 19975 21786
rect 19999 21734 20013 21786
rect 20013 21734 20025 21786
rect 20025 21734 20055 21786
rect 20079 21734 20089 21786
rect 20089 21734 20135 21786
rect 19839 21732 19895 21734
rect 19919 21732 19975 21734
rect 19999 21732 20055 21734
rect 20079 21732 20135 21734
rect 25870 21800 25926 21856
rect 26790 21800 26846 21856
rect 28538 21800 28594 21856
rect 11886 21528 11942 21584
rect 13358 21528 13414 21584
rect 4291 20698 4347 20700
rect 4371 20698 4427 20700
rect 4451 20698 4507 20700
rect 4531 20698 4587 20700
rect 4291 20646 4337 20698
rect 4337 20646 4347 20698
rect 4371 20646 4401 20698
rect 4401 20646 4413 20698
rect 4413 20646 4427 20698
rect 4451 20646 4465 20698
rect 4465 20646 4477 20698
rect 4477 20646 4507 20698
rect 4531 20646 4541 20698
rect 4541 20646 4587 20698
rect 4291 20644 4347 20646
rect 4371 20644 4427 20646
rect 4451 20644 4507 20646
rect 4531 20644 4587 20646
rect 4291 19610 4347 19612
rect 4371 19610 4427 19612
rect 4451 19610 4507 19612
rect 4531 19610 4587 19612
rect 4291 19558 4337 19610
rect 4337 19558 4347 19610
rect 4371 19558 4401 19610
rect 4401 19558 4413 19610
rect 4413 19558 4427 19610
rect 4451 19558 4465 19610
rect 4465 19558 4477 19610
rect 4477 19558 4507 19610
rect 4531 19558 4541 19610
rect 4541 19558 4587 19610
rect 4291 19556 4347 19558
rect 4371 19556 4427 19558
rect 4451 19556 4507 19558
rect 4531 19556 4587 19558
rect 4291 18522 4347 18524
rect 4371 18522 4427 18524
rect 4451 18522 4507 18524
rect 4531 18522 4587 18524
rect 4291 18470 4337 18522
rect 4337 18470 4347 18522
rect 4371 18470 4401 18522
rect 4401 18470 4413 18522
rect 4413 18470 4427 18522
rect 4451 18470 4465 18522
rect 4465 18470 4477 18522
rect 4477 18470 4507 18522
rect 4531 18470 4541 18522
rect 4541 18470 4587 18522
rect 4291 18468 4347 18470
rect 4371 18468 4427 18470
rect 4451 18468 4507 18470
rect 4531 18468 4587 18470
rect 4986 18672 5042 18728
rect 4291 17434 4347 17436
rect 4371 17434 4427 17436
rect 4451 17434 4507 17436
rect 4531 17434 4587 17436
rect 4291 17382 4337 17434
rect 4337 17382 4347 17434
rect 4371 17382 4401 17434
rect 4401 17382 4413 17434
rect 4413 17382 4427 17434
rect 4451 17382 4465 17434
rect 4465 17382 4477 17434
rect 4477 17382 4507 17434
rect 4531 17382 4541 17434
rect 4541 17382 4587 17434
rect 4291 17380 4347 17382
rect 4371 17380 4427 17382
rect 4451 17380 4507 17382
rect 4531 17380 4587 17382
rect 4291 16346 4347 16348
rect 4371 16346 4427 16348
rect 4451 16346 4507 16348
rect 4531 16346 4587 16348
rect 4291 16294 4337 16346
rect 4337 16294 4347 16346
rect 4371 16294 4401 16346
rect 4401 16294 4413 16346
rect 4413 16294 4427 16346
rect 4451 16294 4465 16346
rect 4465 16294 4477 16346
rect 4477 16294 4507 16346
rect 4531 16294 4541 16346
rect 4541 16294 4587 16346
rect 4291 16292 4347 16294
rect 4371 16292 4427 16294
rect 4451 16292 4507 16294
rect 4531 16292 4587 16294
rect 8178 21242 8234 21244
rect 8258 21242 8314 21244
rect 8338 21242 8394 21244
rect 8418 21242 8474 21244
rect 8178 21190 8224 21242
rect 8224 21190 8234 21242
rect 8258 21190 8288 21242
rect 8288 21190 8300 21242
rect 8300 21190 8314 21242
rect 8338 21190 8352 21242
rect 8352 21190 8364 21242
rect 8364 21190 8394 21242
rect 8418 21190 8428 21242
rect 8428 21190 8474 21242
rect 8178 21188 8234 21190
rect 8258 21188 8314 21190
rect 8338 21188 8394 21190
rect 8418 21188 8474 21190
rect 5630 18944 5686 19000
rect 5354 18828 5410 18864
rect 5354 18808 5356 18828
rect 5356 18808 5408 18828
rect 5408 18808 5410 18828
rect 6458 18944 6514 19000
rect 6550 18828 6606 18864
rect 6550 18808 6552 18828
rect 6552 18808 6604 18828
rect 6604 18808 6606 18828
rect 6826 18808 6882 18864
rect 6826 18692 6882 18728
rect 6826 18672 6828 18692
rect 6828 18672 6880 18692
rect 6880 18672 6882 18692
rect 8178 20154 8234 20156
rect 8258 20154 8314 20156
rect 8338 20154 8394 20156
rect 8418 20154 8474 20156
rect 8178 20102 8224 20154
rect 8224 20102 8234 20154
rect 8258 20102 8288 20154
rect 8288 20102 8300 20154
rect 8300 20102 8314 20154
rect 8338 20102 8352 20154
rect 8352 20102 8364 20154
rect 8364 20102 8394 20154
rect 8418 20102 8428 20154
rect 8428 20102 8474 20154
rect 8178 20100 8234 20102
rect 8258 20100 8314 20102
rect 8338 20100 8394 20102
rect 8418 20100 8474 20102
rect 9218 19932 9220 19952
rect 9220 19932 9272 19952
rect 9272 19932 9274 19952
rect 9218 19896 9274 19932
rect 4291 15258 4347 15260
rect 4371 15258 4427 15260
rect 4451 15258 4507 15260
rect 4531 15258 4587 15260
rect 4291 15206 4337 15258
rect 4337 15206 4347 15258
rect 4371 15206 4401 15258
rect 4401 15206 4413 15258
rect 4413 15206 4427 15258
rect 4451 15206 4465 15258
rect 4465 15206 4477 15258
rect 4477 15206 4507 15258
rect 4531 15206 4541 15258
rect 4541 15206 4587 15258
rect 4291 15204 4347 15206
rect 4371 15204 4427 15206
rect 4451 15204 4507 15206
rect 4531 15204 4587 15206
rect 4291 14170 4347 14172
rect 4371 14170 4427 14172
rect 4451 14170 4507 14172
rect 4531 14170 4587 14172
rect 4291 14118 4337 14170
rect 4337 14118 4347 14170
rect 4371 14118 4401 14170
rect 4401 14118 4413 14170
rect 4413 14118 4427 14170
rect 4451 14118 4465 14170
rect 4465 14118 4477 14170
rect 4477 14118 4507 14170
rect 4531 14118 4541 14170
rect 4541 14118 4587 14170
rect 4291 14116 4347 14118
rect 4371 14116 4427 14118
rect 4451 14116 4507 14118
rect 4531 14116 4587 14118
rect 4291 13082 4347 13084
rect 4371 13082 4427 13084
rect 4451 13082 4507 13084
rect 4531 13082 4587 13084
rect 4291 13030 4337 13082
rect 4337 13030 4347 13082
rect 4371 13030 4401 13082
rect 4401 13030 4413 13082
rect 4413 13030 4427 13082
rect 4451 13030 4465 13082
rect 4465 13030 4477 13082
rect 4477 13030 4507 13082
rect 4531 13030 4541 13082
rect 4541 13030 4587 13082
rect 4291 13028 4347 13030
rect 4371 13028 4427 13030
rect 4451 13028 4507 13030
rect 4531 13028 4587 13030
rect 4291 11994 4347 11996
rect 4371 11994 4427 11996
rect 4451 11994 4507 11996
rect 4531 11994 4587 11996
rect 4291 11942 4337 11994
rect 4337 11942 4347 11994
rect 4371 11942 4401 11994
rect 4401 11942 4413 11994
rect 4413 11942 4427 11994
rect 4451 11942 4465 11994
rect 4465 11942 4477 11994
rect 4477 11942 4507 11994
rect 4531 11942 4541 11994
rect 4541 11942 4587 11994
rect 4291 11940 4347 11942
rect 4371 11940 4427 11942
rect 4451 11940 4507 11942
rect 4531 11940 4587 11942
rect 8942 19760 8998 19816
rect 8758 19252 8760 19272
rect 8760 19252 8812 19272
rect 8812 19252 8814 19272
rect 6826 14864 6882 14920
rect 8758 19216 8814 19252
rect 8178 19066 8234 19068
rect 8258 19066 8314 19068
rect 8338 19066 8394 19068
rect 8418 19066 8474 19068
rect 8178 19014 8224 19066
rect 8224 19014 8234 19066
rect 8258 19014 8288 19066
rect 8288 19014 8300 19066
rect 8300 19014 8314 19066
rect 8338 19014 8352 19066
rect 8352 19014 8364 19066
rect 8364 19014 8394 19066
rect 8418 19014 8428 19066
rect 8428 19014 8474 19066
rect 8178 19012 8234 19014
rect 8258 19012 8314 19014
rect 8338 19012 8394 19014
rect 8418 19012 8474 19014
rect 9862 19252 9864 19272
rect 9864 19252 9916 19272
rect 9916 19252 9918 19272
rect 9310 19080 9366 19136
rect 9218 18944 9274 19000
rect 8482 18692 8538 18728
rect 8482 18672 8484 18692
rect 8484 18672 8536 18692
rect 8536 18672 8538 18692
rect 8178 17978 8234 17980
rect 8258 17978 8314 17980
rect 8338 17978 8394 17980
rect 8418 17978 8474 17980
rect 8178 17926 8224 17978
rect 8224 17926 8234 17978
rect 8258 17926 8288 17978
rect 8288 17926 8300 17978
rect 8300 17926 8314 17978
rect 8338 17926 8352 17978
rect 8352 17926 8364 17978
rect 8364 17926 8394 17978
rect 8418 17926 8428 17978
rect 8428 17926 8474 17978
rect 8178 17924 8234 17926
rect 8258 17924 8314 17926
rect 8338 17924 8394 17926
rect 8418 17924 8474 17926
rect 8178 16890 8234 16892
rect 8258 16890 8314 16892
rect 8338 16890 8394 16892
rect 8418 16890 8474 16892
rect 8178 16838 8224 16890
rect 8224 16838 8234 16890
rect 8258 16838 8288 16890
rect 8288 16838 8300 16890
rect 8300 16838 8314 16890
rect 8338 16838 8352 16890
rect 8352 16838 8364 16890
rect 8364 16838 8394 16890
rect 8418 16838 8428 16890
rect 8428 16838 8474 16890
rect 8178 16836 8234 16838
rect 8258 16836 8314 16838
rect 8338 16836 8394 16838
rect 8418 16836 8474 16838
rect 9586 18944 9642 19000
rect 9862 19216 9918 19252
rect 9954 19080 10010 19136
rect 9586 17584 9642 17640
rect 12065 20698 12121 20700
rect 12145 20698 12201 20700
rect 12225 20698 12281 20700
rect 12305 20698 12361 20700
rect 12065 20646 12111 20698
rect 12111 20646 12121 20698
rect 12145 20646 12175 20698
rect 12175 20646 12187 20698
rect 12187 20646 12201 20698
rect 12225 20646 12239 20698
rect 12239 20646 12251 20698
rect 12251 20646 12281 20698
rect 12305 20646 12315 20698
rect 12315 20646 12361 20698
rect 12065 20644 12121 20646
rect 12145 20644 12201 20646
rect 12225 20644 12281 20646
rect 12305 20644 12361 20646
rect 8178 15802 8234 15804
rect 8258 15802 8314 15804
rect 8338 15802 8394 15804
rect 8418 15802 8474 15804
rect 8178 15750 8224 15802
rect 8224 15750 8234 15802
rect 8258 15750 8288 15802
rect 8288 15750 8300 15802
rect 8300 15750 8314 15802
rect 8338 15750 8352 15802
rect 8352 15750 8364 15802
rect 8364 15750 8394 15802
rect 8418 15750 8428 15802
rect 8428 15750 8474 15802
rect 8178 15748 8234 15750
rect 8258 15748 8314 15750
rect 8338 15748 8394 15750
rect 8418 15748 8474 15750
rect 11150 18692 11206 18728
rect 11150 18672 11152 18692
rect 11152 18672 11204 18692
rect 11204 18672 11206 18692
rect 7194 14340 7250 14376
rect 7194 14320 7196 14340
rect 7196 14320 7248 14340
rect 7248 14320 7250 14340
rect 8178 14714 8234 14716
rect 8258 14714 8314 14716
rect 8338 14714 8394 14716
rect 8418 14714 8474 14716
rect 8178 14662 8224 14714
rect 8224 14662 8234 14714
rect 8258 14662 8288 14714
rect 8288 14662 8300 14714
rect 8300 14662 8314 14714
rect 8338 14662 8352 14714
rect 8352 14662 8364 14714
rect 8364 14662 8394 14714
rect 8418 14662 8428 14714
rect 8428 14662 8474 14714
rect 8178 14660 8234 14662
rect 8258 14660 8314 14662
rect 8338 14660 8394 14662
rect 8418 14660 8474 14662
rect 8178 13626 8234 13628
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8178 13574 8224 13626
rect 8224 13574 8234 13626
rect 8258 13574 8288 13626
rect 8288 13574 8300 13626
rect 8300 13574 8314 13626
rect 8338 13574 8352 13626
rect 8352 13574 8364 13626
rect 8364 13574 8394 13626
rect 8418 13574 8428 13626
rect 8428 13574 8474 13626
rect 8178 13572 8234 13574
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 11334 17740 11390 17776
rect 11334 17720 11336 17740
rect 11336 17720 11388 17740
rect 11388 17720 11390 17740
rect 12065 19610 12121 19612
rect 12145 19610 12201 19612
rect 12225 19610 12281 19612
rect 12305 19610 12361 19612
rect 12065 19558 12111 19610
rect 12111 19558 12121 19610
rect 12145 19558 12175 19610
rect 12175 19558 12187 19610
rect 12187 19558 12201 19610
rect 12225 19558 12239 19610
rect 12239 19558 12251 19610
rect 12251 19558 12281 19610
rect 12305 19558 12315 19610
rect 12315 19558 12361 19610
rect 12065 19556 12121 19558
rect 12145 19556 12201 19558
rect 12225 19556 12281 19558
rect 12305 19556 12361 19558
rect 12065 18522 12121 18524
rect 12145 18522 12201 18524
rect 12225 18522 12281 18524
rect 12305 18522 12361 18524
rect 12065 18470 12111 18522
rect 12111 18470 12121 18522
rect 12145 18470 12175 18522
rect 12175 18470 12187 18522
rect 12187 18470 12201 18522
rect 12225 18470 12239 18522
rect 12239 18470 12251 18522
rect 12251 18470 12281 18522
rect 12305 18470 12315 18522
rect 12315 18470 12361 18522
rect 12065 18468 12121 18470
rect 12145 18468 12201 18470
rect 12225 18468 12281 18470
rect 12305 18468 12361 18470
rect 13542 19932 13544 19952
rect 13544 19932 13596 19952
rect 13596 19932 13598 19952
rect 13266 19760 13322 19816
rect 13542 19896 13598 19932
rect 11702 17584 11758 17640
rect 12065 17434 12121 17436
rect 12145 17434 12201 17436
rect 12225 17434 12281 17436
rect 12305 17434 12361 17436
rect 12065 17382 12111 17434
rect 12111 17382 12121 17434
rect 12145 17382 12175 17434
rect 12175 17382 12187 17434
rect 12187 17382 12201 17434
rect 12225 17382 12239 17434
rect 12239 17382 12251 17434
rect 12251 17382 12281 17434
rect 12305 17382 12315 17434
rect 12315 17382 12361 17434
rect 12065 17380 12121 17382
rect 12145 17380 12201 17382
rect 12225 17380 12281 17382
rect 12305 17380 12361 17382
rect 11518 14356 11520 14376
rect 11520 14356 11572 14376
rect 11572 14356 11574 14376
rect 11518 14320 11574 14356
rect 8178 12538 8234 12540
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8178 12486 8224 12538
rect 8224 12486 8234 12538
rect 8258 12486 8288 12538
rect 8288 12486 8300 12538
rect 8300 12486 8314 12538
rect 8338 12486 8352 12538
rect 8352 12486 8364 12538
rect 8364 12486 8394 12538
rect 8418 12486 8428 12538
rect 8428 12486 8474 12538
rect 8178 12484 8234 12486
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 4291 10906 4347 10908
rect 4371 10906 4427 10908
rect 4451 10906 4507 10908
rect 4531 10906 4587 10908
rect 4291 10854 4337 10906
rect 4337 10854 4347 10906
rect 4371 10854 4401 10906
rect 4401 10854 4413 10906
rect 4413 10854 4427 10906
rect 4451 10854 4465 10906
rect 4465 10854 4477 10906
rect 4477 10854 4507 10906
rect 4531 10854 4541 10906
rect 4541 10854 4587 10906
rect 4291 10852 4347 10854
rect 4371 10852 4427 10854
rect 4451 10852 4507 10854
rect 4531 10852 4587 10854
rect 8178 11450 8234 11452
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8178 11398 8224 11450
rect 8224 11398 8234 11450
rect 8258 11398 8288 11450
rect 8288 11398 8300 11450
rect 8300 11398 8314 11450
rect 8338 11398 8352 11450
rect 8352 11398 8364 11450
rect 8364 11398 8394 11450
rect 8418 11398 8428 11450
rect 8428 11398 8474 11450
rect 8178 11396 8234 11398
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 12065 16346 12121 16348
rect 12145 16346 12201 16348
rect 12225 16346 12281 16348
rect 12305 16346 12361 16348
rect 12065 16294 12111 16346
rect 12111 16294 12121 16346
rect 12145 16294 12175 16346
rect 12175 16294 12187 16346
rect 12187 16294 12201 16346
rect 12225 16294 12239 16346
rect 12239 16294 12251 16346
rect 12251 16294 12281 16346
rect 12305 16294 12315 16346
rect 12315 16294 12361 16346
rect 12065 16292 12121 16294
rect 12145 16292 12201 16294
rect 12225 16292 12281 16294
rect 12305 16292 12361 16294
rect 12065 15258 12121 15260
rect 12145 15258 12201 15260
rect 12225 15258 12281 15260
rect 12305 15258 12361 15260
rect 12065 15206 12111 15258
rect 12111 15206 12121 15258
rect 12145 15206 12175 15258
rect 12175 15206 12187 15258
rect 12187 15206 12201 15258
rect 12225 15206 12239 15258
rect 12239 15206 12251 15258
rect 12251 15206 12281 15258
rect 12305 15206 12315 15258
rect 12315 15206 12361 15258
rect 12065 15204 12121 15206
rect 12145 15204 12201 15206
rect 12225 15204 12281 15206
rect 12305 15204 12361 15206
rect 12065 14170 12121 14172
rect 12145 14170 12201 14172
rect 12225 14170 12281 14172
rect 12305 14170 12361 14172
rect 12065 14118 12111 14170
rect 12111 14118 12121 14170
rect 12145 14118 12175 14170
rect 12175 14118 12187 14170
rect 12187 14118 12201 14170
rect 12225 14118 12239 14170
rect 12239 14118 12251 14170
rect 12251 14118 12281 14170
rect 12305 14118 12315 14170
rect 12315 14118 12361 14170
rect 12065 14116 12121 14118
rect 12145 14116 12201 14118
rect 12225 14116 12281 14118
rect 12305 14116 12361 14118
rect 12065 13082 12121 13084
rect 12145 13082 12201 13084
rect 12225 13082 12281 13084
rect 12305 13082 12361 13084
rect 12065 13030 12111 13082
rect 12111 13030 12121 13082
rect 12145 13030 12175 13082
rect 12175 13030 12187 13082
rect 12187 13030 12201 13082
rect 12225 13030 12239 13082
rect 12239 13030 12251 13082
rect 12251 13030 12281 13082
rect 12305 13030 12315 13082
rect 12315 13030 12361 13082
rect 12065 13028 12121 13030
rect 12145 13028 12201 13030
rect 12225 13028 12281 13030
rect 12305 13028 12361 13030
rect 13726 19916 13782 19952
rect 13726 19896 13728 19916
rect 13728 19896 13780 19916
rect 13780 19896 13782 19916
rect 14094 20460 14150 20496
rect 14094 20440 14096 20460
rect 14096 20440 14148 20460
rect 14148 20440 14150 20460
rect 14646 20712 14702 20768
rect 14278 19796 14280 19816
rect 14280 19796 14332 19816
rect 14332 19796 14334 19816
rect 14278 19760 14334 19796
rect 13450 16088 13506 16144
rect 15290 20440 15346 20496
rect 14830 19896 14886 19952
rect 15106 19916 15162 19952
rect 15106 19896 15108 19916
rect 15108 19896 15160 19916
rect 15160 19896 15162 19916
rect 15952 21242 16008 21244
rect 16032 21242 16088 21244
rect 16112 21242 16168 21244
rect 16192 21242 16248 21244
rect 15952 21190 15998 21242
rect 15998 21190 16008 21242
rect 16032 21190 16062 21242
rect 16062 21190 16074 21242
rect 16074 21190 16088 21242
rect 16112 21190 16126 21242
rect 16126 21190 16138 21242
rect 16138 21190 16168 21242
rect 16192 21190 16202 21242
rect 16202 21190 16248 21242
rect 15952 21188 16008 21190
rect 16032 21188 16088 21190
rect 16112 21188 16168 21190
rect 16192 21188 16248 21190
rect 17130 21256 17186 21312
rect 15952 20154 16008 20156
rect 16032 20154 16088 20156
rect 16112 20154 16168 20156
rect 16192 20154 16248 20156
rect 15952 20102 15998 20154
rect 15998 20102 16008 20154
rect 16032 20102 16062 20154
rect 16062 20102 16074 20154
rect 16074 20102 16088 20154
rect 16112 20102 16126 20154
rect 16126 20102 16138 20154
rect 16138 20102 16168 20154
rect 16192 20102 16202 20154
rect 16202 20102 16248 20154
rect 15952 20100 16008 20102
rect 16032 20100 16088 20102
rect 16112 20100 16168 20102
rect 16192 20100 16248 20102
rect 13634 14900 13636 14920
rect 13636 14900 13688 14920
rect 13688 14900 13690 14920
rect 13634 14864 13690 14900
rect 12065 11994 12121 11996
rect 12145 11994 12201 11996
rect 12225 11994 12281 11996
rect 12305 11994 12361 11996
rect 12065 11942 12111 11994
rect 12111 11942 12121 11994
rect 12145 11942 12175 11994
rect 12175 11942 12187 11994
rect 12187 11942 12201 11994
rect 12225 11942 12239 11994
rect 12239 11942 12251 11994
rect 12251 11942 12281 11994
rect 12305 11942 12315 11994
rect 12315 11942 12361 11994
rect 12065 11940 12121 11942
rect 12145 11940 12201 11942
rect 12225 11940 12281 11942
rect 12305 11940 12361 11942
rect 14738 17856 14794 17912
rect 15566 19080 15622 19136
rect 15198 18844 15200 18864
rect 15200 18844 15252 18864
rect 15252 18844 15254 18864
rect 15198 18808 15254 18844
rect 15952 19066 16008 19068
rect 16032 19066 16088 19068
rect 16112 19066 16168 19068
rect 16192 19066 16248 19068
rect 15952 19014 15998 19066
rect 15998 19014 16008 19066
rect 16032 19014 16062 19066
rect 16062 19014 16074 19066
rect 16074 19014 16088 19066
rect 16112 19014 16126 19066
rect 16126 19014 16138 19066
rect 16138 19014 16168 19066
rect 16192 19014 16202 19066
rect 16202 19014 16248 19066
rect 15952 19012 16008 19014
rect 16032 19012 16088 19014
rect 16112 19012 16168 19014
rect 16192 19012 16248 19014
rect 16486 19352 16542 19408
rect 17314 20340 17316 20360
rect 17316 20340 17368 20360
rect 17368 20340 17370 20360
rect 17314 20304 17370 20340
rect 15952 17978 16008 17980
rect 16032 17978 16088 17980
rect 16112 17978 16168 17980
rect 16192 17978 16248 17980
rect 15952 17926 15998 17978
rect 15998 17926 16008 17978
rect 16032 17926 16062 17978
rect 16062 17926 16074 17978
rect 16074 17926 16088 17978
rect 16112 17926 16126 17978
rect 16126 17926 16138 17978
rect 16138 17926 16168 17978
rect 16192 17926 16202 17978
rect 16202 17926 16248 17978
rect 15952 17924 16008 17926
rect 16032 17924 16088 17926
rect 16112 17924 16168 17926
rect 16192 17924 16248 17926
rect 16578 17856 16634 17912
rect 15952 16890 16008 16892
rect 16032 16890 16088 16892
rect 16112 16890 16168 16892
rect 16192 16890 16248 16892
rect 15952 16838 15998 16890
rect 15998 16838 16008 16890
rect 16032 16838 16062 16890
rect 16062 16838 16074 16890
rect 16074 16838 16088 16890
rect 16112 16838 16126 16890
rect 16126 16838 16138 16890
rect 16138 16838 16168 16890
rect 16192 16838 16202 16890
rect 16202 16838 16248 16890
rect 15952 16836 16008 16838
rect 16032 16836 16088 16838
rect 16112 16836 16168 16838
rect 16192 16836 16248 16838
rect 15106 15988 15108 16008
rect 15108 15988 15160 16008
rect 15160 15988 15162 16008
rect 15106 15952 15162 15988
rect 8178 10362 8234 10364
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8178 10310 8224 10362
rect 8224 10310 8234 10362
rect 8258 10310 8288 10362
rect 8288 10310 8300 10362
rect 8300 10310 8314 10362
rect 8338 10310 8352 10362
rect 8352 10310 8364 10362
rect 8364 10310 8394 10362
rect 8418 10310 8428 10362
rect 8428 10310 8474 10362
rect 8178 10308 8234 10310
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 12065 10906 12121 10908
rect 12145 10906 12201 10908
rect 12225 10906 12281 10908
rect 12305 10906 12361 10908
rect 12065 10854 12111 10906
rect 12111 10854 12121 10906
rect 12145 10854 12175 10906
rect 12175 10854 12187 10906
rect 12187 10854 12201 10906
rect 12225 10854 12239 10906
rect 12239 10854 12251 10906
rect 12251 10854 12281 10906
rect 12305 10854 12315 10906
rect 12315 10854 12361 10906
rect 12065 10852 12121 10854
rect 12145 10852 12201 10854
rect 12225 10852 12281 10854
rect 12305 10852 12361 10854
rect 4291 9818 4347 9820
rect 4371 9818 4427 9820
rect 4451 9818 4507 9820
rect 4531 9818 4587 9820
rect 4291 9766 4337 9818
rect 4337 9766 4347 9818
rect 4371 9766 4401 9818
rect 4401 9766 4413 9818
rect 4413 9766 4427 9818
rect 4451 9766 4465 9818
rect 4465 9766 4477 9818
rect 4477 9766 4507 9818
rect 4531 9766 4541 9818
rect 4541 9766 4587 9818
rect 4291 9764 4347 9766
rect 4371 9764 4427 9766
rect 4451 9764 4507 9766
rect 4531 9764 4587 9766
rect 12065 9818 12121 9820
rect 12145 9818 12201 9820
rect 12225 9818 12281 9820
rect 12305 9818 12361 9820
rect 12065 9766 12111 9818
rect 12111 9766 12121 9818
rect 12145 9766 12175 9818
rect 12175 9766 12187 9818
rect 12187 9766 12201 9818
rect 12225 9766 12239 9818
rect 12239 9766 12251 9818
rect 12251 9766 12281 9818
rect 12305 9766 12315 9818
rect 12315 9766 12361 9818
rect 12065 9764 12121 9766
rect 12145 9764 12201 9766
rect 12225 9764 12281 9766
rect 12305 9764 12361 9766
rect 15952 15802 16008 15804
rect 16032 15802 16088 15804
rect 16112 15802 16168 15804
rect 16192 15802 16248 15804
rect 15952 15750 15998 15802
rect 15998 15750 16008 15802
rect 16032 15750 16062 15802
rect 16062 15750 16074 15802
rect 16074 15750 16088 15802
rect 16112 15750 16126 15802
rect 16126 15750 16138 15802
rect 16138 15750 16168 15802
rect 16192 15750 16202 15802
rect 16202 15750 16248 15802
rect 15952 15748 16008 15750
rect 16032 15748 16088 15750
rect 16112 15748 16168 15750
rect 16192 15748 16248 15750
rect 15952 14714 16008 14716
rect 16032 14714 16088 14716
rect 16112 14714 16168 14716
rect 16192 14714 16248 14716
rect 15952 14662 15998 14714
rect 15998 14662 16008 14714
rect 16032 14662 16062 14714
rect 16062 14662 16074 14714
rect 16074 14662 16088 14714
rect 16112 14662 16126 14714
rect 16126 14662 16138 14714
rect 16138 14662 16168 14714
rect 16192 14662 16202 14714
rect 16202 14662 16248 14714
rect 15952 14660 16008 14662
rect 16032 14660 16088 14662
rect 16112 14660 16168 14662
rect 16192 14660 16248 14662
rect 15952 13626 16008 13628
rect 16032 13626 16088 13628
rect 16112 13626 16168 13628
rect 16192 13626 16248 13628
rect 15952 13574 15998 13626
rect 15998 13574 16008 13626
rect 16032 13574 16062 13626
rect 16062 13574 16074 13626
rect 16074 13574 16088 13626
rect 16112 13574 16126 13626
rect 16126 13574 16138 13626
rect 16138 13574 16168 13626
rect 16192 13574 16202 13626
rect 16202 13574 16248 13626
rect 15952 13572 16008 13574
rect 16032 13572 16088 13574
rect 16112 13572 16168 13574
rect 16192 13572 16248 13574
rect 15952 12538 16008 12540
rect 16032 12538 16088 12540
rect 16112 12538 16168 12540
rect 16192 12538 16248 12540
rect 15952 12486 15998 12538
rect 15998 12486 16008 12538
rect 16032 12486 16062 12538
rect 16062 12486 16074 12538
rect 16074 12486 16088 12538
rect 16112 12486 16126 12538
rect 16126 12486 16138 12538
rect 16138 12486 16168 12538
rect 16192 12486 16202 12538
rect 16202 12486 16248 12538
rect 15952 12484 16008 12486
rect 16032 12484 16088 12486
rect 16112 12484 16168 12486
rect 16192 12484 16248 12486
rect 17958 20168 18014 20224
rect 19154 20168 19210 20224
rect 19839 20698 19895 20700
rect 19919 20698 19975 20700
rect 19999 20698 20055 20700
rect 20079 20698 20135 20700
rect 19839 20646 19885 20698
rect 19885 20646 19895 20698
rect 19919 20646 19949 20698
rect 19949 20646 19961 20698
rect 19961 20646 19975 20698
rect 19999 20646 20013 20698
rect 20013 20646 20025 20698
rect 20025 20646 20055 20698
rect 20079 20646 20089 20698
rect 20089 20646 20135 20698
rect 19839 20644 19895 20646
rect 19919 20644 19975 20646
rect 19999 20644 20055 20646
rect 20079 20644 20135 20646
rect 20258 20304 20314 20360
rect 19982 20032 20038 20088
rect 20074 19896 20130 19952
rect 19839 19610 19895 19612
rect 19919 19610 19975 19612
rect 19999 19610 20055 19612
rect 20079 19610 20135 19612
rect 19839 19558 19885 19610
rect 19885 19558 19895 19610
rect 19919 19558 19949 19610
rect 19949 19558 19961 19610
rect 19961 19558 19975 19610
rect 19999 19558 20013 19610
rect 20013 19558 20025 19610
rect 20025 19558 20055 19610
rect 20079 19558 20089 19610
rect 20089 19558 20135 19610
rect 19839 19556 19895 19558
rect 19919 19556 19975 19558
rect 19999 19556 20055 19558
rect 20079 19556 20135 19558
rect 19522 18808 19578 18864
rect 18326 17312 18382 17368
rect 18142 16904 18198 16960
rect 18142 16652 18198 16688
rect 18142 16632 18144 16652
rect 18144 16632 18196 16652
rect 18196 16632 18198 16652
rect 18510 16496 18566 16552
rect 17498 15988 17500 16008
rect 17500 15988 17552 16008
rect 17552 15988 17554 16008
rect 17498 15952 17554 15988
rect 18786 16904 18842 16960
rect 18970 17060 19026 17096
rect 18970 17040 18972 17060
rect 18972 17040 19024 17060
rect 19024 17040 19026 17060
rect 15952 11450 16008 11452
rect 16032 11450 16088 11452
rect 16112 11450 16168 11452
rect 16192 11450 16248 11452
rect 15952 11398 15998 11450
rect 15998 11398 16008 11450
rect 16032 11398 16062 11450
rect 16062 11398 16074 11450
rect 16074 11398 16088 11450
rect 16112 11398 16126 11450
rect 16126 11398 16138 11450
rect 16138 11398 16168 11450
rect 16192 11398 16202 11450
rect 16202 11398 16248 11450
rect 15952 11396 16008 11398
rect 16032 11396 16088 11398
rect 16112 11396 16168 11398
rect 16192 11396 16248 11398
rect 15952 10362 16008 10364
rect 16032 10362 16088 10364
rect 16112 10362 16168 10364
rect 16192 10362 16248 10364
rect 15952 10310 15998 10362
rect 15998 10310 16008 10362
rect 16032 10310 16062 10362
rect 16062 10310 16074 10362
rect 16074 10310 16088 10362
rect 16112 10310 16126 10362
rect 16126 10310 16138 10362
rect 16138 10310 16168 10362
rect 16192 10310 16202 10362
rect 16202 10310 16248 10362
rect 15952 10308 16008 10310
rect 16032 10308 16088 10310
rect 16112 10308 16168 10310
rect 16192 10308 16248 10310
rect 19338 18284 19394 18320
rect 19338 18264 19340 18284
rect 19340 18264 19392 18284
rect 19392 18264 19394 18284
rect 19522 18692 19578 18728
rect 19522 18672 19524 18692
rect 19524 18672 19576 18692
rect 19576 18672 19578 18692
rect 19522 18128 19578 18184
rect 19246 17312 19302 17368
rect 20350 19216 20406 19272
rect 19839 18522 19895 18524
rect 19919 18522 19975 18524
rect 19999 18522 20055 18524
rect 20079 18522 20135 18524
rect 19839 18470 19885 18522
rect 19885 18470 19895 18522
rect 19919 18470 19949 18522
rect 19949 18470 19961 18522
rect 19961 18470 19975 18522
rect 19999 18470 20013 18522
rect 20013 18470 20025 18522
rect 20025 18470 20055 18522
rect 20079 18470 20089 18522
rect 20089 18470 20135 18522
rect 19839 18468 19895 18470
rect 19919 18468 19975 18470
rect 19999 18468 20055 18470
rect 20079 18468 20135 18470
rect 19839 17434 19895 17436
rect 19919 17434 19975 17436
rect 19999 17434 20055 17436
rect 20079 17434 20135 17436
rect 19839 17382 19885 17434
rect 19885 17382 19895 17434
rect 19919 17382 19949 17434
rect 19949 17382 19961 17434
rect 19961 17382 19975 17434
rect 19999 17382 20013 17434
rect 20013 17382 20025 17434
rect 20025 17382 20055 17434
rect 20079 17382 20089 17434
rect 20089 17382 20135 17434
rect 19839 17380 19895 17382
rect 19919 17380 19975 17382
rect 19999 17380 20055 17382
rect 20079 17380 20135 17382
rect 19839 16346 19895 16348
rect 19919 16346 19975 16348
rect 19999 16346 20055 16348
rect 20079 16346 20135 16348
rect 19839 16294 19885 16346
rect 19885 16294 19895 16346
rect 19919 16294 19949 16346
rect 19949 16294 19961 16346
rect 19961 16294 19975 16346
rect 19999 16294 20013 16346
rect 20013 16294 20025 16346
rect 20025 16294 20055 16346
rect 20079 16294 20089 16346
rect 20089 16294 20135 16346
rect 19839 16292 19895 16294
rect 19919 16292 19975 16294
rect 19999 16292 20055 16294
rect 20079 16292 20135 16294
rect 20074 15988 20076 16008
rect 20076 15988 20128 16008
rect 20128 15988 20130 16008
rect 20074 15952 20130 15988
rect 19839 15258 19895 15260
rect 19919 15258 19975 15260
rect 19999 15258 20055 15260
rect 20079 15258 20135 15260
rect 19839 15206 19885 15258
rect 19885 15206 19895 15258
rect 19919 15206 19949 15258
rect 19949 15206 19961 15258
rect 19961 15206 19975 15258
rect 19999 15206 20013 15258
rect 20013 15206 20025 15258
rect 20025 15206 20055 15258
rect 20079 15206 20089 15258
rect 20089 15206 20135 15258
rect 19839 15204 19895 15206
rect 19919 15204 19975 15206
rect 19999 15204 20055 15206
rect 20079 15204 20135 15206
rect 20258 18300 20260 18320
rect 20260 18300 20312 18320
rect 20312 18300 20314 18320
rect 20258 18264 20314 18300
rect 21086 20340 21088 20360
rect 21088 20340 21140 20360
rect 21140 20340 21142 20360
rect 21086 20304 21142 20340
rect 20534 18808 20590 18864
rect 20994 19216 21050 19272
rect 19839 14170 19895 14172
rect 19919 14170 19975 14172
rect 19999 14170 20055 14172
rect 20079 14170 20135 14172
rect 19839 14118 19885 14170
rect 19885 14118 19895 14170
rect 19919 14118 19949 14170
rect 19949 14118 19961 14170
rect 19961 14118 19975 14170
rect 19999 14118 20013 14170
rect 20013 14118 20025 14170
rect 20025 14118 20055 14170
rect 20079 14118 20089 14170
rect 20089 14118 20135 14170
rect 19839 14116 19895 14118
rect 19919 14116 19975 14118
rect 19999 14116 20055 14118
rect 20079 14116 20135 14118
rect 19839 13082 19895 13084
rect 19919 13082 19975 13084
rect 19999 13082 20055 13084
rect 20079 13082 20135 13084
rect 19839 13030 19885 13082
rect 19885 13030 19895 13082
rect 19919 13030 19949 13082
rect 19949 13030 19961 13082
rect 19961 13030 19975 13082
rect 19999 13030 20013 13082
rect 20013 13030 20025 13082
rect 20025 13030 20055 13082
rect 20079 13030 20089 13082
rect 20089 13030 20135 13082
rect 19839 13028 19895 13030
rect 19919 13028 19975 13030
rect 19999 13028 20055 13030
rect 20079 13028 20135 13030
rect 19839 11994 19895 11996
rect 19919 11994 19975 11996
rect 19999 11994 20055 11996
rect 20079 11994 20135 11996
rect 19839 11942 19885 11994
rect 19885 11942 19895 11994
rect 19919 11942 19949 11994
rect 19949 11942 19961 11994
rect 19961 11942 19975 11994
rect 19999 11942 20013 11994
rect 20013 11942 20025 11994
rect 20025 11942 20055 11994
rect 20079 11942 20089 11994
rect 20089 11942 20135 11994
rect 19839 11940 19895 11942
rect 19919 11940 19975 11942
rect 19999 11940 20055 11942
rect 20079 11940 20135 11942
rect 19839 10906 19895 10908
rect 19919 10906 19975 10908
rect 19999 10906 20055 10908
rect 20079 10906 20135 10908
rect 19839 10854 19885 10906
rect 19885 10854 19895 10906
rect 19919 10854 19949 10906
rect 19949 10854 19961 10906
rect 19961 10854 19975 10906
rect 19999 10854 20013 10906
rect 20013 10854 20025 10906
rect 20025 10854 20055 10906
rect 20079 10854 20089 10906
rect 20089 10854 20135 10906
rect 19839 10852 19895 10854
rect 19919 10852 19975 10854
rect 19999 10852 20055 10854
rect 20079 10852 20135 10854
rect 23726 21242 23782 21244
rect 23806 21242 23862 21244
rect 23886 21242 23942 21244
rect 23966 21242 24022 21244
rect 23726 21190 23772 21242
rect 23772 21190 23782 21242
rect 23806 21190 23836 21242
rect 23836 21190 23848 21242
rect 23848 21190 23862 21242
rect 23886 21190 23900 21242
rect 23900 21190 23912 21242
rect 23912 21190 23942 21242
rect 23966 21190 23976 21242
rect 23976 21190 24022 21242
rect 23726 21188 23782 21190
rect 23806 21188 23862 21190
rect 23886 21188 23942 21190
rect 23966 21188 24022 21190
rect 27613 21786 27669 21788
rect 27693 21786 27749 21788
rect 27773 21786 27829 21788
rect 27853 21786 27909 21788
rect 27613 21734 27659 21786
rect 27659 21734 27669 21786
rect 27693 21734 27723 21786
rect 27723 21734 27735 21786
rect 27735 21734 27749 21786
rect 27773 21734 27787 21786
rect 27787 21734 27799 21786
rect 27799 21734 27829 21786
rect 27853 21734 27863 21786
rect 27863 21734 27909 21786
rect 27613 21732 27669 21734
rect 27693 21732 27749 21734
rect 27773 21732 27829 21734
rect 27853 21732 27909 21734
rect 22834 20168 22890 20224
rect 22650 18300 22652 18320
rect 22652 18300 22704 18320
rect 22704 18300 22706 18320
rect 22650 18264 22706 18300
rect 22374 15952 22430 16008
rect 20994 11500 20996 11520
rect 20996 11500 21048 11520
rect 21048 11500 21050 11520
rect 20994 11464 21050 11500
rect 21730 11464 21786 11520
rect 23202 16496 23258 16552
rect 23726 20154 23782 20156
rect 23806 20154 23862 20156
rect 23886 20154 23942 20156
rect 23966 20154 24022 20156
rect 23726 20102 23772 20154
rect 23772 20102 23782 20154
rect 23806 20102 23836 20154
rect 23836 20102 23848 20154
rect 23848 20102 23862 20154
rect 23886 20102 23900 20154
rect 23900 20102 23912 20154
rect 23912 20102 23942 20154
rect 23966 20102 23976 20154
rect 23976 20102 24022 20154
rect 23726 20100 23782 20102
rect 23806 20100 23862 20102
rect 23886 20100 23942 20102
rect 23966 20100 24022 20102
rect 24490 20476 24492 20496
rect 24492 20476 24544 20496
rect 24544 20476 24546 20496
rect 24490 20440 24546 20476
rect 23754 19352 23810 19408
rect 23726 19066 23782 19068
rect 23806 19066 23862 19068
rect 23886 19066 23942 19068
rect 23966 19066 24022 19068
rect 23726 19014 23772 19066
rect 23772 19014 23782 19066
rect 23806 19014 23836 19066
rect 23836 19014 23848 19066
rect 23848 19014 23862 19066
rect 23886 19014 23900 19066
rect 23900 19014 23912 19066
rect 23912 19014 23942 19066
rect 23966 19014 23976 19066
rect 23976 19014 24022 19066
rect 23726 19012 23782 19014
rect 23806 19012 23862 19014
rect 23886 19012 23942 19014
rect 23966 19012 24022 19014
rect 23570 18708 23572 18728
rect 23572 18708 23624 18728
rect 23624 18708 23626 18728
rect 23570 18672 23626 18708
rect 23570 18264 23626 18320
rect 23726 17978 23782 17980
rect 23806 17978 23862 17980
rect 23886 17978 23942 17980
rect 23966 17978 24022 17980
rect 23726 17926 23772 17978
rect 23772 17926 23782 17978
rect 23806 17926 23836 17978
rect 23836 17926 23848 17978
rect 23848 17926 23862 17978
rect 23886 17926 23900 17978
rect 23900 17926 23912 17978
rect 23912 17926 23942 17978
rect 23966 17926 23976 17978
rect 23976 17926 24022 17978
rect 23726 17924 23782 17926
rect 23806 17924 23862 17926
rect 23886 17924 23942 17926
rect 23966 17924 24022 17926
rect 23726 16890 23782 16892
rect 23806 16890 23862 16892
rect 23886 16890 23942 16892
rect 23966 16890 24022 16892
rect 23726 16838 23772 16890
rect 23772 16838 23782 16890
rect 23806 16838 23836 16890
rect 23836 16838 23848 16890
rect 23848 16838 23862 16890
rect 23886 16838 23900 16890
rect 23900 16838 23912 16890
rect 23912 16838 23942 16890
rect 23966 16838 23976 16890
rect 23976 16838 24022 16890
rect 23726 16836 23782 16838
rect 23806 16836 23862 16838
rect 23886 16836 23942 16838
rect 23966 16836 24022 16838
rect 24490 18128 24546 18184
rect 23478 16088 23534 16144
rect 24030 16088 24086 16144
rect 24858 19916 24914 19952
rect 24858 19896 24860 19916
rect 24860 19896 24912 19916
rect 24912 19896 24914 19916
rect 23726 15802 23782 15804
rect 23806 15802 23862 15804
rect 23886 15802 23942 15804
rect 23966 15802 24022 15804
rect 23726 15750 23772 15802
rect 23772 15750 23782 15802
rect 23806 15750 23836 15802
rect 23836 15750 23848 15802
rect 23848 15750 23862 15802
rect 23886 15750 23900 15802
rect 23900 15750 23912 15802
rect 23912 15750 23942 15802
rect 23966 15750 23976 15802
rect 23976 15750 24022 15802
rect 23726 15748 23782 15750
rect 23806 15748 23862 15750
rect 23886 15748 23942 15750
rect 23966 15748 24022 15750
rect 23726 14714 23782 14716
rect 23806 14714 23862 14716
rect 23886 14714 23942 14716
rect 23966 14714 24022 14716
rect 23726 14662 23772 14714
rect 23772 14662 23782 14714
rect 23806 14662 23836 14714
rect 23836 14662 23848 14714
rect 23848 14662 23862 14714
rect 23886 14662 23900 14714
rect 23900 14662 23912 14714
rect 23912 14662 23942 14714
rect 23966 14662 23976 14714
rect 23976 14662 24022 14714
rect 23726 14660 23782 14662
rect 23806 14660 23862 14662
rect 23886 14660 23942 14662
rect 23966 14660 24022 14662
rect 23726 13626 23782 13628
rect 23806 13626 23862 13628
rect 23886 13626 23942 13628
rect 23966 13626 24022 13628
rect 23726 13574 23772 13626
rect 23772 13574 23782 13626
rect 23806 13574 23836 13626
rect 23836 13574 23848 13626
rect 23848 13574 23862 13626
rect 23886 13574 23900 13626
rect 23900 13574 23912 13626
rect 23912 13574 23942 13626
rect 23966 13574 23976 13626
rect 23976 13574 24022 13626
rect 23726 13572 23782 13574
rect 23806 13572 23862 13574
rect 23886 13572 23942 13574
rect 23966 13572 24022 13574
rect 23726 12538 23782 12540
rect 23806 12538 23862 12540
rect 23886 12538 23942 12540
rect 23966 12538 24022 12540
rect 23726 12486 23772 12538
rect 23772 12486 23782 12538
rect 23806 12486 23836 12538
rect 23836 12486 23848 12538
rect 23848 12486 23862 12538
rect 23886 12486 23900 12538
rect 23900 12486 23912 12538
rect 23912 12486 23942 12538
rect 23966 12486 23976 12538
rect 23976 12486 24022 12538
rect 23726 12484 23782 12486
rect 23806 12484 23862 12486
rect 23886 12484 23942 12486
rect 23966 12484 24022 12486
rect 23726 11450 23782 11452
rect 23806 11450 23862 11452
rect 23886 11450 23942 11452
rect 23966 11450 24022 11452
rect 23726 11398 23772 11450
rect 23772 11398 23782 11450
rect 23806 11398 23836 11450
rect 23836 11398 23848 11450
rect 23848 11398 23862 11450
rect 23886 11398 23900 11450
rect 23900 11398 23912 11450
rect 23912 11398 23942 11450
rect 23966 11398 23976 11450
rect 23976 11398 24022 11450
rect 23726 11396 23782 11398
rect 23806 11396 23862 11398
rect 23886 11396 23942 11398
rect 23966 11396 24022 11398
rect 25686 16496 25742 16552
rect 27158 20440 27214 20496
rect 27613 20698 27669 20700
rect 27693 20698 27749 20700
rect 27773 20698 27829 20700
rect 27853 20698 27909 20700
rect 27613 20646 27659 20698
rect 27659 20646 27669 20698
rect 27693 20646 27723 20698
rect 27723 20646 27735 20698
rect 27735 20646 27749 20698
rect 27773 20646 27787 20698
rect 27787 20646 27799 20698
rect 27799 20646 27829 20698
rect 27853 20646 27863 20698
rect 27863 20646 27909 20698
rect 27613 20644 27669 20646
rect 27693 20644 27749 20646
rect 27773 20644 27829 20646
rect 27853 20644 27909 20646
rect 27526 20440 27582 20496
rect 27613 19610 27669 19612
rect 27693 19610 27749 19612
rect 27773 19610 27829 19612
rect 27853 19610 27909 19612
rect 27613 19558 27659 19610
rect 27659 19558 27669 19610
rect 27693 19558 27723 19610
rect 27723 19558 27735 19610
rect 27735 19558 27749 19610
rect 27773 19558 27787 19610
rect 27787 19558 27799 19610
rect 27799 19558 27829 19610
rect 27853 19558 27863 19610
rect 27863 19558 27909 19610
rect 27613 19556 27669 19558
rect 27693 19556 27749 19558
rect 27773 19556 27829 19558
rect 27853 19556 27909 19558
rect 27613 18522 27669 18524
rect 27693 18522 27749 18524
rect 27773 18522 27829 18524
rect 27853 18522 27909 18524
rect 27613 18470 27659 18522
rect 27659 18470 27669 18522
rect 27693 18470 27723 18522
rect 27723 18470 27735 18522
rect 27735 18470 27749 18522
rect 27773 18470 27787 18522
rect 27787 18470 27799 18522
rect 27799 18470 27829 18522
rect 27853 18470 27863 18522
rect 27863 18470 27909 18522
rect 27613 18468 27669 18470
rect 27693 18468 27749 18470
rect 27773 18468 27829 18470
rect 27853 18468 27909 18470
rect 26330 17720 26386 17776
rect 26330 16088 26386 16144
rect 27613 17434 27669 17436
rect 27693 17434 27749 17436
rect 27773 17434 27829 17436
rect 27853 17434 27909 17436
rect 27613 17382 27659 17434
rect 27659 17382 27669 17434
rect 27693 17382 27723 17434
rect 27723 17382 27735 17434
rect 27735 17382 27749 17434
rect 27773 17382 27787 17434
rect 27787 17382 27799 17434
rect 27799 17382 27829 17434
rect 27853 17382 27863 17434
rect 27863 17382 27909 17434
rect 27613 17380 27669 17382
rect 27693 17380 27749 17382
rect 27773 17380 27829 17382
rect 27853 17380 27909 17382
rect 30010 21800 30066 21856
rect 29550 21664 29606 21720
rect 31500 21242 31556 21244
rect 31580 21242 31636 21244
rect 31660 21242 31716 21244
rect 31740 21242 31796 21244
rect 31500 21190 31546 21242
rect 31546 21190 31556 21242
rect 31580 21190 31610 21242
rect 31610 21190 31622 21242
rect 31622 21190 31636 21242
rect 31660 21190 31674 21242
rect 31674 21190 31686 21242
rect 31686 21190 31716 21242
rect 31740 21190 31750 21242
rect 31750 21190 31796 21242
rect 31500 21188 31556 21190
rect 31580 21188 31636 21190
rect 31660 21188 31716 21190
rect 31740 21188 31796 21190
rect 28630 20304 28686 20360
rect 31500 20154 31556 20156
rect 31580 20154 31636 20156
rect 31660 20154 31716 20156
rect 31740 20154 31796 20156
rect 31500 20102 31546 20154
rect 31546 20102 31556 20154
rect 31580 20102 31610 20154
rect 31610 20102 31622 20154
rect 31622 20102 31636 20154
rect 31660 20102 31674 20154
rect 31674 20102 31686 20154
rect 31686 20102 31716 20154
rect 31740 20102 31750 20154
rect 31750 20102 31796 20154
rect 31500 20100 31556 20102
rect 31580 20100 31636 20102
rect 31660 20100 31716 20102
rect 31740 20100 31796 20102
rect 29090 19216 29146 19272
rect 29550 19230 29552 19272
rect 29552 19230 29604 19272
rect 29604 19230 29606 19272
rect 29550 19216 29606 19230
rect 27613 16346 27669 16348
rect 27693 16346 27749 16348
rect 27773 16346 27829 16348
rect 27853 16346 27909 16348
rect 27613 16294 27659 16346
rect 27659 16294 27669 16346
rect 27693 16294 27723 16346
rect 27723 16294 27735 16346
rect 27735 16294 27749 16346
rect 27773 16294 27787 16346
rect 27787 16294 27799 16346
rect 27799 16294 27829 16346
rect 27853 16294 27863 16346
rect 27863 16294 27909 16346
rect 27613 16292 27669 16294
rect 27693 16292 27749 16294
rect 27773 16292 27829 16294
rect 27853 16292 27909 16294
rect 27613 15258 27669 15260
rect 27693 15258 27749 15260
rect 27773 15258 27829 15260
rect 27853 15258 27909 15260
rect 27613 15206 27659 15258
rect 27659 15206 27669 15258
rect 27693 15206 27723 15258
rect 27723 15206 27735 15258
rect 27735 15206 27749 15258
rect 27773 15206 27787 15258
rect 27787 15206 27799 15258
rect 27799 15206 27829 15258
rect 27853 15206 27863 15258
rect 27863 15206 27909 15258
rect 27613 15204 27669 15206
rect 27693 15204 27749 15206
rect 27773 15204 27829 15206
rect 27853 15204 27909 15206
rect 27613 14170 27669 14172
rect 27693 14170 27749 14172
rect 27773 14170 27829 14172
rect 27853 14170 27909 14172
rect 27613 14118 27659 14170
rect 27659 14118 27669 14170
rect 27693 14118 27723 14170
rect 27723 14118 27735 14170
rect 27735 14118 27749 14170
rect 27773 14118 27787 14170
rect 27787 14118 27799 14170
rect 27799 14118 27829 14170
rect 27853 14118 27863 14170
rect 27863 14118 27909 14170
rect 27613 14116 27669 14118
rect 27693 14116 27749 14118
rect 27773 14116 27829 14118
rect 27853 14116 27909 14118
rect 27613 13082 27669 13084
rect 27693 13082 27749 13084
rect 27773 13082 27829 13084
rect 27853 13082 27909 13084
rect 27613 13030 27659 13082
rect 27659 13030 27669 13082
rect 27693 13030 27723 13082
rect 27723 13030 27735 13082
rect 27735 13030 27749 13082
rect 27773 13030 27787 13082
rect 27787 13030 27799 13082
rect 27799 13030 27829 13082
rect 27853 13030 27863 13082
rect 27863 13030 27909 13082
rect 27613 13028 27669 13030
rect 27693 13028 27749 13030
rect 27773 13028 27829 13030
rect 27853 13028 27909 13030
rect 23726 10362 23782 10364
rect 23806 10362 23862 10364
rect 23886 10362 23942 10364
rect 23966 10362 24022 10364
rect 23726 10310 23772 10362
rect 23772 10310 23782 10362
rect 23806 10310 23836 10362
rect 23836 10310 23848 10362
rect 23848 10310 23862 10362
rect 23886 10310 23900 10362
rect 23900 10310 23912 10362
rect 23912 10310 23942 10362
rect 23966 10310 23976 10362
rect 23976 10310 24022 10362
rect 23726 10308 23782 10310
rect 23806 10308 23862 10310
rect 23886 10308 23942 10310
rect 23966 10308 24022 10310
rect 27613 11994 27669 11996
rect 27693 11994 27749 11996
rect 27773 11994 27829 11996
rect 27853 11994 27909 11996
rect 27613 11942 27659 11994
rect 27659 11942 27669 11994
rect 27693 11942 27723 11994
rect 27723 11942 27735 11994
rect 27735 11942 27749 11994
rect 27773 11942 27787 11994
rect 27787 11942 27799 11994
rect 27799 11942 27829 11994
rect 27853 11942 27863 11994
rect 27863 11942 27909 11994
rect 27613 11940 27669 11942
rect 27693 11940 27749 11942
rect 27773 11940 27829 11942
rect 27853 11940 27909 11942
rect 31500 19066 31556 19068
rect 31580 19066 31636 19068
rect 31660 19066 31716 19068
rect 31740 19066 31796 19068
rect 31500 19014 31546 19066
rect 31546 19014 31556 19066
rect 31580 19014 31610 19066
rect 31610 19014 31622 19066
rect 31622 19014 31636 19066
rect 31660 19014 31674 19066
rect 31674 19014 31686 19066
rect 31686 19014 31716 19066
rect 31740 19014 31750 19066
rect 31750 19014 31796 19066
rect 31500 19012 31556 19014
rect 31580 19012 31636 19014
rect 31660 19012 31716 19014
rect 31740 19012 31796 19014
rect 31500 17978 31556 17980
rect 31580 17978 31636 17980
rect 31660 17978 31716 17980
rect 31740 17978 31796 17980
rect 31500 17926 31546 17978
rect 31546 17926 31556 17978
rect 31580 17926 31610 17978
rect 31610 17926 31622 17978
rect 31622 17926 31636 17978
rect 31660 17926 31674 17978
rect 31674 17926 31686 17978
rect 31686 17926 31716 17978
rect 31740 17926 31750 17978
rect 31750 17926 31796 17978
rect 31500 17924 31556 17926
rect 31580 17924 31636 17926
rect 31660 17924 31716 17926
rect 31740 17924 31796 17926
rect 31022 17040 31078 17096
rect 31500 16890 31556 16892
rect 31580 16890 31636 16892
rect 31660 16890 31716 16892
rect 31740 16890 31796 16892
rect 31500 16838 31546 16890
rect 31546 16838 31556 16890
rect 31580 16838 31610 16890
rect 31610 16838 31622 16890
rect 31622 16838 31636 16890
rect 31660 16838 31674 16890
rect 31674 16838 31686 16890
rect 31686 16838 31716 16890
rect 31740 16838 31750 16890
rect 31750 16838 31796 16890
rect 31500 16836 31556 16838
rect 31580 16836 31636 16838
rect 31660 16836 31716 16838
rect 31740 16836 31796 16838
rect 31298 16632 31354 16688
rect 31500 15802 31556 15804
rect 31580 15802 31636 15804
rect 31660 15802 31716 15804
rect 31740 15802 31796 15804
rect 31500 15750 31546 15802
rect 31546 15750 31556 15802
rect 31580 15750 31610 15802
rect 31610 15750 31622 15802
rect 31622 15750 31636 15802
rect 31660 15750 31674 15802
rect 31674 15750 31686 15802
rect 31686 15750 31716 15802
rect 31740 15750 31750 15802
rect 31750 15750 31796 15802
rect 31500 15748 31556 15750
rect 31580 15748 31636 15750
rect 31660 15748 31716 15750
rect 31740 15748 31796 15750
rect 31500 14714 31556 14716
rect 31580 14714 31636 14716
rect 31660 14714 31716 14716
rect 31740 14714 31796 14716
rect 31500 14662 31546 14714
rect 31546 14662 31556 14714
rect 31580 14662 31610 14714
rect 31610 14662 31622 14714
rect 31622 14662 31636 14714
rect 31660 14662 31674 14714
rect 31674 14662 31686 14714
rect 31686 14662 31716 14714
rect 31740 14662 31750 14714
rect 31750 14662 31796 14714
rect 31500 14660 31556 14662
rect 31580 14660 31636 14662
rect 31660 14660 31716 14662
rect 31740 14660 31796 14662
rect 31500 13626 31556 13628
rect 31580 13626 31636 13628
rect 31660 13626 31716 13628
rect 31740 13626 31796 13628
rect 31500 13574 31546 13626
rect 31546 13574 31556 13626
rect 31580 13574 31610 13626
rect 31610 13574 31622 13626
rect 31622 13574 31636 13626
rect 31660 13574 31674 13626
rect 31674 13574 31686 13626
rect 31686 13574 31716 13626
rect 31740 13574 31750 13626
rect 31750 13574 31796 13626
rect 31500 13572 31556 13574
rect 31580 13572 31636 13574
rect 31660 13572 31716 13574
rect 31740 13572 31796 13574
rect 31500 12538 31556 12540
rect 31580 12538 31636 12540
rect 31660 12538 31716 12540
rect 31740 12538 31796 12540
rect 31500 12486 31546 12538
rect 31546 12486 31556 12538
rect 31580 12486 31610 12538
rect 31610 12486 31622 12538
rect 31622 12486 31636 12538
rect 31660 12486 31674 12538
rect 31674 12486 31686 12538
rect 31686 12486 31716 12538
rect 31740 12486 31750 12538
rect 31750 12486 31796 12538
rect 31500 12484 31556 12486
rect 31580 12484 31636 12486
rect 31660 12484 31716 12486
rect 31740 12484 31796 12486
rect 31500 11450 31556 11452
rect 31580 11450 31636 11452
rect 31660 11450 31716 11452
rect 31740 11450 31796 11452
rect 31500 11398 31546 11450
rect 31546 11398 31556 11450
rect 31580 11398 31610 11450
rect 31610 11398 31622 11450
rect 31622 11398 31636 11450
rect 31660 11398 31674 11450
rect 31674 11398 31686 11450
rect 31686 11398 31716 11450
rect 31740 11398 31750 11450
rect 31750 11398 31796 11450
rect 31500 11396 31556 11398
rect 31580 11396 31636 11398
rect 31660 11396 31716 11398
rect 31740 11396 31796 11398
rect 27613 10906 27669 10908
rect 27693 10906 27749 10908
rect 27773 10906 27829 10908
rect 27853 10906 27909 10908
rect 27613 10854 27659 10906
rect 27659 10854 27669 10906
rect 27693 10854 27723 10906
rect 27723 10854 27735 10906
rect 27735 10854 27749 10906
rect 27773 10854 27787 10906
rect 27787 10854 27799 10906
rect 27799 10854 27829 10906
rect 27853 10854 27863 10906
rect 27863 10854 27909 10906
rect 27613 10852 27669 10854
rect 27693 10852 27749 10854
rect 27773 10852 27829 10854
rect 27853 10852 27909 10854
rect 31500 10362 31556 10364
rect 31580 10362 31636 10364
rect 31660 10362 31716 10364
rect 31740 10362 31796 10364
rect 31500 10310 31546 10362
rect 31546 10310 31556 10362
rect 31580 10310 31610 10362
rect 31610 10310 31622 10362
rect 31622 10310 31636 10362
rect 31660 10310 31674 10362
rect 31674 10310 31686 10362
rect 31686 10310 31716 10362
rect 31740 10310 31750 10362
rect 31750 10310 31796 10362
rect 31500 10308 31556 10310
rect 31580 10308 31636 10310
rect 31660 10308 31716 10310
rect 31740 10308 31796 10310
rect 19839 9818 19895 9820
rect 19919 9818 19975 9820
rect 19999 9818 20055 9820
rect 20079 9818 20135 9820
rect 19839 9766 19885 9818
rect 19885 9766 19895 9818
rect 19919 9766 19949 9818
rect 19949 9766 19961 9818
rect 19961 9766 19975 9818
rect 19999 9766 20013 9818
rect 20013 9766 20025 9818
rect 20025 9766 20055 9818
rect 20079 9766 20089 9818
rect 20089 9766 20135 9818
rect 19839 9764 19895 9766
rect 19919 9764 19975 9766
rect 19999 9764 20055 9766
rect 20079 9764 20135 9766
rect 27613 9818 27669 9820
rect 27693 9818 27749 9820
rect 27773 9818 27829 9820
rect 27853 9818 27909 9820
rect 27613 9766 27659 9818
rect 27659 9766 27669 9818
rect 27693 9766 27723 9818
rect 27723 9766 27735 9818
rect 27735 9766 27749 9818
rect 27773 9766 27787 9818
rect 27787 9766 27799 9818
rect 27799 9766 27829 9818
rect 27853 9766 27863 9818
rect 27863 9766 27909 9818
rect 27613 9764 27669 9766
rect 27693 9764 27749 9766
rect 27773 9764 27829 9766
rect 27853 9764 27909 9766
rect 8178 9274 8234 9276
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8178 9222 8224 9274
rect 8224 9222 8234 9274
rect 8258 9222 8288 9274
rect 8288 9222 8300 9274
rect 8300 9222 8314 9274
rect 8338 9222 8352 9274
rect 8352 9222 8364 9274
rect 8364 9222 8394 9274
rect 8418 9222 8428 9274
rect 8428 9222 8474 9274
rect 8178 9220 8234 9222
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 15952 9274 16008 9276
rect 16032 9274 16088 9276
rect 16112 9274 16168 9276
rect 16192 9274 16248 9276
rect 15952 9222 15998 9274
rect 15998 9222 16008 9274
rect 16032 9222 16062 9274
rect 16062 9222 16074 9274
rect 16074 9222 16088 9274
rect 16112 9222 16126 9274
rect 16126 9222 16138 9274
rect 16138 9222 16168 9274
rect 16192 9222 16202 9274
rect 16202 9222 16248 9274
rect 15952 9220 16008 9222
rect 16032 9220 16088 9222
rect 16112 9220 16168 9222
rect 16192 9220 16248 9222
rect 23726 9274 23782 9276
rect 23806 9274 23862 9276
rect 23886 9274 23942 9276
rect 23966 9274 24022 9276
rect 23726 9222 23772 9274
rect 23772 9222 23782 9274
rect 23806 9222 23836 9274
rect 23836 9222 23848 9274
rect 23848 9222 23862 9274
rect 23886 9222 23900 9274
rect 23900 9222 23912 9274
rect 23912 9222 23942 9274
rect 23966 9222 23976 9274
rect 23976 9222 24022 9274
rect 23726 9220 23782 9222
rect 23806 9220 23862 9222
rect 23886 9220 23942 9222
rect 23966 9220 24022 9222
rect 31500 9274 31556 9276
rect 31580 9274 31636 9276
rect 31660 9274 31716 9276
rect 31740 9274 31796 9276
rect 31500 9222 31546 9274
rect 31546 9222 31556 9274
rect 31580 9222 31610 9274
rect 31610 9222 31622 9274
rect 31622 9222 31636 9274
rect 31660 9222 31674 9274
rect 31674 9222 31686 9274
rect 31686 9222 31716 9274
rect 31740 9222 31750 9274
rect 31750 9222 31796 9274
rect 31500 9220 31556 9222
rect 31580 9220 31636 9222
rect 31660 9220 31716 9222
rect 31740 9220 31796 9222
rect 4291 8730 4347 8732
rect 4371 8730 4427 8732
rect 4451 8730 4507 8732
rect 4531 8730 4587 8732
rect 4291 8678 4337 8730
rect 4337 8678 4347 8730
rect 4371 8678 4401 8730
rect 4401 8678 4413 8730
rect 4413 8678 4427 8730
rect 4451 8678 4465 8730
rect 4465 8678 4477 8730
rect 4477 8678 4507 8730
rect 4531 8678 4541 8730
rect 4541 8678 4587 8730
rect 4291 8676 4347 8678
rect 4371 8676 4427 8678
rect 4451 8676 4507 8678
rect 4531 8676 4587 8678
rect 12065 8730 12121 8732
rect 12145 8730 12201 8732
rect 12225 8730 12281 8732
rect 12305 8730 12361 8732
rect 12065 8678 12111 8730
rect 12111 8678 12121 8730
rect 12145 8678 12175 8730
rect 12175 8678 12187 8730
rect 12187 8678 12201 8730
rect 12225 8678 12239 8730
rect 12239 8678 12251 8730
rect 12251 8678 12281 8730
rect 12305 8678 12315 8730
rect 12315 8678 12361 8730
rect 12065 8676 12121 8678
rect 12145 8676 12201 8678
rect 12225 8676 12281 8678
rect 12305 8676 12361 8678
rect 19839 8730 19895 8732
rect 19919 8730 19975 8732
rect 19999 8730 20055 8732
rect 20079 8730 20135 8732
rect 19839 8678 19885 8730
rect 19885 8678 19895 8730
rect 19919 8678 19949 8730
rect 19949 8678 19961 8730
rect 19961 8678 19975 8730
rect 19999 8678 20013 8730
rect 20013 8678 20025 8730
rect 20025 8678 20055 8730
rect 20079 8678 20089 8730
rect 20089 8678 20135 8730
rect 19839 8676 19895 8678
rect 19919 8676 19975 8678
rect 19999 8676 20055 8678
rect 20079 8676 20135 8678
rect 27613 8730 27669 8732
rect 27693 8730 27749 8732
rect 27773 8730 27829 8732
rect 27853 8730 27909 8732
rect 27613 8678 27659 8730
rect 27659 8678 27669 8730
rect 27693 8678 27723 8730
rect 27723 8678 27735 8730
rect 27735 8678 27749 8730
rect 27773 8678 27787 8730
rect 27787 8678 27799 8730
rect 27799 8678 27829 8730
rect 27853 8678 27863 8730
rect 27863 8678 27909 8730
rect 27613 8676 27669 8678
rect 27693 8676 27749 8678
rect 27773 8676 27829 8678
rect 27853 8676 27909 8678
rect 8178 8186 8234 8188
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8178 8134 8224 8186
rect 8224 8134 8234 8186
rect 8258 8134 8288 8186
rect 8288 8134 8300 8186
rect 8300 8134 8314 8186
rect 8338 8134 8352 8186
rect 8352 8134 8364 8186
rect 8364 8134 8394 8186
rect 8418 8134 8428 8186
rect 8428 8134 8474 8186
rect 8178 8132 8234 8134
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 15952 8186 16008 8188
rect 16032 8186 16088 8188
rect 16112 8186 16168 8188
rect 16192 8186 16248 8188
rect 15952 8134 15998 8186
rect 15998 8134 16008 8186
rect 16032 8134 16062 8186
rect 16062 8134 16074 8186
rect 16074 8134 16088 8186
rect 16112 8134 16126 8186
rect 16126 8134 16138 8186
rect 16138 8134 16168 8186
rect 16192 8134 16202 8186
rect 16202 8134 16248 8186
rect 15952 8132 16008 8134
rect 16032 8132 16088 8134
rect 16112 8132 16168 8134
rect 16192 8132 16248 8134
rect 23726 8186 23782 8188
rect 23806 8186 23862 8188
rect 23886 8186 23942 8188
rect 23966 8186 24022 8188
rect 23726 8134 23772 8186
rect 23772 8134 23782 8186
rect 23806 8134 23836 8186
rect 23836 8134 23848 8186
rect 23848 8134 23862 8186
rect 23886 8134 23900 8186
rect 23900 8134 23912 8186
rect 23912 8134 23942 8186
rect 23966 8134 23976 8186
rect 23976 8134 24022 8186
rect 23726 8132 23782 8134
rect 23806 8132 23862 8134
rect 23886 8132 23942 8134
rect 23966 8132 24022 8134
rect 31500 8186 31556 8188
rect 31580 8186 31636 8188
rect 31660 8186 31716 8188
rect 31740 8186 31796 8188
rect 31500 8134 31546 8186
rect 31546 8134 31556 8186
rect 31580 8134 31610 8186
rect 31610 8134 31622 8186
rect 31622 8134 31636 8186
rect 31660 8134 31674 8186
rect 31674 8134 31686 8186
rect 31686 8134 31716 8186
rect 31740 8134 31750 8186
rect 31750 8134 31796 8186
rect 31500 8132 31556 8134
rect 31580 8132 31636 8134
rect 31660 8132 31716 8134
rect 31740 8132 31796 8134
rect 4291 7642 4347 7644
rect 4371 7642 4427 7644
rect 4451 7642 4507 7644
rect 4531 7642 4587 7644
rect 4291 7590 4337 7642
rect 4337 7590 4347 7642
rect 4371 7590 4401 7642
rect 4401 7590 4413 7642
rect 4413 7590 4427 7642
rect 4451 7590 4465 7642
rect 4465 7590 4477 7642
rect 4477 7590 4507 7642
rect 4531 7590 4541 7642
rect 4541 7590 4587 7642
rect 4291 7588 4347 7590
rect 4371 7588 4427 7590
rect 4451 7588 4507 7590
rect 4531 7588 4587 7590
rect 12065 7642 12121 7644
rect 12145 7642 12201 7644
rect 12225 7642 12281 7644
rect 12305 7642 12361 7644
rect 12065 7590 12111 7642
rect 12111 7590 12121 7642
rect 12145 7590 12175 7642
rect 12175 7590 12187 7642
rect 12187 7590 12201 7642
rect 12225 7590 12239 7642
rect 12239 7590 12251 7642
rect 12251 7590 12281 7642
rect 12305 7590 12315 7642
rect 12315 7590 12361 7642
rect 12065 7588 12121 7590
rect 12145 7588 12201 7590
rect 12225 7588 12281 7590
rect 12305 7588 12361 7590
rect 19839 7642 19895 7644
rect 19919 7642 19975 7644
rect 19999 7642 20055 7644
rect 20079 7642 20135 7644
rect 19839 7590 19885 7642
rect 19885 7590 19895 7642
rect 19919 7590 19949 7642
rect 19949 7590 19961 7642
rect 19961 7590 19975 7642
rect 19999 7590 20013 7642
rect 20013 7590 20025 7642
rect 20025 7590 20055 7642
rect 20079 7590 20089 7642
rect 20089 7590 20135 7642
rect 19839 7588 19895 7590
rect 19919 7588 19975 7590
rect 19999 7588 20055 7590
rect 20079 7588 20135 7590
rect 27613 7642 27669 7644
rect 27693 7642 27749 7644
rect 27773 7642 27829 7644
rect 27853 7642 27909 7644
rect 27613 7590 27659 7642
rect 27659 7590 27669 7642
rect 27693 7590 27723 7642
rect 27723 7590 27735 7642
rect 27735 7590 27749 7642
rect 27773 7590 27787 7642
rect 27787 7590 27799 7642
rect 27799 7590 27829 7642
rect 27853 7590 27863 7642
rect 27863 7590 27909 7642
rect 27613 7588 27669 7590
rect 27693 7588 27749 7590
rect 27773 7588 27829 7590
rect 27853 7588 27909 7590
rect 8178 7098 8234 7100
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8178 7046 8224 7098
rect 8224 7046 8234 7098
rect 8258 7046 8288 7098
rect 8288 7046 8300 7098
rect 8300 7046 8314 7098
rect 8338 7046 8352 7098
rect 8352 7046 8364 7098
rect 8364 7046 8394 7098
rect 8418 7046 8428 7098
rect 8428 7046 8474 7098
rect 8178 7044 8234 7046
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 15952 7098 16008 7100
rect 16032 7098 16088 7100
rect 16112 7098 16168 7100
rect 16192 7098 16248 7100
rect 15952 7046 15998 7098
rect 15998 7046 16008 7098
rect 16032 7046 16062 7098
rect 16062 7046 16074 7098
rect 16074 7046 16088 7098
rect 16112 7046 16126 7098
rect 16126 7046 16138 7098
rect 16138 7046 16168 7098
rect 16192 7046 16202 7098
rect 16202 7046 16248 7098
rect 15952 7044 16008 7046
rect 16032 7044 16088 7046
rect 16112 7044 16168 7046
rect 16192 7044 16248 7046
rect 23726 7098 23782 7100
rect 23806 7098 23862 7100
rect 23886 7098 23942 7100
rect 23966 7098 24022 7100
rect 23726 7046 23772 7098
rect 23772 7046 23782 7098
rect 23806 7046 23836 7098
rect 23836 7046 23848 7098
rect 23848 7046 23862 7098
rect 23886 7046 23900 7098
rect 23900 7046 23912 7098
rect 23912 7046 23942 7098
rect 23966 7046 23976 7098
rect 23976 7046 24022 7098
rect 23726 7044 23782 7046
rect 23806 7044 23862 7046
rect 23886 7044 23942 7046
rect 23966 7044 24022 7046
rect 31500 7098 31556 7100
rect 31580 7098 31636 7100
rect 31660 7098 31716 7100
rect 31740 7098 31796 7100
rect 31500 7046 31546 7098
rect 31546 7046 31556 7098
rect 31580 7046 31610 7098
rect 31610 7046 31622 7098
rect 31622 7046 31636 7098
rect 31660 7046 31674 7098
rect 31674 7046 31686 7098
rect 31686 7046 31716 7098
rect 31740 7046 31750 7098
rect 31750 7046 31796 7098
rect 31500 7044 31556 7046
rect 31580 7044 31636 7046
rect 31660 7044 31716 7046
rect 31740 7044 31796 7046
rect 4291 6554 4347 6556
rect 4371 6554 4427 6556
rect 4451 6554 4507 6556
rect 4531 6554 4587 6556
rect 4291 6502 4337 6554
rect 4337 6502 4347 6554
rect 4371 6502 4401 6554
rect 4401 6502 4413 6554
rect 4413 6502 4427 6554
rect 4451 6502 4465 6554
rect 4465 6502 4477 6554
rect 4477 6502 4507 6554
rect 4531 6502 4541 6554
rect 4541 6502 4587 6554
rect 4291 6500 4347 6502
rect 4371 6500 4427 6502
rect 4451 6500 4507 6502
rect 4531 6500 4587 6502
rect 12065 6554 12121 6556
rect 12145 6554 12201 6556
rect 12225 6554 12281 6556
rect 12305 6554 12361 6556
rect 12065 6502 12111 6554
rect 12111 6502 12121 6554
rect 12145 6502 12175 6554
rect 12175 6502 12187 6554
rect 12187 6502 12201 6554
rect 12225 6502 12239 6554
rect 12239 6502 12251 6554
rect 12251 6502 12281 6554
rect 12305 6502 12315 6554
rect 12315 6502 12361 6554
rect 12065 6500 12121 6502
rect 12145 6500 12201 6502
rect 12225 6500 12281 6502
rect 12305 6500 12361 6502
rect 19839 6554 19895 6556
rect 19919 6554 19975 6556
rect 19999 6554 20055 6556
rect 20079 6554 20135 6556
rect 19839 6502 19885 6554
rect 19885 6502 19895 6554
rect 19919 6502 19949 6554
rect 19949 6502 19961 6554
rect 19961 6502 19975 6554
rect 19999 6502 20013 6554
rect 20013 6502 20025 6554
rect 20025 6502 20055 6554
rect 20079 6502 20089 6554
rect 20089 6502 20135 6554
rect 19839 6500 19895 6502
rect 19919 6500 19975 6502
rect 19999 6500 20055 6502
rect 20079 6500 20135 6502
rect 27613 6554 27669 6556
rect 27693 6554 27749 6556
rect 27773 6554 27829 6556
rect 27853 6554 27909 6556
rect 27613 6502 27659 6554
rect 27659 6502 27669 6554
rect 27693 6502 27723 6554
rect 27723 6502 27735 6554
rect 27735 6502 27749 6554
rect 27773 6502 27787 6554
rect 27787 6502 27799 6554
rect 27799 6502 27829 6554
rect 27853 6502 27863 6554
rect 27863 6502 27909 6554
rect 27613 6500 27669 6502
rect 27693 6500 27749 6502
rect 27773 6500 27829 6502
rect 27853 6500 27909 6502
rect 8178 6010 8234 6012
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8178 5958 8224 6010
rect 8224 5958 8234 6010
rect 8258 5958 8288 6010
rect 8288 5958 8300 6010
rect 8300 5958 8314 6010
rect 8338 5958 8352 6010
rect 8352 5958 8364 6010
rect 8364 5958 8394 6010
rect 8418 5958 8428 6010
rect 8428 5958 8474 6010
rect 8178 5956 8234 5958
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 15952 6010 16008 6012
rect 16032 6010 16088 6012
rect 16112 6010 16168 6012
rect 16192 6010 16248 6012
rect 15952 5958 15998 6010
rect 15998 5958 16008 6010
rect 16032 5958 16062 6010
rect 16062 5958 16074 6010
rect 16074 5958 16088 6010
rect 16112 5958 16126 6010
rect 16126 5958 16138 6010
rect 16138 5958 16168 6010
rect 16192 5958 16202 6010
rect 16202 5958 16248 6010
rect 15952 5956 16008 5958
rect 16032 5956 16088 5958
rect 16112 5956 16168 5958
rect 16192 5956 16248 5958
rect 23726 6010 23782 6012
rect 23806 6010 23862 6012
rect 23886 6010 23942 6012
rect 23966 6010 24022 6012
rect 23726 5958 23772 6010
rect 23772 5958 23782 6010
rect 23806 5958 23836 6010
rect 23836 5958 23848 6010
rect 23848 5958 23862 6010
rect 23886 5958 23900 6010
rect 23900 5958 23912 6010
rect 23912 5958 23942 6010
rect 23966 5958 23976 6010
rect 23976 5958 24022 6010
rect 23726 5956 23782 5958
rect 23806 5956 23862 5958
rect 23886 5956 23942 5958
rect 23966 5956 24022 5958
rect 31500 6010 31556 6012
rect 31580 6010 31636 6012
rect 31660 6010 31716 6012
rect 31740 6010 31796 6012
rect 31500 5958 31546 6010
rect 31546 5958 31556 6010
rect 31580 5958 31610 6010
rect 31610 5958 31622 6010
rect 31622 5958 31636 6010
rect 31660 5958 31674 6010
rect 31674 5958 31686 6010
rect 31686 5958 31716 6010
rect 31740 5958 31750 6010
rect 31750 5958 31796 6010
rect 31500 5956 31556 5958
rect 31580 5956 31636 5958
rect 31660 5956 31716 5958
rect 31740 5956 31796 5958
rect 4291 5466 4347 5468
rect 4371 5466 4427 5468
rect 4451 5466 4507 5468
rect 4531 5466 4587 5468
rect 4291 5414 4337 5466
rect 4337 5414 4347 5466
rect 4371 5414 4401 5466
rect 4401 5414 4413 5466
rect 4413 5414 4427 5466
rect 4451 5414 4465 5466
rect 4465 5414 4477 5466
rect 4477 5414 4507 5466
rect 4531 5414 4541 5466
rect 4541 5414 4587 5466
rect 4291 5412 4347 5414
rect 4371 5412 4427 5414
rect 4451 5412 4507 5414
rect 4531 5412 4587 5414
rect 12065 5466 12121 5468
rect 12145 5466 12201 5468
rect 12225 5466 12281 5468
rect 12305 5466 12361 5468
rect 12065 5414 12111 5466
rect 12111 5414 12121 5466
rect 12145 5414 12175 5466
rect 12175 5414 12187 5466
rect 12187 5414 12201 5466
rect 12225 5414 12239 5466
rect 12239 5414 12251 5466
rect 12251 5414 12281 5466
rect 12305 5414 12315 5466
rect 12315 5414 12361 5466
rect 12065 5412 12121 5414
rect 12145 5412 12201 5414
rect 12225 5412 12281 5414
rect 12305 5412 12361 5414
rect 19839 5466 19895 5468
rect 19919 5466 19975 5468
rect 19999 5466 20055 5468
rect 20079 5466 20135 5468
rect 19839 5414 19885 5466
rect 19885 5414 19895 5466
rect 19919 5414 19949 5466
rect 19949 5414 19961 5466
rect 19961 5414 19975 5466
rect 19999 5414 20013 5466
rect 20013 5414 20025 5466
rect 20025 5414 20055 5466
rect 20079 5414 20089 5466
rect 20089 5414 20135 5466
rect 19839 5412 19895 5414
rect 19919 5412 19975 5414
rect 19999 5412 20055 5414
rect 20079 5412 20135 5414
rect 27613 5466 27669 5468
rect 27693 5466 27749 5468
rect 27773 5466 27829 5468
rect 27853 5466 27909 5468
rect 27613 5414 27659 5466
rect 27659 5414 27669 5466
rect 27693 5414 27723 5466
rect 27723 5414 27735 5466
rect 27735 5414 27749 5466
rect 27773 5414 27787 5466
rect 27787 5414 27799 5466
rect 27799 5414 27829 5466
rect 27853 5414 27863 5466
rect 27863 5414 27909 5466
rect 27613 5412 27669 5414
rect 27693 5412 27749 5414
rect 27773 5412 27829 5414
rect 27853 5412 27909 5414
rect 8178 4922 8234 4924
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8178 4870 8224 4922
rect 8224 4870 8234 4922
rect 8258 4870 8288 4922
rect 8288 4870 8300 4922
rect 8300 4870 8314 4922
rect 8338 4870 8352 4922
rect 8352 4870 8364 4922
rect 8364 4870 8394 4922
rect 8418 4870 8428 4922
rect 8428 4870 8474 4922
rect 8178 4868 8234 4870
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 15952 4922 16008 4924
rect 16032 4922 16088 4924
rect 16112 4922 16168 4924
rect 16192 4922 16248 4924
rect 15952 4870 15998 4922
rect 15998 4870 16008 4922
rect 16032 4870 16062 4922
rect 16062 4870 16074 4922
rect 16074 4870 16088 4922
rect 16112 4870 16126 4922
rect 16126 4870 16138 4922
rect 16138 4870 16168 4922
rect 16192 4870 16202 4922
rect 16202 4870 16248 4922
rect 15952 4868 16008 4870
rect 16032 4868 16088 4870
rect 16112 4868 16168 4870
rect 16192 4868 16248 4870
rect 23726 4922 23782 4924
rect 23806 4922 23862 4924
rect 23886 4922 23942 4924
rect 23966 4922 24022 4924
rect 23726 4870 23772 4922
rect 23772 4870 23782 4922
rect 23806 4870 23836 4922
rect 23836 4870 23848 4922
rect 23848 4870 23862 4922
rect 23886 4870 23900 4922
rect 23900 4870 23912 4922
rect 23912 4870 23942 4922
rect 23966 4870 23976 4922
rect 23976 4870 24022 4922
rect 23726 4868 23782 4870
rect 23806 4868 23862 4870
rect 23886 4868 23942 4870
rect 23966 4868 24022 4870
rect 31500 4922 31556 4924
rect 31580 4922 31636 4924
rect 31660 4922 31716 4924
rect 31740 4922 31796 4924
rect 31500 4870 31546 4922
rect 31546 4870 31556 4922
rect 31580 4870 31610 4922
rect 31610 4870 31622 4922
rect 31622 4870 31636 4922
rect 31660 4870 31674 4922
rect 31674 4870 31686 4922
rect 31686 4870 31716 4922
rect 31740 4870 31750 4922
rect 31750 4870 31796 4922
rect 31500 4868 31556 4870
rect 31580 4868 31636 4870
rect 31660 4868 31716 4870
rect 31740 4868 31796 4870
rect 4291 4378 4347 4380
rect 4371 4378 4427 4380
rect 4451 4378 4507 4380
rect 4531 4378 4587 4380
rect 4291 4326 4337 4378
rect 4337 4326 4347 4378
rect 4371 4326 4401 4378
rect 4401 4326 4413 4378
rect 4413 4326 4427 4378
rect 4451 4326 4465 4378
rect 4465 4326 4477 4378
rect 4477 4326 4507 4378
rect 4531 4326 4541 4378
rect 4541 4326 4587 4378
rect 4291 4324 4347 4326
rect 4371 4324 4427 4326
rect 4451 4324 4507 4326
rect 4531 4324 4587 4326
rect 12065 4378 12121 4380
rect 12145 4378 12201 4380
rect 12225 4378 12281 4380
rect 12305 4378 12361 4380
rect 12065 4326 12111 4378
rect 12111 4326 12121 4378
rect 12145 4326 12175 4378
rect 12175 4326 12187 4378
rect 12187 4326 12201 4378
rect 12225 4326 12239 4378
rect 12239 4326 12251 4378
rect 12251 4326 12281 4378
rect 12305 4326 12315 4378
rect 12315 4326 12361 4378
rect 12065 4324 12121 4326
rect 12145 4324 12201 4326
rect 12225 4324 12281 4326
rect 12305 4324 12361 4326
rect 19839 4378 19895 4380
rect 19919 4378 19975 4380
rect 19999 4378 20055 4380
rect 20079 4378 20135 4380
rect 19839 4326 19885 4378
rect 19885 4326 19895 4378
rect 19919 4326 19949 4378
rect 19949 4326 19961 4378
rect 19961 4326 19975 4378
rect 19999 4326 20013 4378
rect 20013 4326 20025 4378
rect 20025 4326 20055 4378
rect 20079 4326 20089 4378
rect 20089 4326 20135 4378
rect 19839 4324 19895 4326
rect 19919 4324 19975 4326
rect 19999 4324 20055 4326
rect 20079 4324 20135 4326
rect 27613 4378 27669 4380
rect 27693 4378 27749 4380
rect 27773 4378 27829 4380
rect 27853 4378 27909 4380
rect 27613 4326 27659 4378
rect 27659 4326 27669 4378
rect 27693 4326 27723 4378
rect 27723 4326 27735 4378
rect 27735 4326 27749 4378
rect 27773 4326 27787 4378
rect 27787 4326 27799 4378
rect 27799 4326 27829 4378
rect 27853 4326 27863 4378
rect 27863 4326 27909 4378
rect 27613 4324 27669 4326
rect 27693 4324 27749 4326
rect 27773 4324 27829 4326
rect 27853 4324 27909 4326
rect 8178 3834 8234 3836
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8178 3782 8224 3834
rect 8224 3782 8234 3834
rect 8258 3782 8288 3834
rect 8288 3782 8300 3834
rect 8300 3782 8314 3834
rect 8338 3782 8352 3834
rect 8352 3782 8364 3834
rect 8364 3782 8394 3834
rect 8418 3782 8428 3834
rect 8428 3782 8474 3834
rect 8178 3780 8234 3782
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 15952 3834 16008 3836
rect 16032 3834 16088 3836
rect 16112 3834 16168 3836
rect 16192 3834 16248 3836
rect 15952 3782 15998 3834
rect 15998 3782 16008 3834
rect 16032 3782 16062 3834
rect 16062 3782 16074 3834
rect 16074 3782 16088 3834
rect 16112 3782 16126 3834
rect 16126 3782 16138 3834
rect 16138 3782 16168 3834
rect 16192 3782 16202 3834
rect 16202 3782 16248 3834
rect 15952 3780 16008 3782
rect 16032 3780 16088 3782
rect 16112 3780 16168 3782
rect 16192 3780 16248 3782
rect 23726 3834 23782 3836
rect 23806 3834 23862 3836
rect 23886 3834 23942 3836
rect 23966 3834 24022 3836
rect 23726 3782 23772 3834
rect 23772 3782 23782 3834
rect 23806 3782 23836 3834
rect 23836 3782 23848 3834
rect 23848 3782 23862 3834
rect 23886 3782 23900 3834
rect 23900 3782 23912 3834
rect 23912 3782 23942 3834
rect 23966 3782 23976 3834
rect 23976 3782 24022 3834
rect 23726 3780 23782 3782
rect 23806 3780 23862 3782
rect 23886 3780 23942 3782
rect 23966 3780 24022 3782
rect 31500 3834 31556 3836
rect 31580 3834 31636 3836
rect 31660 3834 31716 3836
rect 31740 3834 31796 3836
rect 31500 3782 31546 3834
rect 31546 3782 31556 3834
rect 31580 3782 31610 3834
rect 31610 3782 31622 3834
rect 31622 3782 31636 3834
rect 31660 3782 31674 3834
rect 31674 3782 31686 3834
rect 31686 3782 31716 3834
rect 31740 3782 31750 3834
rect 31750 3782 31796 3834
rect 31500 3780 31556 3782
rect 31580 3780 31636 3782
rect 31660 3780 31716 3782
rect 31740 3780 31796 3782
rect 4291 3290 4347 3292
rect 4371 3290 4427 3292
rect 4451 3290 4507 3292
rect 4531 3290 4587 3292
rect 4291 3238 4337 3290
rect 4337 3238 4347 3290
rect 4371 3238 4401 3290
rect 4401 3238 4413 3290
rect 4413 3238 4427 3290
rect 4451 3238 4465 3290
rect 4465 3238 4477 3290
rect 4477 3238 4507 3290
rect 4531 3238 4541 3290
rect 4541 3238 4587 3290
rect 4291 3236 4347 3238
rect 4371 3236 4427 3238
rect 4451 3236 4507 3238
rect 4531 3236 4587 3238
rect 12065 3290 12121 3292
rect 12145 3290 12201 3292
rect 12225 3290 12281 3292
rect 12305 3290 12361 3292
rect 12065 3238 12111 3290
rect 12111 3238 12121 3290
rect 12145 3238 12175 3290
rect 12175 3238 12187 3290
rect 12187 3238 12201 3290
rect 12225 3238 12239 3290
rect 12239 3238 12251 3290
rect 12251 3238 12281 3290
rect 12305 3238 12315 3290
rect 12315 3238 12361 3290
rect 12065 3236 12121 3238
rect 12145 3236 12201 3238
rect 12225 3236 12281 3238
rect 12305 3236 12361 3238
rect 19839 3290 19895 3292
rect 19919 3290 19975 3292
rect 19999 3290 20055 3292
rect 20079 3290 20135 3292
rect 19839 3238 19885 3290
rect 19885 3238 19895 3290
rect 19919 3238 19949 3290
rect 19949 3238 19961 3290
rect 19961 3238 19975 3290
rect 19999 3238 20013 3290
rect 20013 3238 20025 3290
rect 20025 3238 20055 3290
rect 20079 3238 20089 3290
rect 20089 3238 20135 3290
rect 19839 3236 19895 3238
rect 19919 3236 19975 3238
rect 19999 3236 20055 3238
rect 20079 3236 20135 3238
rect 27613 3290 27669 3292
rect 27693 3290 27749 3292
rect 27773 3290 27829 3292
rect 27853 3290 27909 3292
rect 27613 3238 27659 3290
rect 27659 3238 27669 3290
rect 27693 3238 27723 3290
rect 27723 3238 27735 3290
rect 27735 3238 27749 3290
rect 27773 3238 27787 3290
rect 27787 3238 27799 3290
rect 27799 3238 27829 3290
rect 27853 3238 27863 3290
rect 27863 3238 27909 3290
rect 27613 3236 27669 3238
rect 27693 3236 27749 3238
rect 27773 3236 27829 3238
rect 27853 3236 27909 3238
rect 8178 2746 8234 2748
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8178 2694 8224 2746
rect 8224 2694 8234 2746
rect 8258 2694 8288 2746
rect 8288 2694 8300 2746
rect 8300 2694 8314 2746
rect 8338 2694 8352 2746
rect 8352 2694 8364 2746
rect 8364 2694 8394 2746
rect 8418 2694 8428 2746
rect 8428 2694 8474 2746
rect 8178 2692 8234 2694
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 15952 2746 16008 2748
rect 16032 2746 16088 2748
rect 16112 2746 16168 2748
rect 16192 2746 16248 2748
rect 15952 2694 15998 2746
rect 15998 2694 16008 2746
rect 16032 2694 16062 2746
rect 16062 2694 16074 2746
rect 16074 2694 16088 2746
rect 16112 2694 16126 2746
rect 16126 2694 16138 2746
rect 16138 2694 16168 2746
rect 16192 2694 16202 2746
rect 16202 2694 16248 2746
rect 15952 2692 16008 2694
rect 16032 2692 16088 2694
rect 16112 2692 16168 2694
rect 16192 2692 16248 2694
rect 23726 2746 23782 2748
rect 23806 2746 23862 2748
rect 23886 2746 23942 2748
rect 23966 2746 24022 2748
rect 23726 2694 23772 2746
rect 23772 2694 23782 2746
rect 23806 2694 23836 2746
rect 23836 2694 23848 2746
rect 23848 2694 23862 2746
rect 23886 2694 23900 2746
rect 23900 2694 23912 2746
rect 23912 2694 23942 2746
rect 23966 2694 23976 2746
rect 23976 2694 24022 2746
rect 23726 2692 23782 2694
rect 23806 2692 23862 2694
rect 23886 2692 23942 2694
rect 23966 2692 24022 2694
rect 31500 2746 31556 2748
rect 31580 2746 31636 2748
rect 31660 2746 31716 2748
rect 31740 2746 31796 2748
rect 31500 2694 31546 2746
rect 31546 2694 31556 2746
rect 31580 2694 31610 2746
rect 31610 2694 31622 2746
rect 31622 2694 31636 2746
rect 31660 2694 31674 2746
rect 31674 2694 31686 2746
rect 31686 2694 31716 2746
rect 31740 2694 31750 2746
rect 31750 2694 31796 2746
rect 31500 2692 31556 2694
rect 31580 2692 31636 2694
rect 31660 2692 31716 2694
rect 31740 2692 31796 2694
rect 4291 2202 4347 2204
rect 4371 2202 4427 2204
rect 4451 2202 4507 2204
rect 4531 2202 4587 2204
rect 4291 2150 4337 2202
rect 4337 2150 4347 2202
rect 4371 2150 4401 2202
rect 4401 2150 4413 2202
rect 4413 2150 4427 2202
rect 4451 2150 4465 2202
rect 4465 2150 4477 2202
rect 4477 2150 4507 2202
rect 4531 2150 4541 2202
rect 4541 2150 4587 2202
rect 4291 2148 4347 2150
rect 4371 2148 4427 2150
rect 4451 2148 4507 2150
rect 4531 2148 4587 2150
rect 12065 2202 12121 2204
rect 12145 2202 12201 2204
rect 12225 2202 12281 2204
rect 12305 2202 12361 2204
rect 12065 2150 12111 2202
rect 12111 2150 12121 2202
rect 12145 2150 12175 2202
rect 12175 2150 12187 2202
rect 12187 2150 12201 2202
rect 12225 2150 12239 2202
rect 12239 2150 12251 2202
rect 12251 2150 12281 2202
rect 12305 2150 12315 2202
rect 12315 2150 12361 2202
rect 12065 2148 12121 2150
rect 12145 2148 12201 2150
rect 12225 2148 12281 2150
rect 12305 2148 12361 2150
rect 19839 2202 19895 2204
rect 19919 2202 19975 2204
rect 19999 2202 20055 2204
rect 20079 2202 20135 2204
rect 19839 2150 19885 2202
rect 19885 2150 19895 2202
rect 19919 2150 19949 2202
rect 19949 2150 19961 2202
rect 19961 2150 19975 2202
rect 19999 2150 20013 2202
rect 20013 2150 20025 2202
rect 20025 2150 20055 2202
rect 20079 2150 20089 2202
rect 20089 2150 20135 2202
rect 19839 2148 19895 2150
rect 19919 2148 19975 2150
rect 19999 2148 20055 2150
rect 20079 2148 20135 2150
rect 27613 2202 27669 2204
rect 27693 2202 27749 2204
rect 27773 2202 27829 2204
rect 27853 2202 27909 2204
rect 27613 2150 27659 2202
rect 27659 2150 27669 2202
rect 27693 2150 27723 2202
rect 27723 2150 27735 2202
rect 27735 2150 27749 2202
rect 27773 2150 27787 2202
rect 27787 2150 27799 2202
rect 27799 2150 27829 2202
rect 27853 2150 27863 2202
rect 27863 2150 27909 2202
rect 27613 2148 27669 2150
rect 27693 2148 27749 2150
rect 27773 2148 27829 2150
rect 27853 2148 27909 2150
rect 8178 1658 8234 1660
rect 8258 1658 8314 1660
rect 8338 1658 8394 1660
rect 8418 1658 8474 1660
rect 8178 1606 8224 1658
rect 8224 1606 8234 1658
rect 8258 1606 8288 1658
rect 8288 1606 8300 1658
rect 8300 1606 8314 1658
rect 8338 1606 8352 1658
rect 8352 1606 8364 1658
rect 8364 1606 8394 1658
rect 8418 1606 8428 1658
rect 8428 1606 8474 1658
rect 8178 1604 8234 1606
rect 8258 1604 8314 1606
rect 8338 1604 8394 1606
rect 8418 1604 8474 1606
rect 15952 1658 16008 1660
rect 16032 1658 16088 1660
rect 16112 1658 16168 1660
rect 16192 1658 16248 1660
rect 15952 1606 15998 1658
rect 15998 1606 16008 1658
rect 16032 1606 16062 1658
rect 16062 1606 16074 1658
rect 16074 1606 16088 1658
rect 16112 1606 16126 1658
rect 16126 1606 16138 1658
rect 16138 1606 16168 1658
rect 16192 1606 16202 1658
rect 16202 1606 16248 1658
rect 15952 1604 16008 1606
rect 16032 1604 16088 1606
rect 16112 1604 16168 1606
rect 16192 1604 16248 1606
rect 23726 1658 23782 1660
rect 23806 1658 23862 1660
rect 23886 1658 23942 1660
rect 23966 1658 24022 1660
rect 23726 1606 23772 1658
rect 23772 1606 23782 1658
rect 23806 1606 23836 1658
rect 23836 1606 23848 1658
rect 23848 1606 23862 1658
rect 23886 1606 23900 1658
rect 23900 1606 23912 1658
rect 23912 1606 23942 1658
rect 23966 1606 23976 1658
rect 23976 1606 24022 1658
rect 23726 1604 23782 1606
rect 23806 1604 23862 1606
rect 23886 1604 23942 1606
rect 23966 1604 24022 1606
rect 31500 1658 31556 1660
rect 31580 1658 31636 1660
rect 31660 1658 31716 1660
rect 31740 1658 31796 1660
rect 31500 1606 31546 1658
rect 31546 1606 31556 1658
rect 31580 1606 31610 1658
rect 31610 1606 31622 1658
rect 31622 1606 31636 1658
rect 31660 1606 31674 1658
rect 31674 1606 31686 1658
rect 31686 1606 31716 1658
rect 31740 1606 31750 1658
rect 31750 1606 31796 1658
rect 31500 1604 31556 1606
rect 31580 1604 31636 1606
rect 31660 1604 31716 1606
rect 31740 1604 31796 1606
rect 4291 1114 4347 1116
rect 4371 1114 4427 1116
rect 4451 1114 4507 1116
rect 4531 1114 4587 1116
rect 4291 1062 4337 1114
rect 4337 1062 4347 1114
rect 4371 1062 4401 1114
rect 4401 1062 4413 1114
rect 4413 1062 4427 1114
rect 4451 1062 4465 1114
rect 4465 1062 4477 1114
rect 4477 1062 4507 1114
rect 4531 1062 4541 1114
rect 4541 1062 4587 1114
rect 4291 1060 4347 1062
rect 4371 1060 4427 1062
rect 4451 1060 4507 1062
rect 4531 1060 4587 1062
rect 12065 1114 12121 1116
rect 12145 1114 12201 1116
rect 12225 1114 12281 1116
rect 12305 1114 12361 1116
rect 12065 1062 12111 1114
rect 12111 1062 12121 1114
rect 12145 1062 12175 1114
rect 12175 1062 12187 1114
rect 12187 1062 12201 1114
rect 12225 1062 12239 1114
rect 12239 1062 12251 1114
rect 12251 1062 12281 1114
rect 12305 1062 12315 1114
rect 12315 1062 12361 1114
rect 12065 1060 12121 1062
rect 12145 1060 12201 1062
rect 12225 1060 12281 1062
rect 12305 1060 12361 1062
rect 19839 1114 19895 1116
rect 19919 1114 19975 1116
rect 19999 1114 20055 1116
rect 20079 1114 20135 1116
rect 19839 1062 19885 1114
rect 19885 1062 19895 1114
rect 19919 1062 19949 1114
rect 19949 1062 19961 1114
rect 19961 1062 19975 1114
rect 19999 1062 20013 1114
rect 20013 1062 20025 1114
rect 20025 1062 20055 1114
rect 20079 1062 20089 1114
rect 20089 1062 20135 1114
rect 19839 1060 19895 1062
rect 19919 1060 19975 1062
rect 19999 1060 20055 1062
rect 20079 1060 20135 1062
rect 27613 1114 27669 1116
rect 27693 1114 27749 1116
rect 27773 1114 27829 1116
rect 27853 1114 27909 1116
rect 27613 1062 27659 1114
rect 27659 1062 27669 1114
rect 27693 1062 27723 1114
rect 27723 1062 27735 1114
rect 27735 1062 27749 1114
rect 27773 1062 27787 1114
rect 27787 1062 27799 1114
rect 27799 1062 27829 1114
rect 27853 1062 27863 1114
rect 27863 1062 27909 1114
rect 27613 1060 27669 1062
rect 27693 1060 27749 1062
rect 27773 1060 27829 1062
rect 27853 1060 27909 1062
rect 8178 570 8234 572
rect 8258 570 8314 572
rect 8338 570 8394 572
rect 8418 570 8474 572
rect 8178 518 8224 570
rect 8224 518 8234 570
rect 8258 518 8288 570
rect 8288 518 8300 570
rect 8300 518 8314 570
rect 8338 518 8352 570
rect 8352 518 8364 570
rect 8364 518 8394 570
rect 8418 518 8428 570
rect 8428 518 8474 570
rect 8178 516 8234 518
rect 8258 516 8314 518
rect 8338 516 8394 518
rect 8418 516 8474 518
rect 15952 570 16008 572
rect 16032 570 16088 572
rect 16112 570 16168 572
rect 16192 570 16248 572
rect 15952 518 15998 570
rect 15998 518 16008 570
rect 16032 518 16062 570
rect 16062 518 16074 570
rect 16074 518 16088 570
rect 16112 518 16126 570
rect 16126 518 16138 570
rect 16138 518 16168 570
rect 16192 518 16202 570
rect 16202 518 16248 570
rect 15952 516 16008 518
rect 16032 516 16088 518
rect 16112 516 16168 518
rect 16192 516 16248 518
rect 23726 570 23782 572
rect 23806 570 23862 572
rect 23886 570 23942 572
rect 23966 570 24022 572
rect 23726 518 23772 570
rect 23772 518 23782 570
rect 23806 518 23836 570
rect 23836 518 23848 570
rect 23848 518 23862 570
rect 23886 518 23900 570
rect 23900 518 23912 570
rect 23912 518 23942 570
rect 23966 518 23976 570
rect 23976 518 24022 570
rect 23726 516 23782 518
rect 23806 516 23862 518
rect 23886 516 23942 518
rect 23966 516 24022 518
rect 31500 570 31556 572
rect 31580 570 31636 572
rect 31660 570 31716 572
rect 31740 570 31796 572
rect 31500 518 31546 570
rect 31546 518 31556 570
rect 31580 518 31610 570
rect 31610 518 31622 570
rect 31622 518 31636 570
rect 31660 518 31674 570
rect 31674 518 31686 570
rect 31686 518 31716 570
rect 31740 518 31750 570
rect 31750 518 31796 570
rect 31500 516 31556 518
rect 31580 516 31636 518
rect 31660 516 31716 518
rect 31740 516 31796 518
<< metal3 >>
rect 4521 21996 4587 21997
rect 8201 21996 8267 21997
rect 4470 21932 4476 21996
rect 4540 21994 4587 21996
rect 4540 21992 4632 21994
rect 4582 21936 4632 21992
rect 4540 21934 4632 21936
rect 4540 21932 4587 21934
rect 8150 21932 8156 21996
rect 8220 21994 8267 21996
rect 8220 21992 8312 21994
rect 8262 21936 8312 21992
rect 8220 21934 8312 21936
rect 8220 21932 8267 21934
rect 27470 21932 27476 21996
rect 27540 21994 27546 21996
rect 28993 21994 29059 21997
rect 27540 21992 29059 21994
rect 27540 21936 28998 21992
rect 29054 21936 29059 21992
rect 27540 21934 29059 21936
rect 27540 21932 27546 21934
rect 4521 21931 4587 21932
rect 8201 21931 8267 21932
rect 28993 21931 29059 21934
rect 841 21860 907 21861
rect 1577 21860 1643 21861
rect 2313 21860 2379 21861
rect 790 21796 796 21860
rect 860 21858 907 21860
rect 860 21856 952 21858
rect 902 21800 952 21856
rect 860 21798 952 21800
rect 860 21796 907 21798
rect 1526 21796 1532 21860
rect 1596 21858 1643 21860
rect 1596 21856 1688 21858
rect 1638 21800 1688 21856
rect 1596 21798 1688 21800
rect 1596 21796 1643 21798
rect 2262 21796 2268 21860
rect 2332 21858 2379 21860
rect 2332 21856 2424 21858
rect 2374 21800 2424 21856
rect 2332 21798 2424 21800
rect 2332 21796 2379 21798
rect 2998 21796 3004 21860
rect 3068 21858 3074 21860
rect 3233 21858 3299 21861
rect 3785 21860 3851 21861
rect 5257 21860 5323 21861
rect 5993 21860 6059 21861
rect 6729 21860 6795 21861
rect 7465 21860 7531 21861
rect 3068 21856 3299 21858
rect 3068 21800 3238 21856
rect 3294 21800 3299 21856
rect 3068 21798 3299 21800
rect 3068 21796 3074 21798
rect 841 21795 907 21796
rect 1577 21795 1643 21796
rect 2313 21795 2379 21796
rect 3233 21795 3299 21798
rect 3734 21796 3740 21860
rect 3804 21858 3851 21860
rect 3804 21856 3896 21858
rect 3846 21800 3896 21856
rect 3804 21798 3896 21800
rect 3804 21796 3851 21798
rect 5206 21796 5212 21860
rect 5276 21858 5323 21860
rect 5276 21856 5368 21858
rect 5318 21800 5368 21856
rect 5276 21798 5368 21800
rect 5276 21796 5323 21798
rect 5942 21796 5948 21860
rect 6012 21858 6059 21860
rect 6012 21856 6104 21858
rect 6054 21800 6104 21856
rect 6012 21798 6104 21800
rect 6012 21796 6059 21798
rect 6678 21796 6684 21860
rect 6748 21858 6795 21860
rect 6748 21856 6840 21858
rect 6790 21800 6840 21856
rect 6748 21798 6840 21800
rect 6748 21796 6795 21798
rect 7414 21796 7420 21860
rect 7484 21858 7531 21860
rect 8753 21858 8819 21861
rect 9673 21860 9739 21861
rect 10409 21860 10475 21861
rect 11145 21860 11211 21861
rect 25865 21860 25931 21861
rect 8886 21858 8892 21860
rect 7484 21856 7576 21858
rect 7526 21800 7576 21856
rect 7484 21798 7576 21800
rect 8753 21856 8892 21858
rect 8753 21800 8758 21856
rect 8814 21800 8892 21856
rect 8753 21798 8892 21800
rect 7484 21796 7531 21798
rect 3785 21795 3851 21796
rect 5257 21795 5323 21796
rect 5993 21795 6059 21796
rect 6729 21795 6795 21796
rect 7465 21795 7531 21796
rect 8753 21795 8819 21798
rect 8886 21796 8892 21798
rect 8956 21796 8962 21860
rect 9622 21796 9628 21860
rect 9692 21858 9739 21860
rect 9692 21856 9784 21858
rect 9734 21800 9784 21856
rect 9692 21798 9784 21800
rect 9692 21796 9739 21798
rect 10358 21796 10364 21860
rect 10428 21858 10475 21860
rect 10428 21856 10520 21858
rect 10470 21800 10520 21856
rect 10428 21798 10520 21800
rect 10428 21796 10475 21798
rect 11094 21796 11100 21860
rect 11164 21858 11211 21860
rect 25814 21858 25820 21860
rect 11164 21856 11256 21858
rect 11206 21800 11256 21856
rect 11164 21798 11256 21800
rect 25774 21798 25820 21858
rect 25884 21856 25931 21860
rect 25926 21800 25931 21856
rect 11164 21796 11211 21798
rect 25814 21796 25820 21798
rect 25884 21796 25931 21800
rect 26550 21796 26556 21860
rect 26620 21858 26626 21860
rect 26785 21858 26851 21861
rect 26620 21856 26851 21858
rect 26620 21800 26790 21856
rect 26846 21800 26851 21856
rect 26620 21798 26851 21800
rect 26620 21796 26626 21798
rect 9673 21795 9739 21796
rect 10409 21795 10475 21796
rect 11145 21795 11211 21796
rect 25865 21795 25931 21796
rect 26785 21795 26851 21798
rect 28022 21796 28028 21860
rect 28092 21858 28098 21860
rect 28533 21858 28599 21861
rect 28092 21856 28599 21858
rect 28092 21800 28538 21856
rect 28594 21800 28599 21856
rect 28092 21798 28599 21800
rect 28092 21796 28098 21798
rect 28533 21795 28599 21798
rect 29494 21796 29500 21860
rect 29564 21858 29570 21860
rect 30005 21858 30071 21861
rect 29564 21856 30071 21858
rect 29564 21800 30010 21856
rect 30066 21800 30071 21856
rect 29564 21798 30071 21800
rect 29564 21796 29570 21798
rect 30005 21795 30071 21798
rect 4281 21792 4597 21793
rect 4281 21728 4287 21792
rect 4351 21728 4367 21792
rect 4431 21728 4447 21792
rect 4511 21728 4527 21792
rect 4591 21728 4597 21792
rect 4281 21727 4597 21728
rect 12055 21792 12371 21793
rect 12055 21728 12061 21792
rect 12125 21728 12141 21792
rect 12205 21728 12221 21792
rect 12285 21728 12301 21792
rect 12365 21728 12371 21792
rect 12055 21727 12371 21728
rect 19829 21792 20145 21793
rect 19829 21728 19835 21792
rect 19899 21728 19915 21792
rect 19979 21728 19995 21792
rect 20059 21728 20075 21792
rect 20139 21728 20145 21792
rect 19829 21727 20145 21728
rect 27603 21792 27919 21793
rect 27603 21728 27609 21792
rect 27673 21728 27689 21792
rect 27753 21728 27769 21792
rect 27833 21728 27849 21792
rect 27913 21728 27919 21792
rect 27603 21727 27919 21728
rect 28758 21660 28764 21724
rect 28828 21722 28834 21724
rect 29545 21722 29611 21725
rect 28828 21720 29611 21722
rect 28828 21664 29550 21720
rect 29606 21664 29611 21720
rect 28828 21662 29611 21664
rect 28828 21660 28834 21662
rect 29545 21659 29611 21662
rect 11881 21588 11947 21589
rect 13353 21588 13419 21589
rect 11830 21524 11836 21588
rect 11900 21586 11947 21588
rect 13302 21586 13308 21588
rect 11900 21584 11992 21586
rect 11942 21528 11992 21584
rect 11900 21526 11992 21528
rect 13262 21526 13308 21586
rect 13372 21584 13419 21588
rect 13414 21528 13419 21584
rect 11900 21524 11947 21526
rect 13302 21524 13308 21526
rect 13372 21524 13419 21528
rect 11881 21523 11947 21524
rect 13353 21523 13419 21524
rect 16982 21252 16988 21316
rect 17052 21314 17058 21316
rect 17125 21314 17191 21317
rect 17052 21312 17191 21314
rect 17052 21256 17130 21312
rect 17186 21256 17191 21312
rect 17052 21254 17191 21256
rect 17052 21252 17058 21254
rect 17125 21251 17191 21254
rect 8168 21248 8484 21249
rect 8168 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8484 21248
rect 8168 21183 8484 21184
rect 15942 21248 16258 21249
rect 15942 21184 15948 21248
rect 16012 21184 16028 21248
rect 16092 21184 16108 21248
rect 16172 21184 16188 21248
rect 16252 21184 16258 21248
rect 15942 21183 16258 21184
rect 23716 21248 24032 21249
rect 23716 21184 23722 21248
rect 23786 21184 23802 21248
rect 23866 21184 23882 21248
rect 23946 21184 23962 21248
rect 24026 21184 24032 21248
rect 23716 21183 24032 21184
rect 31490 21248 31806 21249
rect 31490 21184 31496 21248
rect 31560 21184 31576 21248
rect 31640 21184 31656 21248
rect 31720 21184 31736 21248
rect 31800 21184 31806 21248
rect 31490 21183 31806 21184
rect 14038 20708 14044 20772
rect 14108 20770 14114 20772
rect 14641 20770 14707 20773
rect 14108 20768 14707 20770
rect 14108 20712 14646 20768
rect 14702 20712 14707 20768
rect 14108 20710 14707 20712
rect 14108 20708 14114 20710
rect 14641 20707 14707 20710
rect 4281 20704 4597 20705
rect 4281 20640 4287 20704
rect 4351 20640 4367 20704
rect 4431 20640 4447 20704
rect 4511 20640 4527 20704
rect 4591 20640 4597 20704
rect 4281 20639 4597 20640
rect 12055 20704 12371 20705
rect 12055 20640 12061 20704
rect 12125 20640 12141 20704
rect 12205 20640 12221 20704
rect 12285 20640 12301 20704
rect 12365 20640 12371 20704
rect 12055 20639 12371 20640
rect 19829 20704 20145 20705
rect 19829 20640 19835 20704
rect 19899 20640 19915 20704
rect 19979 20640 19995 20704
rect 20059 20640 20075 20704
rect 20139 20640 20145 20704
rect 19829 20639 20145 20640
rect 27603 20704 27919 20705
rect 27603 20640 27609 20704
rect 27673 20640 27689 20704
rect 27753 20640 27769 20704
rect 27833 20640 27849 20704
rect 27913 20640 27919 20704
rect 27603 20639 27919 20640
rect 12934 20436 12940 20500
rect 13004 20498 13010 20500
rect 14089 20498 14155 20501
rect 13004 20496 14155 20498
rect 13004 20440 14094 20496
rect 14150 20440 14155 20496
rect 13004 20438 14155 20440
rect 13004 20436 13010 20438
rect 14089 20435 14155 20438
rect 15285 20498 15351 20501
rect 24485 20498 24551 20501
rect 15285 20496 24551 20498
rect 15285 20440 15290 20496
rect 15346 20440 24490 20496
rect 24546 20440 24551 20496
rect 15285 20438 24551 20440
rect 15285 20435 15351 20438
rect 24485 20435 24551 20438
rect 27153 20498 27219 20501
rect 27521 20498 27587 20501
rect 27153 20496 27587 20498
rect 27153 20440 27158 20496
rect 27214 20440 27526 20496
rect 27582 20440 27587 20496
rect 27153 20438 27587 20440
rect 27153 20435 27219 20438
rect 27521 20435 27587 20438
rect 17309 20362 17375 20365
rect 20253 20362 20319 20365
rect 21081 20362 21147 20365
rect 28625 20362 28691 20365
rect 17309 20360 21147 20362
rect 17309 20304 17314 20360
rect 17370 20304 20258 20360
rect 20314 20304 21086 20360
rect 21142 20304 21147 20360
rect 17309 20302 21147 20304
rect 17309 20299 17375 20302
rect 20253 20299 20319 20302
rect 21081 20299 21147 20302
rect 23062 20360 28691 20362
rect 23062 20304 28630 20360
rect 28686 20304 28691 20360
rect 23062 20302 28691 20304
rect 17953 20226 18019 20229
rect 19149 20226 19215 20229
rect 22829 20226 22895 20229
rect 17953 20224 22895 20226
rect 17953 20168 17958 20224
rect 18014 20168 19154 20224
rect 19210 20168 22834 20224
rect 22890 20168 22895 20224
rect 17953 20166 22895 20168
rect 17953 20163 18019 20166
rect 19149 20163 19215 20166
rect 22829 20163 22895 20166
rect 8168 20160 8484 20161
rect 8168 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8484 20160
rect 8168 20095 8484 20096
rect 15942 20160 16258 20161
rect 15942 20096 15948 20160
rect 16012 20096 16028 20160
rect 16092 20096 16108 20160
rect 16172 20096 16188 20160
rect 16252 20096 16258 20160
rect 15942 20095 16258 20096
rect 19977 20090 20043 20093
rect 23062 20090 23122 20302
rect 28625 20299 28691 20302
rect 23716 20160 24032 20161
rect 23716 20096 23722 20160
rect 23786 20096 23802 20160
rect 23866 20096 23882 20160
rect 23946 20096 23962 20160
rect 24026 20096 24032 20160
rect 23716 20095 24032 20096
rect 31490 20160 31806 20161
rect 31490 20096 31496 20160
rect 31560 20096 31576 20160
rect 31640 20096 31656 20160
rect 31720 20096 31736 20160
rect 31800 20096 31806 20160
rect 31490 20095 31806 20096
rect 19977 20088 23122 20090
rect 19977 20032 19982 20088
rect 20038 20032 23122 20088
rect 19977 20030 23122 20032
rect 19977 20027 20043 20030
rect 9213 19954 9279 19957
rect 13537 19954 13603 19957
rect 9213 19952 13603 19954
rect 9213 19896 9218 19952
rect 9274 19896 13542 19952
rect 13598 19896 13603 19952
rect 9213 19894 13603 19896
rect 9213 19891 9279 19894
rect 13537 19891 13603 19894
rect 13721 19954 13787 19957
rect 14825 19954 14891 19957
rect 13721 19952 14891 19954
rect 13721 19896 13726 19952
rect 13782 19896 14830 19952
rect 14886 19896 14891 19952
rect 13721 19894 14891 19896
rect 13721 19891 13787 19894
rect 14825 19891 14891 19894
rect 15101 19954 15167 19957
rect 20069 19954 20135 19957
rect 24853 19954 24919 19957
rect 15101 19952 20135 19954
rect 15101 19896 15106 19952
rect 15162 19896 20074 19952
rect 20130 19896 20135 19952
rect 15101 19894 20135 19896
rect 15101 19891 15167 19894
rect 20069 19891 20135 19894
rect 20302 19952 24919 19954
rect 20302 19896 24858 19952
rect 24914 19896 24919 19952
rect 20302 19894 24919 19896
rect 8937 19818 9003 19821
rect 13261 19818 13327 19821
rect 8937 19816 13327 19818
rect 8937 19760 8942 19816
rect 8998 19760 13266 19816
rect 13322 19760 13327 19816
rect 8937 19758 13327 19760
rect 8937 19755 9003 19758
rect 13261 19755 13327 19758
rect 14273 19818 14339 19821
rect 20302 19818 20362 19894
rect 24853 19891 24919 19894
rect 14273 19816 20362 19818
rect 14273 19760 14278 19816
rect 14334 19760 20362 19816
rect 14273 19758 20362 19760
rect 14273 19755 14339 19758
rect 4281 19616 4597 19617
rect 4281 19552 4287 19616
rect 4351 19552 4367 19616
rect 4431 19552 4447 19616
rect 4511 19552 4527 19616
rect 4591 19552 4597 19616
rect 4281 19551 4597 19552
rect 12055 19616 12371 19617
rect 12055 19552 12061 19616
rect 12125 19552 12141 19616
rect 12205 19552 12221 19616
rect 12285 19552 12301 19616
rect 12365 19552 12371 19616
rect 12055 19551 12371 19552
rect 19829 19616 20145 19617
rect 19829 19552 19835 19616
rect 19899 19552 19915 19616
rect 19979 19552 19995 19616
rect 20059 19552 20075 19616
rect 20139 19552 20145 19616
rect 19829 19551 20145 19552
rect 27603 19616 27919 19617
rect 27603 19552 27609 19616
rect 27673 19552 27689 19616
rect 27753 19552 27769 19616
rect 27833 19552 27849 19616
rect 27913 19552 27919 19616
rect 27603 19551 27919 19552
rect 16481 19410 16547 19413
rect 23749 19410 23815 19413
rect 16481 19408 23815 19410
rect 16481 19352 16486 19408
rect 16542 19352 23754 19408
rect 23810 19352 23815 19408
rect 16481 19350 23815 19352
rect 16481 19347 16547 19350
rect 23749 19347 23815 19350
rect 8753 19274 8819 19277
rect 9857 19274 9923 19277
rect 8753 19272 9923 19274
rect 8753 19216 8758 19272
rect 8814 19216 9862 19272
rect 9918 19216 9923 19272
rect 8753 19214 9923 19216
rect 8753 19211 8819 19214
rect 9857 19211 9923 19214
rect 20345 19274 20411 19277
rect 20989 19274 21055 19277
rect 20345 19272 21055 19274
rect 20345 19216 20350 19272
rect 20406 19216 20994 19272
rect 21050 19216 21055 19272
rect 20345 19214 21055 19216
rect 20345 19211 20411 19214
rect 20989 19211 21055 19214
rect 29085 19274 29151 19277
rect 29545 19274 29611 19277
rect 29085 19272 29611 19274
rect 29085 19216 29090 19272
rect 29146 19216 29550 19272
rect 29606 19216 29611 19272
rect 29085 19214 29611 19216
rect 29085 19211 29151 19214
rect 29545 19211 29611 19214
rect 9305 19138 9371 19141
rect 9949 19138 10015 19141
rect 15561 19140 15627 19141
rect 9305 19136 10015 19138
rect 9305 19080 9310 19136
rect 9366 19080 9954 19136
rect 10010 19080 10015 19136
rect 9305 19078 10015 19080
rect 9305 19075 9371 19078
rect 9949 19075 10015 19078
rect 15510 19076 15516 19140
rect 15580 19138 15627 19140
rect 15580 19136 15672 19138
rect 15622 19080 15672 19136
rect 15580 19078 15672 19080
rect 15580 19076 15627 19078
rect 15561 19075 15627 19076
rect 8168 19072 8484 19073
rect 8168 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8484 19072
rect 8168 19007 8484 19008
rect 15942 19072 16258 19073
rect 15942 19008 15948 19072
rect 16012 19008 16028 19072
rect 16092 19008 16108 19072
rect 16172 19008 16188 19072
rect 16252 19008 16258 19072
rect 15942 19007 16258 19008
rect 23716 19072 24032 19073
rect 23716 19008 23722 19072
rect 23786 19008 23802 19072
rect 23866 19008 23882 19072
rect 23946 19008 23962 19072
rect 24026 19008 24032 19072
rect 23716 19007 24032 19008
rect 31490 19072 31806 19073
rect 31490 19008 31496 19072
rect 31560 19008 31576 19072
rect 31640 19008 31656 19072
rect 31720 19008 31736 19072
rect 31800 19008 31806 19072
rect 31490 19007 31806 19008
rect 5625 19002 5691 19005
rect 6453 19002 6519 19005
rect 5625 19000 6519 19002
rect 5625 18944 5630 19000
rect 5686 18944 6458 19000
rect 6514 18944 6519 19000
rect 5625 18942 6519 18944
rect 5625 18939 5691 18942
rect 6453 18939 6519 18942
rect 9213 19002 9279 19005
rect 9581 19002 9647 19005
rect 9213 19000 9647 19002
rect 9213 18944 9218 19000
rect 9274 18944 9586 19000
rect 9642 18944 9647 19000
rect 9213 18942 9647 18944
rect 9213 18939 9279 18942
rect 9581 18939 9647 18942
rect 5349 18866 5415 18869
rect 6545 18866 6611 18869
rect 5349 18864 6611 18866
rect 5349 18808 5354 18864
rect 5410 18808 6550 18864
rect 6606 18808 6611 18864
rect 5349 18806 6611 18808
rect 5349 18803 5415 18806
rect 6545 18803 6611 18806
rect 6821 18866 6887 18869
rect 15193 18866 15259 18869
rect 6821 18864 15259 18866
rect 6821 18808 6826 18864
rect 6882 18808 15198 18864
rect 15254 18808 15259 18864
rect 6821 18806 15259 18808
rect 6821 18803 6887 18806
rect 15193 18803 15259 18806
rect 19517 18866 19583 18869
rect 20529 18866 20595 18869
rect 19517 18864 20595 18866
rect 19517 18808 19522 18864
rect 19578 18808 20534 18864
rect 20590 18808 20595 18864
rect 19517 18806 20595 18808
rect 19517 18803 19583 18806
rect 20529 18803 20595 18806
rect 4981 18730 5047 18733
rect 6821 18730 6887 18733
rect 4981 18728 6887 18730
rect 4981 18672 4986 18728
rect 5042 18672 6826 18728
rect 6882 18672 6887 18728
rect 4981 18670 6887 18672
rect 4981 18667 5047 18670
rect 6821 18667 6887 18670
rect 8477 18730 8543 18733
rect 11145 18730 11211 18733
rect 8477 18728 11211 18730
rect 8477 18672 8482 18728
rect 8538 18672 11150 18728
rect 11206 18672 11211 18728
rect 8477 18670 11211 18672
rect 8477 18667 8543 18670
rect 11145 18667 11211 18670
rect 19517 18730 19583 18733
rect 23565 18730 23631 18733
rect 19517 18728 23631 18730
rect 19517 18672 19522 18728
rect 19578 18672 23570 18728
rect 23626 18672 23631 18728
rect 19517 18670 23631 18672
rect 19517 18667 19583 18670
rect 23565 18667 23631 18670
rect 4281 18528 4597 18529
rect 4281 18464 4287 18528
rect 4351 18464 4367 18528
rect 4431 18464 4447 18528
rect 4511 18464 4527 18528
rect 4591 18464 4597 18528
rect 4281 18463 4597 18464
rect 12055 18528 12371 18529
rect 12055 18464 12061 18528
rect 12125 18464 12141 18528
rect 12205 18464 12221 18528
rect 12285 18464 12301 18528
rect 12365 18464 12371 18528
rect 12055 18463 12371 18464
rect 19829 18528 20145 18529
rect 19829 18464 19835 18528
rect 19899 18464 19915 18528
rect 19979 18464 19995 18528
rect 20059 18464 20075 18528
rect 20139 18464 20145 18528
rect 19829 18463 20145 18464
rect 27603 18528 27919 18529
rect 27603 18464 27609 18528
rect 27673 18464 27689 18528
rect 27753 18464 27769 18528
rect 27833 18464 27849 18528
rect 27913 18464 27919 18528
rect 27603 18463 27919 18464
rect 19333 18322 19399 18325
rect 20253 18322 20319 18325
rect 19333 18320 20319 18322
rect 19333 18264 19338 18320
rect 19394 18264 20258 18320
rect 20314 18264 20319 18320
rect 19333 18262 20319 18264
rect 19333 18259 19399 18262
rect 20253 18259 20319 18262
rect 22645 18322 22711 18325
rect 23565 18322 23631 18325
rect 22645 18320 23631 18322
rect 22645 18264 22650 18320
rect 22706 18264 23570 18320
rect 23626 18264 23631 18320
rect 22645 18262 23631 18264
rect 22645 18259 22711 18262
rect 23565 18259 23631 18262
rect 19517 18186 19583 18189
rect 24485 18186 24551 18189
rect 19517 18184 24551 18186
rect 19517 18128 19522 18184
rect 19578 18128 24490 18184
rect 24546 18128 24551 18184
rect 19517 18126 24551 18128
rect 19517 18123 19583 18126
rect 24485 18123 24551 18126
rect 8168 17984 8484 17985
rect 8168 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8484 17984
rect 8168 17919 8484 17920
rect 15942 17984 16258 17985
rect 15942 17920 15948 17984
rect 16012 17920 16028 17984
rect 16092 17920 16108 17984
rect 16172 17920 16188 17984
rect 16252 17920 16258 17984
rect 15942 17919 16258 17920
rect 23716 17984 24032 17985
rect 23716 17920 23722 17984
rect 23786 17920 23802 17984
rect 23866 17920 23882 17984
rect 23946 17920 23962 17984
rect 24026 17920 24032 17984
rect 23716 17919 24032 17920
rect 31490 17984 31806 17985
rect 31490 17920 31496 17984
rect 31560 17920 31576 17984
rect 31640 17920 31656 17984
rect 31720 17920 31736 17984
rect 31800 17920 31806 17984
rect 31490 17919 31806 17920
rect 14733 17916 14799 17917
rect 14733 17912 14780 17916
rect 14844 17914 14850 17916
rect 14733 17856 14738 17912
rect 14733 17852 14780 17856
rect 14844 17854 14890 17914
rect 14844 17852 14850 17854
rect 16430 17852 16436 17916
rect 16500 17914 16506 17916
rect 16573 17914 16639 17917
rect 16500 17912 16639 17914
rect 16500 17856 16578 17912
rect 16634 17856 16639 17912
rect 16500 17854 16639 17856
rect 16500 17852 16506 17854
rect 14733 17851 14799 17852
rect 16573 17851 16639 17854
rect 11329 17778 11395 17781
rect 26325 17778 26391 17781
rect 11329 17776 26391 17778
rect 11329 17720 11334 17776
rect 11390 17720 26330 17776
rect 26386 17720 26391 17776
rect 11329 17718 26391 17720
rect 11329 17715 11395 17718
rect 26325 17715 26391 17718
rect 9581 17642 9647 17645
rect 11697 17642 11763 17645
rect 9581 17640 11763 17642
rect 9581 17584 9586 17640
rect 9642 17584 11702 17640
rect 11758 17584 11763 17640
rect 9581 17582 11763 17584
rect 9581 17579 9647 17582
rect 11697 17579 11763 17582
rect 4281 17440 4597 17441
rect 4281 17376 4287 17440
rect 4351 17376 4367 17440
rect 4431 17376 4447 17440
rect 4511 17376 4527 17440
rect 4591 17376 4597 17440
rect 4281 17375 4597 17376
rect 12055 17440 12371 17441
rect 12055 17376 12061 17440
rect 12125 17376 12141 17440
rect 12205 17376 12221 17440
rect 12285 17376 12301 17440
rect 12365 17376 12371 17440
rect 12055 17375 12371 17376
rect 19829 17440 20145 17441
rect 19829 17376 19835 17440
rect 19899 17376 19915 17440
rect 19979 17376 19995 17440
rect 20059 17376 20075 17440
rect 20139 17376 20145 17440
rect 19829 17375 20145 17376
rect 27603 17440 27919 17441
rect 27603 17376 27609 17440
rect 27673 17376 27689 17440
rect 27753 17376 27769 17440
rect 27833 17376 27849 17440
rect 27913 17376 27919 17440
rect 27603 17375 27919 17376
rect 18321 17370 18387 17373
rect 19241 17370 19307 17373
rect 18321 17368 19307 17370
rect 18321 17312 18326 17368
rect 18382 17312 19246 17368
rect 19302 17312 19307 17368
rect 18321 17310 19307 17312
rect 18321 17307 18387 17310
rect 19241 17307 19307 17310
rect 18965 17098 19031 17101
rect 31017 17098 31083 17101
rect 18965 17096 31083 17098
rect 18965 17040 18970 17096
rect 19026 17040 31022 17096
rect 31078 17040 31083 17096
rect 18965 17038 31083 17040
rect 18965 17035 19031 17038
rect 31017 17035 31083 17038
rect 18137 16962 18203 16965
rect 18781 16962 18847 16965
rect 18137 16960 18847 16962
rect 18137 16904 18142 16960
rect 18198 16904 18786 16960
rect 18842 16904 18847 16960
rect 18137 16902 18847 16904
rect 18137 16899 18203 16902
rect 18781 16899 18847 16902
rect 8168 16896 8484 16897
rect 8168 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8484 16896
rect 8168 16831 8484 16832
rect 15942 16896 16258 16897
rect 15942 16832 15948 16896
rect 16012 16832 16028 16896
rect 16092 16832 16108 16896
rect 16172 16832 16188 16896
rect 16252 16832 16258 16896
rect 15942 16831 16258 16832
rect 23716 16896 24032 16897
rect 23716 16832 23722 16896
rect 23786 16832 23802 16896
rect 23866 16832 23882 16896
rect 23946 16832 23962 16896
rect 24026 16832 24032 16896
rect 23716 16831 24032 16832
rect 31490 16896 31806 16897
rect 31490 16832 31496 16896
rect 31560 16832 31576 16896
rect 31640 16832 31656 16896
rect 31720 16832 31736 16896
rect 31800 16832 31806 16896
rect 31490 16831 31806 16832
rect 18137 16690 18203 16693
rect 31293 16690 31359 16693
rect 18137 16688 31359 16690
rect 18137 16632 18142 16688
rect 18198 16632 31298 16688
rect 31354 16632 31359 16688
rect 18137 16630 31359 16632
rect 18137 16627 18203 16630
rect 31293 16627 31359 16630
rect 17718 16492 17724 16556
rect 17788 16554 17794 16556
rect 18505 16554 18571 16557
rect 17788 16552 18571 16554
rect 17788 16496 18510 16552
rect 18566 16496 18571 16552
rect 17788 16494 18571 16496
rect 17788 16492 17794 16494
rect 18505 16491 18571 16494
rect 23197 16554 23263 16557
rect 25681 16554 25747 16557
rect 23197 16552 25747 16554
rect 23197 16496 23202 16552
rect 23258 16496 25686 16552
rect 25742 16496 25747 16552
rect 23197 16494 25747 16496
rect 23197 16491 23263 16494
rect 25681 16491 25747 16494
rect 4281 16352 4597 16353
rect 4281 16288 4287 16352
rect 4351 16288 4367 16352
rect 4431 16288 4447 16352
rect 4511 16288 4527 16352
rect 4591 16288 4597 16352
rect 4281 16287 4597 16288
rect 12055 16352 12371 16353
rect 12055 16288 12061 16352
rect 12125 16288 12141 16352
rect 12205 16288 12221 16352
rect 12285 16288 12301 16352
rect 12365 16288 12371 16352
rect 12055 16287 12371 16288
rect 19829 16352 20145 16353
rect 19829 16288 19835 16352
rect 19899 16288 19915 16352
rect 19979 16288 19995 16352
rect 20059 16288 20075 16352
rect 20139 16288 20145 16352
rect 19829 16287 20145 16288
rect 27603 16352 27919 16353
rect 27603 16288 27609 16352
rect 27673 16288 27689 16352
rect 27753 16288 27769 16352
rect 27833 16288 27849 16352
rect 27913 16288 27919 16352
rect 27603 16287 27919 16288
rect 13445 16146 13511 16149
rect 23473 16146 23539 16149
rect 13445 16144 23539 16146
rect 13445 16088 13450 16144
rect 13506 16088 23478 16144
rect 23534 16088 23539 16144
rect 13445 16086 23539 16088
rect 13445 16083 13511 16086
rect 23473 16083 23539 16086
rect 24025 16146 24091 16149
rect 26325 16146 26391 16149
rect 24025 16144 26391 16146
rect 24025 16088 24030 16144
rect 24086 16088 26330 16144
rect 26386 16088 26391 16144
rect 24025 16086 26391 16088
rect 24025 16083 24091 16086
rect 26325 16083 26391 16086
rect 15101 16010 15167 16013
rect 17493 16010 17559 16013
rect 15101 16008 17559 16010
rect 15101 15952 15106 16008
rect 15162 15952 17498 16008
rect 17554 15952 17559 16008
rect 15101 15950 17559 15952
rect 15101 15947 15167 15950
rect 17493 15947 17559 15950
rect 20069 16010 20135 16013
rect 22369 16010 22435 16013
rect 20069 16008 22435 16010
rect 20069 15952 20074 16008
rect 20130 15952 22374 16008
rect 22430 15952 22435 16008
rect 20069 15950 22435 15952
rect 20069 15947 20135 15950
rect 22369 15947 22435 15950
rect 8168 15808 8484 15809
rect 8168 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8484 15808
rect 8168 15743 8484 15744
rect 15942 15808 16258 15809
rect 15942 15744 15948 15808
rect 16012 15744 16028 15808
rect 16092 15744 16108 15808
rect 16172 15744 16188 15808
rect 16252 15744 16258 15808
rect 15942 15743 16258 15744
rect 23716 15808 24032 15809
rect 23716 15744 23722 15808
rect 23786 15744 23802 15808
rect 23866 15744 23882 15808
rect 23946 15744 23962 15808
rect 24026 15744 24032 15808
rect 23716 15743 24032 15744
rect 31490 15808 31806 15809
rect 31490 15744 31496 15808
rect 31560 15744 31576 15808
rect 31640 15744 31656 15808
rect 31720 15744 31736 15808
rect 31800 15744 31806 15808
rect 31490 15743 31806 15744
rect 4281 15264 4597 15265
rect 4281 15200 4287 15264
rect 4351 15200 4367 15264
rect 4431 15200 4447 15264
rect 4511 15200 4527 15264
rect 4591 15200 4597 15264
rect 4281 15199 4597 15200
rect 12055 15264 12371 15265
rect 12055 15200 12061 15264
rect 12125 15200 12141 15264
rect 12205 15200 12221 15264
rect 12285 15200 12301 15264
rect 12365 15200 12371 15264
rect 12055 15199 12371 15200
rect 19829 15264 20145 15265
rect 19829 15200 19835 15264
rect 19899 15200 19915 15264
rect 19979 15200 19995 15264
rect 20059 15200 20075 15264
rect 20139 15200 20145 15264
rect 19829 15199 20145 15200
rect 27603 15264 27919 15265
rect 27603 15200 27609 15264
rect 27673 15200 27689 15264
rect 27753 15200 27769 15264
rect 27833 15200 27849 15264
rect 27913 15200 27919 15264
rect 27603 15199 27919 15200
rect 6821 14922 6887 14925
rect 13629 14922 13695 14925
rect 6821 14920 13695 14922
rect 6821 14864 6826 14920
rect 6882 14864 13634 14920
rect 13690 14864 13695 14920
rect 6821 14862 13695 14864
rect 6821 14859 6887 14862
rect 13629 14859 13695 14862
rect 8168 14720 8484 14721
rect 8168 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8484 14720
rect 8168 14655 8484 14656
rect 15942 14720 16258 14721
rect 15942 14656 15948 14720
rect 16012 14656 16028 14720
rect 16092 14656 16108 14720
rect 16172 14656 16188 14720
rect 16252 14656 16258 14720
rect 15942 14655 16258 14656
rect 23716 14720 24032 14721
rect 23716 14656 23722 14720
rect 23786 14656 23802 14720
rect 23866 14656 23882 14720
rect 23946 14656 23962 14720
rect 24026 14656 24032 14720
rect 23716 14655 24032 14656
rect 31490 14720 31806 14721
rect 31490 14656 31496 14720
rect 31560 14656 31576 14720
rect 31640 14656 31656 14720
rect 31720 14656 31736 14720
rect 31800 14656 31806 14720
rect 31490 14655 31806 14656
rect 7189 14378 7255 14381
rect 11513 14378 11579 14381
rect 7189 14376 11579 14378
rect 7189 14320 7194 14376
rect 7250 14320 11518 14376
rect 11574 14320 11579 14376
rect 7189 14318 11579 14320
rect 7189 14315 7255 14318
rect 11513 14315 11579 14318
rect 4281 14176 4597 14177
rect 4281 14112 4287 14176
rect 4351 14112 4367 14176
rect 4431 14112 4447 14176
rect 4511 14112 4527 14176
rect 4591 14112 4597 14176
rect 4281 14111 4597 14112
rect 12055 14176 12371 14177
rect 12055 14112 12061 14176
rect 12125 14112 12141 14176
rect 12205 14112 12221 14176
rect 12285 14112 12301 14176
rect 12365 14112 12371 14176
rect 12055 14111 12371 14112
rect 19829 14176 20145 14177
rect 19829 14112 19835 14176
rect 19899 14112 19915 14176
rect 19979 14112 19995 14176
rect 20059 14112 20075 14176
rect 20139 14112 20145 14176
rect 19829 14111 20145 14112
rect 27603 14176 27919 14177
rect 27603 14112 27609 14176
rect 27673 14112 27689 14176
rect 27753 14112 27769 14176
rect 27833 14112 27849 14176
rect 27913 14112 27919 14176
rect 27603 14111 27919 14112
rect 8168 13632 8484 13633
rect 8168 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8484 13632
rect 8168 13567 8484 13568
rect 15942 13632 16258 13633
rect 15942 13568 15948 13632
rect 16012 13568 16028 13632
rect 16092 13568 16108 13632
rect 16172 13568 16188 13632
rect 16252 13568 16258 13632
rect 15942 13567 16258 13568
rect 23716 13632 24032 13633
rect 23716 13568 23722 13632
rect 23786 13568 23802 13632
rect 23866 13568 23882 13632
rect 23946 13568 23962 13632
rect 24026 13568 24032 13632
rect 23716 13567 24032 13568
rect 31490 13632 31806 13633
rect 31490 13568 31496 13632
rect 31560 13568 31576 13632
rect 31640 13568 31656 13632
rect 31720 13568 31736 13632
rect 31800 13568 31806 13632
rect 31490 13567 31806 13568
rect 4281 13088 4597 13089
rect 4281 13024 4287 13088
rect 4351 13024 4367 13088
rect 4431 13024 4447 13088
rect 4511 13024 4527 13088
rect 4591 13024 4597 13088
rect 4281 13023 4597 13024
rect 12055 13088 12371 13089
rect 12055 13024 12061 13088
rect 12125 13024 12141 13088
rect 12205 13024 12221 13088
rect 12285 13024 12301 13088
rect 12365 13024 12371 13088
rect 12055 13023 12371 13024
rect 19829 13088 20145 13089
rect 19829 13024 19835 13088
rect 19899 13024 19915 13088
rect 19979 13024 19995 13088
rect 20059 13024 20075 13088
rect 20139 13024 20145 13088
rect 19829 13023 20145 13024
rect 27603 13088 27919 13089
rect 27603 13024 27609 13088
rect 27673 13024 27689 13088
rect 27753 13024 27769 13088
rect 27833 13024 27849 13088
rect 27913 13024 27919 13088
rect 27603 13023 27919 13024
rect 8168 12544 8484 12545
rect 8168 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8484 12544
rect 8168 12479 8484 12480
rect 15942 12544 16258 12545
rect 15942 12480 15948 12544
rect 16012 12480 16028 12544
rect 16092 12480 16108 12544
rect 16172 12480 16188 12544
rect 16252 12480 16258 12544
rect 15942 12479 16258 12480
rect 23716 12544 24032 12545
rect 23716 12480 23722 12544
rect 23786 12480 23802 12544
rect 23866 12480 23882 12544
rect 23946 12480 23962 12544
rect 24026 12480 24032 12544
rect 23716 12479 24032 12480
rect 31490 12544 31806 12545
rect 31490 12480 31496 12544
rect 31560 12480 31576 12544
rect 31640 12480 31656 12544
rect 31720 12480 31736 12544
rect 31800 12480 31806 12544
rect 31490 12479 31806 12480
rect 4281 12000 4597 12001
rect 4281 11936 4287 12000
rect 4351 11936 4367 12000
rect 4431 11936 4447 12000
rect 4511 11936 4527 12000
rect 4591 11936 4597 12000
rect 4281 11935 4597 11936
rect 12055 12000 12371 12001
rect 12055 11936 12061 12000
rect 12125 11936 12141 12000
rect 12205 11936 12221 12000
rect 12285 11936 12301 12000
rect 12365 11936 12371 12000
rect 12055 11935 12371 11936
rect 19829 12000 20145 12001
rect 19829 11936 19835 12000
rect 19899 11936 19915 12000
rect 19979 11936 19995 12000
rect 20059 11936 20075 12000
rect 20139 11936 20145 12000
rect 19829 11935 20145 11936
rect 27603 12000 27919 12001
rect 27603 11936 27609 12000
rect 27673 11936 27689 12000
rect 27753 11936 27769 12000
rect 27833 11936 27849 12000
rect 27913 11936 27919 12000
rect 27603 11935 27919 11936
rect 20989 11522 21055 11525
rect 21725 11522 21791 11525
rect 20989 11520 21791 11522
rect 20989 11464 20994 11520
rect 21050 11464 21730 11520
rect 21786 11464 21791 11520
rect 20989 11462 21791 11464
rect 20989 11459 21055 11462
rect 21725 11459 21791 11462
rect 8168 11456 8484 11457
rect 8168 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8484 11456
rect 8168 11391 8484 11392
rect 15942 11456 16258 11457
rect 15942 11392 15948 11456
rect 16012 11392 16028 11456
rect 16092 11392 16108 11456
rect 16172 11392 16188 11456
rect 16252 11392 16258 11456
rect 15942 11391 16258 11392
rect 23716 11456 24032 11457
rect 23716 11392 23722 11456
rect 23786 11392 23802 11456
rect 23866 11392 23882 11456
rect 23946 11392 23962 11456
rect 24026 11392 24032 11456
rect 23716 11391 24032 11392
rect 31490 11456 31806 11457
rect 31490 11392 31496 11456
rect 31560 11392 31576 11456
rect 31640 11392 31656 11456
rect 31720 11392 31736 11456
rect 31800 11392 31806 11456
rect 31490 11391 31806 11392
rect 4281 10912 4597 10913
rect 4281 10848 4287 10912
rect 4351 10848 4367 10912
rect 4431 10848 4447 10912
rect 4511 10848 4527 10912
rect 4591 10848 4597 10912
rect 4281 10847 4597 10848
rect 12055 10912 12371 10913
rect 12055 10848 12061 10912
rect 12125 10848 12141 10912
rect 12205 10848 12221 10912
rect 12285 10848 12301 10912
rect 12365 10848 12371 10912
rect 12055 10847 12371 10848
rect 19829 10912 20145 10913
rect 19829 10848 19835 10912
rect 19899 10848 19915 10912
rect 19979 10848 19995 10912
rect 20059 10848 20075 10912
rect 20139 10848 20145 10912
rect 19829 10847 20145 10848
rect 27603 10912 27919 10913
rect 27603 10848 27609 10912
rect 27673 10848 27689 10912
rect 27753 10848 27769 10912
rect 27833 10848 27849 10912
rect 27913 10848 27919 10912
rect 27603 10847 27919 10848
rect 8168 10368 8484 10369
rect 8168 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8484 10368
rect 8168 10303 8484 10304
rect 15942 10368 16258 10369
rect 15942 10304 15948 10368
rect 16012 10304 16028 10368
rect 16092 10304 16108 10368
rect 16172 10304 16188 10368
rect 16252 10304 16258 10368
rect 15942 10303 16258 10304
rect 23716 10368 24032 10369
rect 23716 10304 23722 10368
rect 23786 10304 23802 10368
rect 23866 10304 23882 10368
rect 23946 10304 23962 10368
rect 24026 10304 24032 10368
rect 23716 10303 24032 10304
rect 31490 10368 31806 10369
rect 31490 10304 31496 10368
rect 31560 10304 31576 10368
rect 31640 10304 31656 10368
rect 31720 10304 31736 10368
rect 31800 10304 31806 10368
rect 31490 10303 31806 10304
rect 4281 9824 4597 9825
rect 4281 9760 4287 9824
rect 4351 9760 4367 9824
rect 4431 9760 4447 9824
rect 4511 9760 4527 9824
rect 4591 9760 4597 9824
rect 4281 9759 4597 9760
rect 12055 9824 12371 9825
rect 12055 9760 12061 9824
rect 12125 9760 12141 9824
rect 12205 9760 12221 9824
rect 12285 9760 12301 9824
rect 12365 9760 12371 9824
rect 12055 9759 12371 9760
rect 19829 9824 20145 9825
rect 19829 9760 19835 9824
rect 19899 9760 19915 9824
rect 19979 9760 19995 9824
rect 20059 9760 20075 9824
rect 20139 9760 20145 9824
rect 19829 9759 20145 9760
rect 27603 9824 27919 9825
rect 27603 9760 27609 9824
rect 27673 9760 27689 9824
rect 27753 9760 27769 9824
rect 27833 9760 27849 9824
rect 27913 9760 27919 9824
rect 27603 9759 27919 9760
rect 8168 9280 8484 9281
rect 8168 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8484 9280
rect 8168 9215 8484 9216
rect 15942 9280 16258 9281
rect 15942 9216 15948 9280
rect 16012 9216 16028 9280
rect 16092 9216 16108 9280
rect 16172 9216 16188 9280
rect 16252 9216 16258 9280
rect 15942 9215 16258 9216
rect 23716 9280 24032 9281
rect 23716 9216 23722 9280
rect 23786 9216 23802 9280
rect 23866 9216 23882 9280
rect 23946 9216 23962 9280
rect 24026 9216 24032 9280
rect 23716 9215 24032 9216
rect 31490 9280 31806 9281
rect 31490 9216 31496 9280
rect 31560 9216 31576 9280
rect 31640 9216 31656 9280
rect 31720 9216 31736 9280
rect 31800 9216 31806 9280
rect 31490 9215 31806 9216
rect 4281 8736 4597 8737
rect 4281 8672 4287 8736
rect 4351 8672 4367 8736
rect 4431 8672 4447 8736
rect 4511 8672 4527 8736
rect 4591 8672 4597 8736
rect 4281 8671 4597 8672
rect 12055 8736 12371 8737
rect 12055 8672 12061 8736
rect 12125 8672 12141 8736
rect 12205 8672 12221 8736
rect 12285 8672 12301 8736
rect 12365 8672 12371 8736
rect 12055 8671 12371 8672
rect 19829 8736 20145 8737
rect 19829 8672 19835 8736
rect 19899 8672 19915 8736
rect 19979 8672 19995 8736
rect 20059 8672 20075 8736
rect 20139 8672 20145 8736
rect 19829 8671 20145 8672
rect 27603 8736 27919 8737
rect 27603 8672 27609 8736
rect 27673 8672 27689 8736
rect 27753 8672 27769 8736
rect 27833 8672 27849 8736
rect 27913 8672 27919 8736
rect 27603 8671 27919 8672
rect 8168 8192 8484 8193
rect 8168 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8484 8192
rect 8168 8127 8484 8128
rect 15942 8192 16258 8193
rect 15942 8128 15948 8192
rect 16012 8128 16028 8192
rect 16092 8128 16108 8192
rect 16172 8128 16188 8192
rect 16252 8128 16258 8192
rect 15942 8127 16258 8128
rect 23716 8192 24032 8193
rect 23716 8128 23722 8192
rect 23786 8128 23802 8192
rect 23866 8128 23882 8192
rect 23946 8128 23962 8192
rect 24026 8128 24032 8192
rect 23716 8127 24032 8128
rect 31490 8192 31806 8193
rect 31490 8128 31496 8192
rect 31560 8128 31576 8192
rect 31640 8128 31656 8192
rect 31720 8128 31736 8192
rect 31800 8128 31806 8192
rect 31490 8127 31806 8128
rect 4281 7648 4597 7649
rect 4281 7584 4287 7648
rect 4351 7584 4367 7648
rect 4431 7584 4447 7648
rect 4511 7584 4527 7648
rect 4591 7584 4597 7648
rect 4281 7583 4597 7584
rect 12055 7648 12371 7649
rect 12055 7584 12061 7648
rect 12125 7584 12141 7648
rect 12205 7584 12221 7648
rect 12285 7584 12301 7648
rect 12365 7584 12371 7648
rect 12055 7583 12371 7584
rect 19829 7648 20145 7649
rect 19829 7584 19835 7648
rect 19899 7584 19915 7648
rect 19979 7584 19995 7648
rect 20059 7584 20075 7648
rect 20139 7584 20145 7648
rect 19829 7583 20145 7584
rect 27603 7648 27919 7649
rect 27603 7584 27609 7648
rect 27673 7584 27689 7648
rect 27753 7584 27769 7648
rect 27833 7584 27849 7648
rect 27913 7584 27919 7648
rect 27603 7583 27919 7584
rect 8168 7104 8484 7105
rect 8168 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8484 7104
rect 8168 7039 8484 7040
rect 15942 7104 16258 7105
rect 15942 7040 15948 7104
rect 16012 7040 16028 7104
rect 16092 7040 16108 7104
rect 16172 7040 16188 7104
rect 16252 7040 16258 7104
rect 15942 7039 16258 7040
rect 23716 7104 24032 7105
rect 23716 7040 23722 7104
rect 23786 7040 23802 7104
rect 23866 7040 23882 7104
rect 23946 7040 23962 7104
rect 24026 7040 24032 7104
rect 23716 7039 24032 7040
rect 31490 7104 31806 7105
rect 31490 7040 31496 7104
rect 31560 7040 31576 7104
rect 31640 7040 31656 7104
rect 31720 7040 31736 7104
rect 31800 7040 31806 7104
rect 31490 7039 31806 7040
rect 4281 6560 4597 6561
rect 4281 6496 4287 6560
rect 4351 6496 4367 6560
rect 4431 6496 4447 6560
rect 4511 6496 4527 6560
rect 4591 6496 4597 6560
rect 4281 6495 4597 6496
rect 12055 6560 12371 6561
rect 12055 6496 12061 6560
rect 12125 6496 12141 6560
rect 12205 6496 12221 6560
rect 12285 6496 12301 6560
rect 12365 6496 12371 6560
rect 12055 6495 12371 6496
rect 19829 6560 20145 6561
rect 19829 6496 19835 6560
rect 19899 6496 19915 6560
rect 19979 6496 19995 6560
rect 20059 6496 20075 6560
rect 20139 6496 20145 6560
rect 19829 6495 20145 6496
rect 27603 6560 27919 6561
rect 27603 6496 27609 6560
rect 27673 6496 27689 6560
rect 27753 6496 27769 6560
rect 27833 6496 27849 6560
rect 27913 6496 27919 6560
rect 27603 6495 27919 6496
rect 8168 6016 8484 6017
rect 8168 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8484 6016
rect 8168 5951 8484 5952
rect 15942 6016 16258 6017
rect 15942 5952 15948 6016
rect 16012 5952 16028 6016
rect 16092 5952 16108 6016
rect 16172 5952 16188 6016
rect 16252 5952 16258 6016
rect 15942 5951 16258 5952
rect 23716 6016 24032 6017
rect 23716 5952 23722 6016
rect 23786 5952 23802 6016
rect 23866 5952 23882 6016
rect 23946 5952 23962 6016
rect 24026 5952 24032 6016
rect 23716 5951 24032 5952
rect 31490 6016 31806 6017
rect 31490 5952 31496 6016
rect 31560 5952 31576 6016
rect 31640 5952 31656 6016
rect 31720 5952 31736 6016
rect 31800 5952 31806 6016
rect 31490 5951 31806 5952
rect 4281 5472 4597 5473
rect 4281 5408 4287 5472
rect 4351 5408 4367 5472
rect 4431 5408 4447 5472
rect 4511 5408 4527 5472
rect 4591 5408 4597 5472
rect 4281 5407 4597 5408
rect 12055 5472 12371 5473
rect 12055 5408 12061 5472
rect 12125 5408 12141 5472
rect 12205 5408 12221 5472
rect 12285 5408 12301 5472
rect 12365 5408 12371 5472
rect 12055 5407 12371 5408
rect 19829 5472 20145 5473
rect 19829 5408 19835 5472
rect 19899 5408 19915 5472
rect 19979 5408 19995 5472
rect 20059 5408 20075 5472
rect 20139 5408 20145 5472
rect 19829 5407 20145 5408
rect 27603 5472 27919 5473
rect 27603 5408 27609 5472
rect 27673 5408 27689 5472
rect 27753 5408 27769 5472
rect 27833 5408 27849 5472
rect 27913 5408 27919 5472
rect 27603 5407 27919 5408
rect 8168 4928 8484 4929
rect 8168 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8484 4928
rect 8168 4863 8484 4864
rect 15942 4928 16258 4929
rect 15942 4864 15948 4928
rect 16012 4864 16028 4928
rect 16092 4864 16108 4928
rect 16172 4864 16188 4928
rect 16252 4864 16258 4928
rect 15942 4863 16258 4864
rect 23716 4928 24032 4929
rect 23716 4864 23722 4928
rect 23786 4864 23802 4928
rect 23866 4864 23882 4928
rect 23946 4864 23962 4928
rect 24026 4864 24032 4928
rect 23716 4863 24032 4864
rect 31490 4928 31806 4929
rect 31490 4864 31496 4928
rect 31560 4864 31576 4928
rect 31640 4864 31656 4928
rect 31720 4864 31736 4928
rect 31800 4864 31806 4928
rect 31490 4863 31806 4864
rect 4281 4384 4597 4385
rect 4281 4320 4287 4384
rect 4351 4320 4367 4384
rect 4431 4320 4447 4384
rect 4511 4320 4527 4384
rect 4591 4320 4597 4384
rect 4281 4319 4597 4320
rect 12055 4384 12371 4385
rect 12055 4320 12061 4384
rect 12125 4320 12141 4384
rect 12205 4320 12221 4384
rect 12285 4320 12301 4384
rect 12365 4320 12371 4384
rect 12055 4319 12371 4320
rect 19829 4384 20145 4385
rect 19829 4320 19835 4384
rect 19899 4320 19915 4384
rect 19979 4320 19995 4384
rect 20059 4320 20075 4384
rect 20139 4320 20145 4384
rect 19829 4319 20145 4320
rect 27603 4384 27919 4385
rect 27603 4320 27609 4384
rect 27673 4320 27689 4384
rect 27753 4320 27769 4384
rect 27833 4320 27849 4384
rect 27913 4320 27919 4384
rect 27603 4319 27919 4320
rect 8168 3840 8484 3841
rect 8168 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8484 3840
rect 8168 3775 8484 3776
rect 15942 3840 16258 3841
rect 15942 3776 15948 3840
rect 16012 3776 16028 3840
rect 16092 3776 16108 3840
rect 16172 3776 16188 3840
rect 16252 3776 16258 3840
rect 15942 3775 16258 3776
rect 23716 3840 24032 3841
rect 23716 3776 23722 3840
rect 23786 3776 23802 3840
rect 23866 3776 23882 3840
rect 23946 3776 23962 3840
rect 24026 3776 24032 3840
rect 23716 3775 24032 3776
rect 31490 3840 31806 3841
rect 31490 3776 31496 3840
rect 31560 3776 31576 3840
rect 31640 3776 31656 3840
rect 31720 3776 31736 3840
rect 31800 3776 31806 3840
rect 31490 3775 31806 3776
rect 4281 3296 4597 3297
rect 4281 3232 4287 3296
rect 4351 3232 4367 3296
rect 4431 3232 4447 3296
rect 4511 3232 4527 3296
rect 4591 3232 4597 3296
rect 4281 3231 4597 3232
rect 12055 3296 12371 3297
rect 12055 3232 12061 3296
rect 12125 3232 12141 3296
rect 12205 3232 12221 3296
rect 12285 3232 12301 3296
rect 12365 3232 12371 3296
rect 12055 3231 12371 3232
rect 19829 3296 20145 3297
rect 19829 3232 19835 3296
rect 19899 3232 19915 3296
rect 19979 3232 19995 3296
rect 20059 3232 20075 3296
rect 20139 3232 20145 3296
rect 19829 3231 20145 3232
rect 27603 3296 27919 3297
rect 27603 3232 27609 3296
rect 27673 3232 27689 3296
rect 27753 3232 27769 3296
rect 27833 3232 27849 3296
rect 27913 3232 27919 3296
rect 27603 3231 27919 3232
rect 8168 2752 8484 2753
rect 8168 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8484 2752
rect 8168 2687 8484 2688
rect 15942 2752 16258 2753
rect 15942 2688 15948 2752
rect 16012 2688 16028 2752
rect 16092 2688 16108 2752
rect 16172 2688 16188 2752
rect 16252 2688 16258 2752
rect 15942 2687 16258 2688
rect 23716 2752 24032 2753
rect 23716 2688 23722 2752
rect 23786 2688 23802 2752
rect 23866 2688 23882 2752
rect 23946 2688 23962 2752
rect 24026 2688 24032 2752
rect 23716 2687 24032 2688
rect 31490 2752 31806 2753
rect 31490 2688 31496 2752
rect 31560 2688 31576 2752
rect 31640 2688 31656 2752
rect 31720 2688 31736 2752
rect 31800 2688 31806 2752
rect 31490 2687 31806 2688
rect 4281 2208 4597 2209
rect 4281 2144 4287 2208
rect 4351 2144 4367 2208
rect 4431 2144 4447 2208
rect 4511 2144 4527 2208
rect 4591 2144 4597 2208
rect 4281 2143 4597 2144
rect 12055 2208 12371 2209
rect 12055 2144 12061 2208
rect 12125 2144 12141 2208
rect 12205 2144 12221 2208
rect 12285 2144 12301 2208
rect 12365 2144 12371 2208
rect 12055 2143 12371 2144
rect 19829 2208 20145 2209
rect 19829 2144 19835 2208
rect 19899 2144 19915 2208
rect 19979 2144 19995 2208
rect 20059 2144 20075 2208
rect 20139 2144 20145 2208
rect 19829 2143 20145 2144
rect 27603 2208 27919 2209
rect 27603 2144 27609 2208
rect 27673 2144 27689 2208
rect 27753 2144 27769 2208
rect 27833 2144 27849 2208
rect 27913 2144 27919 2208
rect 27603 2143 27919 2144
rect 8168 1664 8484 1665
rect 8168 1600 8174 1664
rect 8238 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8484 1664
rect 8168 1599 8484 1600
rect 15942 1664 16258 1665
rect 15942 1600 15948 1664
rect 16012 1600 16028 1664
rect 16092 1600 16108 1664
rect 16172 1600 16188 1664
rect 16252 1600 16258 1664
rect 15942 1599 16258 1600
rect 23716 1664 24032 1665
rect 23716 1600 23722 1664
rect 23786 1600 23802 1664
rect 23866 1600 23882 1664
rect 23946 1600 23962 1664
rect 24026 1600 24032 1664
rect 23716 1599 24032 1600
rect 31490 1664 31806 1665
rect 31490 1600 31496 1664
rect 31560 1600 31576 1664
rect 31640 1600 31656 1664
rect 31720 1600 31736 1664
rect 31800 1600 31806 1664
rect 31490 1599 31806 1600
rect 4281 1120 4597 1121
rect 4281 1056 4287 1120
rect 4351 1056 4367 1120
rect 4431 1056 4447 1120
rect 4511 1056 4527 1120
rect 4591 1056 4597 1120
rect 4281 1055 4597 1056
rect 12055 1120 12371 1121
rect 12055 1056 12061 1120
rect 12125 1056 12141 1120
rect 12205 1056 12221 1120
rect 12285 1056 12301 1120
rect 12365 1056 12371 1120
rect 12055 1055 12371 1056
rect 19829 1120 20145 1121
rect 19829 1056 19835 1120
rect 19899 1056 19915 1120
rect 19979 1056 19995 1120
rect 20059 1056 20075 1120
rect 20139 1056 20145 1120
rect 19829 1055 20145 1056
rect 27603 1120 27919 1121
rect 27603 1056 27609 1120
rect 27673 1056 27689 1120
rect 27753 1056 27769 1120
rect 27833 1056 27849 1120
rect 27913 1056 27919 1120
rect 27603 1055 27919 1056
rect 8168 576 8484 577
rect 8168 512 8174 576
rect 8238 512 8254 576
rect 8318 512 8334 576
rect 8398 512 8414 576
rect 8478 512 8484 576
rect 8168 511 8484 512
rect 15942 576 16258 577
rect 15942 512 15948 576
rect 16012 512 16028 576
rect 16092 512 16108 576
rect 16172 512 16188 576
rect 16252 512 16258 576
rect 15942 511 16258 512
rect 23716 576 24032 577
rect 23716 512 23722 576
rect 23786 512 23802 576
rect 23866 512 23882 576
rect 23946 512 23962 576
rect 24026 512 24032 576
rect 23716 511 24032 512
rect 31490 576 31806 577
rect 31490 512 31496 576
rect 31560 512 31576 576
rect 31640 512 31656 576
rect 31720 512 31736 576
rect 31800 512 31806 576
rect 31490 511 31806 512
<< via3 >>
rect 4476 21992 4540 21996
rect 4476 21936 4526 21992
rect 4526 21936 4540 21992
rect 4476 21932 4540 21936
rect 8156 21992 8220 21996
rect 8156 21936 8206 21992
rect 8206 21936 8220 21992
rect 8156 21932 8220 21936
rect 27476 21932 27540 21996
rect 796 21856 860 21860
rect 796 21800 846 21856
rect 846 21800 860 21856
rect 796 21796 860 21800
rect 1532 21856 1596 21860
rect 1532 21800 1582 21856
rect 1582 21800 1596 21856
rect 1532 21796 1596 21800
rect 2268 21856 2332 21860
rect 2268 21800 2318 21856
rect 2318 21800 2332 21856
rect 2268 21796 2332 21800
rect 3004 21796 3068 21860
rect 3740 21856 3804 21860
rect 3740 21800 3790 21856
rect 3790 21800 3804 21856
rect 3740 21796 3804 21800
rect 5212 21856 5276 21860
rect 5212 21800 5262 21856
rect 5262 21800 5276 21856
rect 5212 21796 5276 21800
rect 5948 21856 6012 21860
rect 5948 21800 5998 21856
rect 5998 21800 6012 21856
rect 5948 21796 6012 21800
rect 6684 21856 6748 21860
rect 6684 21800 6734 21856
rect 6734 21800 6748 21856
rect 6684 21796 6748 21800
rect 7420 21856 7484 21860
rect 7420 21800 7470 21856
rect 7470 21800 7484 21856
rect 7420 21796 7484 21800
rect 8892 21796 8956 21860
rect 9628 21856 9692 21860
rect 9628 21800 9678 21856
rect 9678 21800 9692 21856
rect 9628 21796 9692 21800
rect 10364 21856 10428 21860
rect 10364 21800 10414 21856
rect 10414 21800 10428 21856
rect 10364 21796 10428 21800
rect 11100 21856 11164 21860
rect 11100 21800 11150 21856
rect 11150 21800 11164 21856
rect 11100 21796 11164 21800
rect 25820 21856 25884 21860
rect 25820 21800 25870 21856
rect 25870 21800 25884 21856
rect 25820 21796 25884 21800
rect 26556 21796 26620 21860
rect 28028 21796 28092 21860
rect 29500 21796 29564 21860
rect 4287 21788 4351 21792
rect 4287 21732 4291 21788
rect 4291 21732 4347 21788
rect 4347 21732 4351 21788
rect 4287 21728 4351 21732
rect 4367 21788 4431 21792
rect 4367 21732 4371 21788
rect 4371 21732 4427 21788
rect 4427 21732 4431 21788
rect 4367 21728 4431 21732
rect 4447 21788 4511 21792
rect 4447 21732 4451 21788
rect 4451 21732 4507 21788
rect 4507 21732 4511 21788
rect 4447 21728 4511 21732
rect 4527 21788 4591 21792
rect 4527 21732 4531 21788
rect 4531 21732 4587 21788
rect 4587 21732 4591 21788
rect 4527 21728 4591 21732
rect 12061 21788 12125 21792
rect 12061 21732 12065 21788
rect 12065 21732 12121 21788
rect 12121 21732 12125 21788
rect 12061 21728 12125 21732
rect 12141 21788 12205 21792
rect 12141 21732 12145 21788
rect 12145 21732 12201 21788
rect 12201 21732 12205 21788
rect 12141 21728 12205 21732
rect 12221 21788 12285 21792
rect 12221 21732 12225 21788
rect 12225 21732 12281 21788
rect 12281 21732 12285 21788
rect 12221 21728 12285 21732
rect 12301 21788 12365 21792
rect 12301 21732 12305 21788
rect 12305 21732 12361 21788
rect 12361 21732 12365 21788
rect 12301 21728 12365 21732
rect 19835 21788 19899 21792
rect 19835 21732 19839 21788
rect 19839 21732 19895 21788
rect 19895 21732 19899 21788
rect 19835 21728 19899 21732
rect 19915 21788 19979 21792
rect 19915 21732 19919 21788
rect 19919 21732 19975 21788
rect 19975 21732 19979 21788
rect 19915 21728 19979 21732
rect 19995 21788 20059 21792
rect 19995 21732 19999 21788
rect 19999 21732 20055 21788
rect 20055 21732 20059 21788
rect 19995 21728 20059 21732
rect 20075 21788 20139 21792
rect 20075 21732 20079 21788
rect 20079 21732 20135 21788
rect 20135 21732 20139 21788
rect 20075 21728 20139 21732
rect 27609 21788 27673 21792
rect 27609 21732 27613 21788
rect 27613 21732 27669 21788
rect 27669 21732 27673 21788
rect 27609 21728 27673 21732
rect 27689 21788 27753 21792
rect 27689 21732 27693 21788
rect 27693 21732 27749 21788
rect 27749 21732 27753 21788
rect 27689 21728 27753 21732
rect 27769 21788 27833 21792
rect 27769 21732 27773 21788
rect 27773 21732 27829 21788
rect 27829 21732 27833 21788
rect 27769 21728 27833 21732
rect 27849 21788 27913 21792
rect 27849 21732 27853 21788
rect 27853 21732 27909 21788
rect 27909 21732 27913 21788
rect 27849 21728 27913 21732
rect 28764 21660 28828 21724
rect 11836 21584 11900 21588
rect 11836 21528 11886 21584
rect 11886 21528 11900 21584
rect 11836 21524 11900 21528
rect 13308 21584 13372 21588
rect 13308 21528 13358 21584
rect 13358 21528 13372 21584
rect 13308 21524 13372 21528
rect 16988 21252 17052 21316
rect 8174 21244 8238 21248
rect 8174 21188 8178 21244
rect 8178 21188 8234 21244
rect 8234 21188 8238 21244
rect 8174 21184 8238 21188
rect 8254 21244 8318 21248
rect 8254 21188 8258 21244
rect 8258 21188 8314 21244
rect 8314 21188 8318 21244
rect 8254 21184 8318 21188
rect 8334 21244 8398 21248
rect 8334 21188 8338 21244
rect 8338 21188 8394 21244
rect 8394 21188 8398 21244
rect 8334 21184 8398 21188
rect 8414 21244 8478 21248
rect 8414 21188 8418 21244
rect 8418 21188 8474 21244
rect 8474 21188 8478 21244
rect 8414 21184 8478 21188
rect 15948 21244 16012 21248
rect 15948 21188 15952 21244
rect 15952 21188 16008 21244
rect 16008 21188 16012 21244
rect 15948 21184 16012 21188
rect 16028 21244 16092 21248
rect 16028 21188 16032 21244
rect 16032 21188 16088 21244
rect 16088 21188 16092 21244
rect 16028 21184 16092 21188
rect 16108 21244 16172 21248
rect 16108 21188 16112 21244
rect 16112 21188 16168 21244
rect 16168 21188 16172 21244
rect 16108 21184 16172 21188
rect 16188 21244 16252 21248
rect 16188 21188 16192 21244
rect 16192 21188 16248 21244
rect 16248 21188 16252 21244
rect 16188 21184 16252 21188
rect 23722 21244 23786 21248
rect 23722 21188 23726 21244
rect 23726 21188 23782 21244
rect 23782 21188 23786 21244
rect 23722 21184 23786 21188
rect 23802 21244 23866 21248
rect 23802 21188 23806 21244
rect 23806 21188 23862 21244
rect 23862 21188 23866 21244
rect 23802 21184 23866 21188
rect 23882 21244 23946 21248
rect 23882 21188 23886 21244
rect 23886 21188 23942 21244
rect 23942 21188 23946 21244
rect 23882 21184 23946 21188
rect 23962 21244 24026 21248
rect 23962 21188 23966 21244
rect 23966 21188 24022 21244
rect 24022 21188 24026 21244
rect 23962 21184 24026 21188
rect 31496 21244 31560 21248
rect 31496 21188 31500 21244
rect 31500 21188 31556 21244
rect 31556 21188 31560 21244
rect 31496 21184 31560 21188
rect 31576 21244 31640 21248
rect 31576 21188 31580 21244
rect 31580 21188 31636 21244
rect 31636 21188 31640 21244
rect 31576 21184 31640 21188
rect 31656 21244 31720 21248
rect 31656 21188 31660 21244
rect 31660 21188 31716 21244
rect 31716 21188 31720 21244
rect 31656 21184 31720 21188
rect 31736 21244 31800 21248
rect 31736 21188 31740 21244
rect 31740 21188 31796 21244
rect 31796 21188 31800 21244
rect 31736 21184 31800 21188
rect 14044 20708 14108 20772
rect 4287 20700 4351 20704
rect 4287 20644 4291 20700
rect 4291 20644 4347 20700
rect 4347 20644 4351 20700
rect 4287 20640 4351 20644
rect 4367 20700 4431 20704
rect 4367 20644 4371 20700
rect 4371 20644 4427 20700
rect 4427 20644 4431 20700
rect 4367 20640 4431 20644
rect 4447 20700 4511 20704
rect 4447 20644 4451 20700
rect 4451 20644 4507 20700
rect 4507 20644 4511 20700
rect 4447 20640 4511 20644
rect 4527 20700 4591 20704
rect 4527 20644 4531 20700
rect 4531 20644 4587 20700
rect 4587 20644 4591 20700
rect 4527 20640 4591 20644
rect 12061 20700 12125 20704
rect 12061 20644 12065 20700
rect 12065 20644 12121 20700
rect 12121 20644 12125 20700
rect 12061 20640 12125 20644
rect 12141 20700 12205 20704
rect 12141 20644 12145 20700
rect 12145 20644 12201 20700
rect 12201 20644 12205 20700
rect 12141 20640 12205 20644
rect 12221 20700 12285 20704
rect 12221 20644 12225 20700
rect 12225 20644 12281 20700
rect 12281 20644 12285 20700
rect 12221 20640 12285 20644
rect 12301 20700 12365 20704
rect 12301 20644 12305 20700
rect 12305 20644 12361 20700
rect 12361 20644 12365 20700
rect 12301 20640 12365 20644
rect 19835 20700 19899 20704
rect 19835 20644 19839 20700
rect 19839 20644 19895 20700
rect 19895 20644 19899 20700
rect 19835 20640 19899 20644
rect 19915 20700 19979 20704
rect 19915 20644 19919 20700
rect 19919 20644 19975 20700
rect 19975 20644 19979 20700
rect 19915 20640 19979 20644
rect 19995 20700 20059 20704
rect 19995 20644 19999 20700
rect 19999 20644 20055 20700
rect 20055 20644 20059 20700
rect 19995 20640 20059 20644
rect 20075 20700 20139 20704
rect 20075 20644 20079 20700
rect 20079 20644 20135 20700
rect 20135 20644 20139 20700
rect 20075 20640 20139 20644
rect 27609 20700 27673 20704
rect 27609 20644 27613 20700
rect 27613 20644 27669 20700
rect 27669 20644 27673 20700
rect 27609 20640 27673 20644
rect 27689 20700 27753 20704
rect 27689 20644 27693 20700
rect 27693 20644 27749 20700
rect 27749 20644 27753 20700
rect 27689 20640 27753 20644
rect 27769 20700 27833 20704
rect 27769 20644 27773 20700
rect 27773 20644 27829 20700
rect 27829 20644 27833 20700
rect 27769 20640 27833 20644
rect 27849 20700 27913 20704
rect 27849 20644 27853 20700
rect 27853 20644 27909 20700
rect 27909 20644 27913 20700
rect 27849 20640 27913 20644
rect 12940 20436 13004 20500
rect 8174 20156 8238 20160
rect 8174 20100 8178 20156
rect 8178 20100 8234 20156
rect 8234 20100 8238 20156
rect 8174 20096 8238 20100
rect 8254 20156 8318 20160
rect 8254 20100 8258 20156
rect 8258 20100 8314 20156
rect 8314 20100 8318 20156
rect 8254 20096 8318 20100
rect 8334 20156 8398 20160
rect 8334 20100 8338 20156
rect 8338 20100 8394 20156
rect 8394 20100 8398 20156
rect 8334 20096 8398 20100
rect 8414 20156 8478 20160
rect 8414 20100 8418 20156
rect 8418 20100 8474 20156
rect 8474 20100 8478 20156
rect 8414 20096 8478 20100
rect 15948 20156 16012 20160
rect 15948 20100 15952 20156
rect 15952 20100 16008 20156
rect 16008 20100 16012 20156
rect 15948 20096 16012 20100
rect 16028 20156 16092 20160
rect 16028 20100 16032 20156
rect 16032 20100 16088 20156
rect 16088 20100 16092 20156
rect 16028 20096 16092 20100
rect 16108 20156 16172 20160
rect 16108 20100 16112 20156
rect 16112 20100 16168 20156
rect 16168 20100 16172 20156
rect 16108 20096 16172 20100
rect 16188 20156 16252 20160
rect 16188 20100 16192 20156
rect 16192 20100 16248 20156
rect 16248 20100 16252 20156
rect 16188 20096 16252 20100
rect 23722 20156 23786 20160
rect 23722 20100 23726 20156
rect 23726 20100 23782 20156
rect 23782 20100 23786 20156
rect 23722 20096 23786 20100
rect 23802 20156 23866 20160
rect 23802 20100 23806 20156
rect 23806 20100 23862 20156
rect 23862 20100 23866 20156
rect 23802 20096 23866 20100
rect 23882 20156 23946 20160
rect 23882 20100 23886 20156
rect 23886 20100 23942 20156
rect 23942 20100 23946 20156
rect 23882 20096 23946 20100
rect 23962 20156 24026 20160
rect 23962 20100 23966 20156
rect 23966 20100 24022 20156
rect 24022 20100 24026 20156
rect 23962 20096 24026 20100
rect 31496 20156 31560 20160
rect 31496 20100 31500 20156
rect 31500 20100 31556 20156
rect 31556 20100 31560 20156
rect 31496 20096 31560 20100
rect 31576 20156 31640 20160
rect 31576 20100 31580 20156
rect 31580 20100 31636 20156
rect 31636 20100 31640 20156
rect 31576 20096 31640 20100
rect 31656 20156 31720 20160
rect 31656 20100 31660 20156
rect 31660 20100 31716 20156
rect 31716 20100 31720 20156
rect 31656 20096 31720 20100
rect 31736 20156 31800 20160
rect 31736 20100 31740 20156
rect 31740 20100 31796 20156
rect 31796 20100 31800 20156
rect 31736 20096 31800 20100
rect 4287 19612 4351 19616
rect 4287 19556 4291 19612
rect 4291 19556 4347 19612
rect 4347 19556 4351 19612
rect 4287 19552 4351 19556
rect 4367 19612 4431 19616
rect 4367 19556 4371 19612
rect 4371 19556 4427 19612
rect 4427 19556 4431 19612
rect 4367 19552 4431 19556
rect 4447 19612 4511 19616
rect 4447 19556 4451 19612
rect 4451 19556 4507 19612
rect 4507 19556 4511 19612
rect 4447 19552 4511 19556
rect 4527 19612 4591 19616
rect 4527 19556 4531 19612
rect 4531 19556 4587 19612
rect 4587 19556 4591 19612
rect 4527 19552 4591 19556
rect 12061 19612 12125 19616
rect 12061 19556 12065 19612
rect 12065 19556 12121 19612
rect 12121 19556 12125 19612
rect 12061 19552 12125 19556
rect 12141 19612 12205 19616
rect 12141 19556 12145 19612
rect 12145 19556 12201 19612
rect 12201 19556 12205 19612
rect 12141 19552 12205 19556
rect 12221 19612 12285 19616
rect 12221 19556 12225 19612
rect 12225 19556 12281 19612
rect 12281 19556 12285 19612
rect 12221 19552 12285 19556
rect 12301 19612 12365 19616
rect 12301 19556 12305 19612
rect 12305 19556 12361 19612
rect 12361 19556 12365 19612
rect 12301 19552 12365 19556
rect 19835 19612 19899 19616
rect 19835 19556 19839 19612
rect 19839 19556 19895 19612
rect 19895 19556 19899 19612
rect 19835 19552 19899 19556
rect 19915 19612 19979 19616
rect 19915 19556 19919 19612
rect 19919 19556 19975 19612
rect 19975 19556 19979 19612
rect 19915 19552 19979 19556
rect 19995 19612 20059 19616
rect 19995 19556 19999 19612
rect 19999 19556 20055 19612
rect 20055 19556 20059 19612
rect 19995 19552 20059 19556
rect 20075 19612 20139 19616
rect 20075 19556 20079 19612
rect 20079 19556 20135 19612
rect 20135 19556 20139 19612
rect 20075 19552 20139 19556
rect 27609 19612 27673 19616
rect 27609 19556 27613 19612
rect 27613 19556 27669 19612
rect 27669 19556 27673 19612
rect 27609 19552 27673 19556
rect 27689 19612 27753 19616
rect 27689 19556 27693 19612
rect 27693 19556 27749 19612
rect 27749 19556 27753 19612
rect 27689 19552 27753 19556
rect 27769 19612 27833 19616
rect 27769 19556 27773 19612
rect 27773 19556 27829 19612
rect 27829 19556 27833 19612
rect 27769 19552 27833 19556
rect 27849 19612 27913 19616
rect 27849 19556 27853 19612
rect 27853 19556 27909 19612
rect 27909 19556 27913 19612
rect 27849 19552 27913 19556
rect 15516 19136 15580 19140
rect 15516 19080 15566 19136
rect 15566 19080 15580 19136
rect 15516 19076 15580 19080
rect 8174 19068 8238 19072
rect 8174 19012 8178 19068
rect 8178 19012 8234 19068
rect 8234 19012 8238 19068
rect 8174 19008 8238 19012
rect 8254 19068 8318 19072
rect 8254 19012 8258 19068
rect 8258 19012 8314 19068
rect 8314 19012 8318 19068
rect 8254 19008 8318 19012
rect 8334 19068 8398 19072
rect 8334 19012 8338 19068
rect 8338 19012 8394 19068
rect 8394 19012 8398 19068
rect 8334 19008 8398 19012
rect 8414 19068 8478 19072
rect 8414 19012 8418 19068
rect 8418 19012 8474 19068
rect 8474 19012 8478 19068
rect 8414 19008 8478 19012
rect 15948 19068 16012 19072
rect 15948 19012 15952 19068
rect 15952 19012 16008 19068
rect 16008 19012 16012 19068
rect 15948 19008 16012 19012
rect 16028 19068 16092 19072
rect 16028 19012 16032 19068
rect 16032 19012 16088 19068
rect 16088 19012 16092 19068
rect 16028 19008 16092 19012
rect 16108 19068 16172 19072
rect 16108 19012 16112 19068
rect 16112 19012 16168 19068
rect 16168 19012 16172 19068
rect 16108 19008 16172 19012
rect 16188 19068 16252 19072
rect 16188 19012 16192 19068
rect 16192 19012 16248 19068
rect 16248 19012 16252 19068
rect 16188 19008 16252 19012
rect 23722 19068 23786 19072
rect 23722 19012 23726 19068
rect 23726 19012 23782 19068
rect 23782 19012 23786 19068
rect 23722 19008 23786 19012
rect 23802 19068 23866 19072
rect 23802 19012 23806 19068
rect 23806 19012 23862 19068
rect 23862 19012 23866 19068
rect 23802 19008 23866 19012
rect 23882 19068 23946 19072
rect 23882 19012 23886 19068
rect 23886 19012 23942 19068
rect 23942 19012 23946 19068
rect 23882 19008 23946 19012
rect 23962 19068 24026 19072
rect 23962 19012 23966 19068
rect 23966 19012 24022 19068
rect 24022 19012 24026 19068
rect 23962 19008 24026 19012
rect 31496 19068 31560 19072
rect 31496 19012 31500 19068
rect 31500 19012 31556 19068
rect 31556 19012 31560 19068
rect 31496 19008 31560 19012
rect 31576 19068 31640 19072
rect 31576 19012 31580 19068
rect 31580 19012 31636 19068
rect 31636 19012 31640 19068
rect 31576 19008 31640 19012
rect 31656 19068 31720 19072
rect 31656 19012 31660 19068
rect 31660 19012 31716 19068
rect 31716 19012 31720 19068
rect 31656 19008 31720 19012
rect 31736 19068 31800 19072
rect 31736 19012 31740 19068
rect 31740 19012 31796 19068
rect 31796 19012 31800 19068
rect 31736 19008 31800 19012
rect 4287 18524 4351 18528
rect 4287 18468 4291 18524
rect 4291 18468 4347 18524
rect 4347 18468 4351 18524
rect 4287 18464 4351 18468
rect 4367 18524 4431 18528
rect 4367 18468 4371 18524
rect 4371 18468 4427 18524
rect 4427 18468 4431 18524
rect 4367 18464 4431 18468
rect 4447 18524 4511 18528
rect 4447 18468 4451 18524
rect 4451 18468 4507 18524
rect 4507 18468 4511 18524
rect 4447 18464 4511 18468
rect 4527 18524 4591 18528
rect 4527 18468 4531 18524
rect 4531 18468 4587 18524
rect 4587 18468 4591 18524
rect 4527 18464 4591 18468
rect 12061 18524 12125 18528
rect 12061 18468 12065 18524
rect 12065 18468 12121 18524
rect 12121 18468 12125 18524
rect 12061 18464 12125 18468
rect 12141 18524 12205 18528
rect 12141 18468 12145 18524
rect 12145 18468 12201 18524
rect 12201 18468 12205 18524
rect 12141 18464 12205 18468
rect 12221 18524 12285 18528
rect 12221 18468 12225 18524
rect 12225 18468 12281 18524
rect 12281 18468 12285 18524
rect 12221 18464 12285 18468
rect 12301 18524 12365 18528
rect 12301 18468 12305 18524
rect 12305 18468 12361 18524
rect 12361 18468 12365 18524
rect 12301 18464 12365 18468
rect 19835 18524 19899 18528
rect 19835 18468 19839 18524
rect 19839 18468 19895 18524
rect 19895 18468 19899 18524
rect 19835 18464 19899 18468
rect 19915 18524 19979 18528
rect 19915 18468 19919 18524
rect 19919 18468 19975 18524
rect 19975 18468 19979 18524
rect 19915 18464 19979 18468
rect 19995 18524 20059 18528
rect 19995 18468 19999 18524
rect 19999 18468 20055 18524
rect 20055 18468 20059 18524
rect 19995 18464 20059 18468
rect 20075 18524 20139 18528
rect 20075 18468 20079 18524
rect 20079 18468 20135 18524
rect 20135 18468 20139 18524
rect 20075 18464 20139 18468
rect 27609 18524 27673 18528
rect 27609 18468 27613 18524
rect 27613 18468 27669 18524
rect 27669 18468 27673 18524
rect 27609 18464 27673 18468
rect 27689 18524 27753 18528
rect 27689 18468 27693 18524
rect 27693 18468 27749 18524
rect 27749 18468 27753 18524
rect 27689 18464 27753 18468
rect 27769 18524 27833 18528
rect 27769 18468 27773 18524
rect 27773 18468 27829 18524
rect 27829 18468 27833 18524
rect 27769 18464 27833 18468
rect 27849 18524 27913 18528
rect 27849 18468 27853 18524
rect 27853 18468 27909 18524
rect 27909 18468 27913 18524
rect 27849 18464 27913 18468
rect 8174 17980 8238 17984
rect 8174 17924 8178 17980
rect 8178 17924 8234 17980
rect 8234 17924 8238 17980
rect 8174 17920 8238 17924
rect 8254 17980 8318 17984
rect 8254 17924 8258 17980
rect 8258 17924 8314 17980
rect 8314 17924 8318 17980
rect 8254 17920 8318 17924
rect 8334 17980 8398 17984
rect 8334 17924 8338 17980
rect 8338 17924 8394 17980
rect 8394 17924 8398 17980
rect 8334 17920 8398 17924
rect 8414 17980 8478 17984
rect 8414 17924 8418 17980
rect 8418 17924 8474 17980
rect 8474 17924 8478 17980
rect 8414 17920 8478 17924
rect 15948 17980 16012 17984
rect 15948 17924 15952 17980
rect 15952 17924 16008 17980
rect 16008 17924 16012 17980
rect 15948 17920 16012 17924
rect 16028 17980 16092 17984
rect 16028 17924 16032 17980
rect 16032 17924 16088 17980
rect 16088 17924 16092 17980
rect 16028 17920 16092 17924
rect 16108 17980 16172 17984
rect 16108 17924 16112 17980
rect 16112 17924 16168 17980
rect 16168 17924 16172 17980
rect 16108 17920 16172 17924
rect 16188 17980 16252 17984
rect 16188 17924 16192 17980
rect 16192 17924 16248 17980
rect 16248 17924 16252 17980
rect 16188 17920 16252 17924
rect 23722 17980 23786 17984
rect 23722 17924 23726 17980
rect 23726 17924 23782 17980
rect 23782 17924 23786 17980
rect 23722 17920 23786 17924
rect 23802 17980 23866 17984
rect 23802 17924 23806 17980
rect 23806 17924 23862 17980
rect 23862 17924 23866 17980
rect 23802 17920 23866 17924
rect 23882 17980 23946 17984
rect 23882 17924 23886 17980
rect 23886 17924 23942 17980
rect 23942 17924 23946 17980
rect 23882 17920 23946 17924
rect 23962 17980 24026 17984
rect 23962 17924 23966 17980
rect 23966 17924 24022 17980
rect 24022 17924 24026 17980
rect 23962 17920 24026 17924
rect 31496 17980 31560 17984
rect 31496 17924 31500 17980
rect 31500 17924 31556 17980
rect 31556 17924 31560 17980
rect 31496 17920 31560 17924
rect 31576 17980 31640 17984
rect 31576 17924 31580 17980
rect 31580 17924 31636 17980
rect 31636 17924 31640 17980
rect 31576 17920 31640 17924
rect 31656 17980 31720 17984
rect 31656 17924 31660 17980
rect 31660 17924 31716 17980
rect 31716 17924 31720 17980
rect 31656 17920 31720 17924
rect 31736 17980 31800 17984
rect 31736 17924 31740 17980
rect 31740 17924 31796 17980
rect 31796 17924 31800 17980
rect 31736 17920 31800 17924
rect 14780 17912 14844 17916
rect 14780 17856 14794 17912
rect 14794 17856 14844 17912
rect 14780 17852 14844 17856
rect 16436 17852 16500 17916
rect 4287 17436 4351 17440
rect 4287 17380 4291 17436
rect 4291 17380 4347 17436
rect 4347 17380 4351 17436
rect 4287 17376 4351 17380
rect 4367 17436 4431 17440
rect 4367 17380 4371 17436
rect 4371 17380 4427 17436
rect 4427 17380 4431 17436
rect 4367 17376 4431 17380
rect 4447 17436 4511 17440
rect 4447 17380 4451 17436
rect 4451 17380 4507 17436
rect 4507 17380 4511 17436
rect 4447 17376 4511 17380
rect 4527 17436 4591 17440
rect 4527 17380 4531 17436
rect 4531 17380 4587 17436
rect 4587 17380 4591 17436
rect 4527 17376 4591 17380
rect 12061 17436 12125 17440
rect 12061 17380 12065 17436
rect 12065 17380 12121 17436
rect 12121 17380 12125 17436
rect 12061 17376 12125 17380
rect 12141 17436 12205 17440
rect 12141 17380 12145 17436
rect 12145 17380 12201 17436
rect 12201 17380 12205 17436
rect 12141 17376 12205 17380
rect 12221 17436 12285 17440
rect 12221 17380 12225 17436
rect 12225 17380 12281 17436
rect 12281 17380 12285 17436
rect 12221 17376 12285 17380
rect 12301 17436 12365 17440
rect 12301 17380 12305 17436
rect 12305 17380 12361 17436
rect 12361 17380 12365 17436
rect 12301 17376 12365 17380
rect 19835 17436 19899 17440
rect 19835 17380 19839 17436
rect 19839 17380 19895 17436
rect 19895 17380 19899 17436
rect 19835 17376 19899 17380
rect 19915 17436 19979 17440
rect 19915 17380 19919 17436
rect 19919 17380 19975 17436
rect 19975 17380 19979 17436
rect 19915 17376 19979 17380
rect 19995 17436 20059 17440
rect 19995 17380 19999 17436
rect 19999 17380 20055 17436
rect 20055 17380 20059 17436
rect 19995 17376 20059 17380
rect 20075 17436 20139 17440
rect 20075 17380 20079 17436
rect 20079 17380 20135 17436
rect 20135 17380 20139 17436
rect 20075 17376 20139 17380
rect 27609 17436 27673 17440
rect 27609 17380 27613 17436
rect 27613 17380 27669 17436
rect 27669 17380 27673 17436
rect 27609 17376 27673 17380
rect 27689 17436 27753 17440
rect 27689 17380 27693 17436
rect 27693 17380 27749 17436
rect 27749 17380 27753 17436
rect 27689 17376 27753 17380
rect 27769 17436 27833 17440
rect 27769 17380 27773 17436
rect 27773 17380 27829 17436
rect 27829 17380 27833 17436
rect 27769 17376 27833 17380
rect 27849 17436 27913 17440
rect 27849 17380 27853 17436
rect 27853 17380 27909 17436
rect 27909 17380 27913 17436
rect 27849 17376 27913 17380
rect 8174 16892 8238 16896
rect 8174 16836 8178 16892
rect 8178 16836 8234 16892
rect 8234 16836 8238 16892
rect 8174 16832 8238 16836
rect 8254 16892 8318 16896
rect 8254 16836 8258 16892
rect 8258 16836 8314 16892
rect 8314 16836 8318 16892
rect 8254 16832 8318 16836
rect 8334 16892 8398 16896
rect 8334 16836 8338 16892
rect 8338 16836 8394 16892
rect 8394 16836 8398 16892
rect 8334 16832 8398 16836
rect 8414 16892 8478 16896
rect 8414 16836 8418 16892
rect 8418 16836 8474 16892
rect 8474 16836 8478 16892
rect 8414 16832 8478 16836
rect 15948 16892 16012 16896
rect 15948 16836 15952 16892
rect 15952 16836 16008 16892
rect 16008 16836 16012 16892
rect 15948 16832 16012 16836
rect 16028 16892 16092 16896
rect 16028 16836 16032 16892
rect 16032 16836 16088 16892
rect 16088 16836 16092 16892
rect 16028 16832 16092 16836
rect 16108 16892 16172 16896
rect 16108 16836 16112 16892
rect 16112 16836 16168 16892
rect 16168 16836 16172 16892
rect 16108 16832 16172 16836
rect 16188 16892 16252 16896
rect 16188 16836 16192 16892
rect 16192 16836 16248 16892
rect 16248 16836 16252 16892
rect 16188 16832 16252 16836
rect 23722 16892 23786 16896
rect 23722 16836 23726 16892
rect 23726 16836 23782 16892
rect 23782 16836 23786 16892
rect 23722 16832 23786 16836
rect 23802 16892 23866 16896
rect 23802 16836 23806 16892
rect 23806 16836 23862 16892
rect 23862 16836 23866 16892
rect 23802 16832 23866 16836
rect 23882 16892 23946 16896
rect 23882 16836 23886 16892
rect 23886 16836 23942 16892
rect 23942 16836 23946 16892
rect 23882 16832 23946 16836
rect 23962 16892 24026 16896
rect 23962 16836 23966 16892
rect 23966 16836 24022 16892
rect 24022 16836 24026 16892
rect 23962 16832 24026 16836
rect 31496 16892 31560 16896
rect 31496 16836 31500 16892
rect 31500 16836 31556 16892
rect 31556 16836 31560 16892
rect 31496 16832 31560 16836
rect 31576 16892 31640 16896
rect 31576 16836 31580 16892
rect 31580 16836 31636 16892
rect 31636 16836 31640 16892
rect 31576 16832 31640 16836
rect 31656 16892 31720 16896
rect 31656 16836 31660 16892
rect 31660 16836 31716 16892
rect 31716 16836 31720 16892
rect 31656 16832 31720 16836
rect 31736 16892 31800 16896
rect 31736 16836 31740 16892
rect 31740 16836 31796 16892
rect 31796 16836 31800 16892
rect 31736 16832 31800 16836
rect 17724 16492 17788 16556
rect 4287 16348 4351 16352
rect 4287 16292 4291 16348
rect 4291 16292 4347 16348
rect 4347 16292 4351 16348
rect 4287 16288 4351 16292
rect 4367 16348 4431 16352
rect 4367 16292 4371 16348
rect 4371 16292 4427 16348
rect 4427 16292 4431 16348
rect 4367 16288 4431 16292
rect 4447 16348 4511 16352
rect 4447 16292 4451 16348
rect 4451 16292 4507 16348
rect 4507 16292 4511 16348
rect 4447 16288 4511 16292
rect 4527 16348 4591 16352
rect 4527 16292 4531 16348
rect 4531 16292 4587 16348
rect 4587 16292 4591 16348
rect 4527 16288 4591 16292
rect 12061 16348 12125 16352
rect 12061 16292 12065 16348
rect 12065 16292 12121 16348
rect 12121 16292 12125 16348
rect 12061 16288 12125 16292
rect 12141 16348 12205 16352
rect 12141 16292 12145 16348
rect 12145 16292 12201 16348
rect 12201 16292 12205 16348
rect 12141 16288 12205 16292
rect 12221 16348 12285 16352
rect 12221 16292 12225 16348
rect 12225 16292 12281 16348
rect 12281 16292 12285 16348
rect 12221 16288 12285 16292
rect 12301 16348 12365 16352
rect 12301 16292 12305 16348
rect 12305 16292 12361 16348
rect 12361 16292 12365 16348
rect 12301 16288 12365 16292
rect 19835 16348 19899 16352
rect 19835 16292 19839 16348
rect 19839 16292 19895 16348
rect 19895 16292 19899 16348
rect 19835 16288 19899 16292
rect 19915 16348 19979 16352
rect 19915 16292 19919 16348
rect 19919 16292 19975 16348
rect 19975 16292 19979 16348
rect 19915 16288 19979 16292
rect 19995 16348 20059 16352
rect 19995 16292 19999 16348
rect 19999 16292 20055 16348
rect 20055 16292 20059 16348
rect 19995 16288 20059 16292
rect 20075 16348 20139 16352
rect 20075 16292 20079 16348
rect 20079 16292 20135 16348
rect 20135 16292 20139 16348
rect 20075 16288 20139 16292
rect 27609 16348 27673 16352
rect 27609 16292 27613 16348
rect 27613 16292 27669 16348
rect 27669 16292 27673 16348
rect 27609 16288 27673 16292
rect 27689 16348 27753 16352
rect 27689 16292 27693 16348
rect 27693 16292 27749 16348
rect 27749 16292 27753 16348
rect 27689 16288 27753 16292
rect 27769 16348 27833 16352
rect 27769 16292 27773 16348
rect 27773 16292 27829 16348
rect 27829 16292 27833 16348
rect 27769 16288 27833 16292
rect 27849 16348 27913 16352
rect 27849 16292 27853 16348
rect 27853 16292 27909 16348
rect 27909 16292 27913 16348
rect 27849 16288 27913 16292
rect 8174 15804 8238 15808
rect 8174 15748 8178 15804
rect 8178 15748 8234 15804
rect 8234 15748 8238 15804
rect 8174 15744 8238 15748
rect 8254 15804 8318 15808
rect 8254 15748 8258 15804
rect 8258 15748 8314 15804
rect 8314 15748 8318 15804
rect 8254 15744 8318 15748
rect 8334 15804 8398 15808
rect 8334 15748 8338 15804
rect 8338 15748 8394 15804
rect 8394 15748 8398 15804
rect 8334 15744 8398 15748
rect 8414 15804 8478 15808
rect 8414 15748 8418 15804
rect 8418 15748 8474 15804
rect 8474 15748 8478 15804
rect 8414 15744 8478 15748
rect 15948 15804 16012 15808
rect 15948 15748 15952 15804
rect 15952 15748 16008 15804
rect 16008 15748 16012 15804
rect 15948 15744 16012 15748
rect 16028 15804 16092 15808
rect 16028 15748 16032 15804
rect 16032 15748 16088 15804
rect 16088 15748 16092 15804
rect 16028 15744 16092 15748
rect 16108 15804 16172 15808
rect 16108 15748 16112 15804
rect 16112 15748 16168 15804
rect 16168 15748 16172 15804
rect 16108 15744 16172 15748
rect 16188 15804 16252 15808
rect 16188 15748 16192 15804
rect 16192 15748 16248 15804
rect 16248 15748 16252 15804
rect 16188 15744 16252 15748
rect 23722 15804 23786 15808
rect 23722 15748 23726 15804
rect 23726 15748 23782 15804
rect 23782 15748 23786 15804
rect 23722 15744 23786 15748
rect 23802 15804 23866 15808
rect 23802 15748 23806 15804
rect 23806 15748 23862 15804
rect 23862 15748 23866 15804
rect 23802 15744 23866 15748
rect 23882 15804 23946 15808
rect 23882 15748 23886 15804
rect 23886 15748 23942 15804
rect 23942 15748 23946 15804
rect 23882 15744 23946 15748
rect 23962 15804 24026 15808
rect 23962 15748 23966 15804
rect 23966 15748 24022 15804
rect 24022 15748 24026 15804
rect 23962 15744 24026 15748
rect 31496 15804 31560 15808
rect 31496 15748 31500 15804
rect 31500 15748 31556 15804
rect 31556 15748 31560 15804
rect 31496 15744 31560 15748
rect 31576 15804 31640 15808
rect 31576 15748 31580 15804
rect 31580 15748 31636 15804
rect 31636 15748 31640 15804
rect 31576 15744 31640 15748
rect 31656 15804 31720 15808
rect 31656 15748 31660 15804
rect 31660 15748 31716 15804
rect 31716 15748 31720 15804
rect 31656 15744 31720 15748
rect 31736 15804 31800 15808
rect 31736 15748 31740 15804
rect 31740 15748 31796 15804
rect 31796 15748 31800 15804
rect 31736 15744 31800 15748
rect 4287 15260 4351 15264
rect 4287 15204 4291 15260
rect 4291 15204 4347 15260
rect 4347 15204 4351 15260
rect 4287 15200 4351 15204
rect 4367 15260 4431 15264
rect 4367 15204 4371 15260
rect 4371 15204 4427 15260
rect 4427 15204 4431 15260
rect 4367 15200 4431 15204
rect 4447 15260 4511 15264
rect 4447 15204 4451 15260
rect 4451 15204 4507 15260
rect 4507 15204 4511 15260
rect 4447 15200 4511 15204
rect 4527 15260 4591 15264
rect 4527 15204 4531 15260
rect 4531 15204 4587 15260
rect 4587 15204 4591 15260
rect 4527 15200 4591 15204
rect 12061 15260 12125 15264
rect 12061 15204 12065 15260
rect 12065 15204 12121 15260
rect 12121 15204 12125 15260
rect 12061 15200 12125 15204
rect 12141 15260 12205 15264
rect 12141 15204 12145 15260
rect 12145 15204 12201 15260
rect 12201 15204 12205 15260
rect 12141 15200 12205 15204
rect 12221 15260 12285 15264
rect 12221 15204 12225 15260
rect 12225 15204 12281 15260
rect 12281 15204 12285 15260
rect 12221 15200 12285 15204
rect 12301 15260 12365 15264
rect 12301 15204 12305 15260
rect 12305 15204 12361 15260
rect 12361 15204 12365 15260
rect 12301 15200 12365 15204
rect 19835 15260 19899 15264
rect 19835 15204 19839 15260
rect 19839 15204 19895 15260
rect 19895 15204 19899 15260
rect 19835 15200 19899 15204
rect 19915 15260 19979 15264
rect 19915 15204 19919 15260
rect 19919 15204 19975 15260
rect 19975 15204 19979 15260
rect 19915 15200 19979 15204
rect 19995 15260 20059 15264
rect 19995 15204 19999 15260
rect 19999 15204 20055 15260
rect 20055 15204 20059 15260
rect 19995 15200 20059 15204
rect 20075 15260 20139 15264
rect 20075 15204 20079 15260
rect 20079 15204 20135 15260
rect 20135 15204 20139 15260
rect 20075 15200 20139 15204
rect 27609 15260 27673 15264
rect 27609 15204 27613 15260
rect 27613 15204 27669 15260
rect 27669 15204 27673 15260
rect 27609 15200 27673 15204
rect 27689 15260 27753 15264
rect 27689 15204 27693 15260
rect 27693 15204 27749 15260
rect 27749 15204 27753 15260
rect 27689 15200 27753 15204
rect 27769 15260 27833 15264
rect 27769 15204 27773 15260
rect 27773 15204 27829 15260
rect 27829 15204 27833 15260
rect 27769 15200 27833 15204
rect 27849 15260 27913 15264
rect 27849 15204 27853 15260
rect 27853 15204 27909 15260
rect 27909 15204 27913 15260
rect 27849 15200 27913 15204
rect 8174 14716 8238 14720
rect 8174 14660 8178 14716
rect 8178 14660 8234 14716
rect 8234 14660 8238 14716
rect 8174 14656 8238 14660
rect 8254 14716 8318 14720
rect 8254 14660 8258 14716
rect 8258 14660 8314 14716
rect 8314 14660 8318 14716
rect 8254 14656 8318 14660
rect 8334 14716 8398 14720
rect 8334 14660 8338 14716
rect 8338 14660 8394 14716
rect 8394 14660 8398 14716
rect 8334 14656 8398 14660
rect 8414 14716 8478 14720
rect 8414 14660 8418 14716
rect 8418 14660 8474 14716
rect 8474 14660 8478 14716
rect 8414 14656 8478 14660
rect 15948 14716 16012 14720
rect 15948 14660 15952 14716
rect 15952 14660 16008 14716
rect 16008 14660 16012 14716
rect 15948 14656 16012 14660
rect 16028 14716 16092 14720
rect 16028 14660 16032 14716
rect 16032 14660 16088 14716
rect 16088 14660 16092 14716
rect 16028 14656 16092 14660
rect 16108 14716 16172 14720
rect 16108 14660 16112 14716
rect 16112 14660 16168 14716
rect 16168 14660 16172 14716
rect 16108 14656 16172 14660
rect 16188 14716 16252 14720
rect 16188 14660 16192 14716
rect 16192 14660 16248 14716
rect 16248 14660 16252 14716
rect 16188 14656 16252 14660
rect 23722 14716 23786 14720
rect 23722 14660 23726 14716
rect 23726 14660 23782 14716
rect 23782 14660 23786 14716
rect 23722 14656 23786 14660
rect 23802 14716 23866 14720
rect 23802 14660 23806 14716
rect 23806 14660 23862 14716
rect 23862 14660 23866 14716
rect 23802 14656 23866 14660
rect 23882 14716 23946 14720
rect 23882 14660 23886 14716
rect 23886 14660 23942 14716
rect 23942 14660 23946 14716
rect 23882 14656 23946 14660
rect 23962 14716 24026 14720
rect 23962 14660 23966 14716
rect 23966 14660 24022 14716
rect 24022 14660 24026 14716
rect 23962 14656 24026 14660
rect 31496 14716 31560 14720
rect 31496 14660 31500 14716
rect 31500 14660 31556 14716
rect 31556 14660 31560 14716
rect 31496 14656 31560 14660
rect 31576 14716 31640 14720
rect 31576 14660 31580 14716
rect 31580 14660 31636 14716
rect 31636 14660 31640 14716
rect 31576 14656 31640 14660
rect 31656 14716 31720 14720
rect 31656 14660 31660 14716
rect 31660 14660 31716 14716
rect 31716 14660 31720 14716
rect 31656 14656 31720 14660
rect 31736 14716 31800 14720
rect 31736 14660 31740 14716
rect 31740 14660 31796 14716
rect 31796 14660 31800 14716
rect 31736 14656 31800 14660
rect 4287 14172 4351 14176
rect 4287 14116 4291 14172
rect 4291 14116 4347 14172
rect 4347 14116 4351 14172
rect 4287 14112 4351 14116
rect 4367 14172 4431 14176
rect 4367 14116 4371 14172
rect 4371 14116 4427 14172
rect 4427 14116 4431 14172
rect 4367 14112 4431 14116
rect 4447 14172 4511 14176
rect 4447 14116 4451 14172
rect 4451 14116 4507 14172
rect 4507 14116 4511 14172
rect 4447 14112 4511 14116
rect 4527 14172 4591 14176
rect 4527 14116 4531 14172
rect 4531 14116 4587 14172
rect 4587 14116 4591 14172
rect 4527 14112 4591 14116
rect 12061 14172 12125 14176
rect 12061 14116 12065 14172
rect 12065 14116 12121 14172
rect 12121 14116 12125 14172
rect 12061 14112 12125 14116
rect 12141 14172 12205 14176
rect 12141 14116 12145 14172
rect 12145 14116 12201 14172
rect 12201 14116 12205 14172
rect 12141 14112 12205 14116
rect 12221 14172 12285 14176
rect 12221 14116 12225 14172
rect 12225 14116 12281 14172
rect 12281 14116 12285 14172
rect 12221 14112 12285 14116
rect 12301 14172 12365 14176
rect 12301 14116 12305 14172
rect 12305 14116 12361 14172
rect 12361 14116 12365 14172
rect 12301 14112 12365 14116
rect 19835 14172 19899 14176
rect 19835 14116 19839 14172
rect 19839 14116 19895 14172
rect 19895 14116 19899 14172
rect 19835 14112 19899 14116
rect 19915 14172 19979 14176
rect 19915 14116 19919 14172
rect 19919 14116 19975 14172
rect 19975 14116 19979 14172
rect 19915 14112 19979 14116
rect 19995 14172 20059 14176
rect 19995 14116 19999 14172
rect 19999 14116 20055 14172
rect 20055 14116 20059 14172
rect 19995 14112 20059 14116
rect 20075 14172 20139 14176
rect 20075 14116 20079 14172
rect 20079 14116 20135 14172
rect 20135 14116 20139 14172
rect 20075 14112 20139 14116
rect 27609 14172 27673 14176
rect 27609 14116 27613 14172
rect 27613 14116 27669 14172
rect 27669 14116 27673 14172
rect 27609 14112 27673 14116
rect 27689 14172 27753 14176
rect 27689 14116 27693 14172
rect 27693 14116 27749 14172
rect 27749 14116 27753 14172
rect 27689 14112 27753 14116
rect 27769 14172 27833 14176
rect 27769 14116 27773 14172
rect 27773 14116 27829 14172
rect 27829 14116 27833 14172
rect 27769 14112 27833 14116
rect 27849 14172 27913 14176
rect 27849 14116 27853 14172
rect 27853 14116 27909 14172
rect 27909 14116 27913 14172
rect 27849 14112 27913 14116
rect 8174 13628 8238 13632
rect 8174 13572 8178 13628
rect 8178 13572 8234 13628
rect 8234 13572 8238 13628
rect 8174 13568 8238 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 15948 13628 16012 13632
rect 15948 13572 15952 13628
rect 15952 13572 16008 13628
rect 16008 13572 16012 13628
rect 15948 13568 16012 13572
rect 16028 13628 16092 13632
rect 16028 13572 16032 13628
rect 16032 13572 16088 13628
rect 16088 13572 16092 13628
rect 16028 13568 16092 13572
rect 16108 13628 16172 13632
rect 16108 13572 16112 13628
rect 16112 13572 16168 13628
rect 16168 13572 16172 13628
rect 16108 13568 16172 13572
rect 16188 13628 16252 13632
rect 16188 13572 16192 13628
rect 16192 13572 16248 13628
rect 16248 13572 16252 13628
rect 16188 13568 16252 13572
rect 23722 13628 23786 13632
rect 23722 13572 23726 13628
rect 23726 13572 23782 13628
rect 23782 13572 23786 13628
rect 23722 13568 23786 13572
rect 23802 13628 23866 13632
rect 23802 13572 23806 13628
rect 23806 13572 23862 13628
rect 23862 13572 23866 13628
rect 23802 13568 23866 13572
rect 23882 13628 23946 13632
rect 23882 13572 23886 13628
rect 23886 13572 23942 13628
rect 23942 13572 23946 13628
rect 23882 13568 23946 13572
rect 23962 13628 24026 13632
rect 23962 13572 23966 13628
rect 23966 13572 24022 13628
rect 24022 13572 24026 13628
rect 23962 13568 24026 13572
rect 31496 13628 31560 13632
rect 31496 13572 31500 13628
rect 31500 13572 31556 13628
rect 31556 13572 31560 13628
rect 31496 13568 31560 13572
rect 31576 13628 31640 13632
rect 31576 13572 31580 13628
rect 31580 13572 31636 13628
rect 31636 13572 31640 13628
rect 31576 13568 31640 13572
rect 31656 13628 31720 13632
rect 31656 13572 31660 13628
rect 31660 13572 31716 13628
rect 31716 13572 31720 13628
rect 31656 13568 31720 13572
rect 31736 13628 31800 13632
rect 31736 13572 31740 13628
rect 31740 13572 31796 13628
rect 31796 13572 31800 13628
rect 31736 13568 31800 13572
rect 4287 13084 4351 13088
rect 4287 13028 4291 13084
rect 4291 13028 4347 13084
rect 4347 13028 4351 13084
rect 4287 13024 4351 13028
rect 4367 13084 4431 13088
rect 4367 13028 4371 13084
rect 4371 13028 4427 13084
rect 4427 13028 4431 13084
rect 4367 13024 4431 13028
rect 4447 13084 4511 13088
rect 4447 13028 4451 13084
rect 4451 13028 4507 13084
rect 4507 13028 4511 13084
rect 4447 13024 4511 13028
rect 4527 13084 4591 13088
rect 4527 13028 4531 13084
rect 4531 13028 4587 13084
rect 4587 13028 4591 13084
rect 4527 13024 4591 13028
rect 12061 13084 12125 13088
rect 12061 13028 12065 13084
rect 12065 13028 12121 13084
rect 12121 13028 12125 13084
rect 12061 13024 12125 13028
rect 12141 13084 12205 13088
rect 12141 13028 12145 13084
rect 12145 13028 12201 13084
rect 12201 13028 12205 13084
rect 12141 13024 12205 13028
rect 12221 13084 12285 13088
rect 12221 13028 12225 13084
rect 12225 13028 12281 13084
rect 12281 13028 12285 13084
rect 12221 13024 12285 13028
rect 12301 13084 12365 13088
rect 12301 13028 12305 13084
rect 12305 13028 12361 13084
rect 12361 13028 12365 13084
rect 12301 13024 12365 13028
rect 19835 13084 19899 13088
rect 19835 13028 19839 13084
rect 19839 13028 19895 13084
rect 19895 13028 19899 13084
rect 19835 13024 19899 13028
rect 19915 13084 19979 13088
rect 19915 13028 19919 13084
rect 19919 13028 19975 13084
rect 19975 13028 19979 13084
rect 19915 13024 19979 13028
rect 19995 13084 20059 13088
rect 19995 13028 19999 13084
rect 19999 13028 20055 13084
rect 20055 13028 20059 13084
rect 19995 13024 20059 13028
rect 20075 13084 20139 13088
rect 20075 13028 20079 13084
rect 20079 13028 20135 13084
rect 20135 13028 20139 13084
rect 20075 13024 20139 13028
rect 27609 13084 27673 13088
rect 27609 13028 27613 13084
rect 27613 13028 27669 13084
rect 27669 13028 27673 13084
rect 27609 13024 27673 13028
rect 27689 13084 27753 13088
rect 27689 13028 27693 13084
rect 27693 13028 27749 13084
rect 27749 13028 27753 13084
rect 27689 13024 27753 13028
rect 27769 13084 27833 13088
rect 27769 13028 27773 13084
rect 27773 13028 27829 13084
rect 27829 13028 27833 13084
rect 27769 13024 27833 13028
rect 27849 13084 27913 13088
rect 27849 13028 27853 13084
rect 27853 13028 27909 13084
rect 27909 13028 27913 13084
rect 27849 13024 27913 13028
rect 8174 12540 8238 12544
rect 8174 12484 8178 12540
rect 8178 12484 8234 12540
rect 8234 12484 8238 12540
rect 8174 12480 8238 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 15948 12540 16012 12544
rect 15948 12484 15952 12540
rect 15952 12484 16008 12540
rect 16008 12484 16012 12540
rect 15948 12480 16012 12484
rect 16028 12540 16092 12544
rect 16028 12484 16032 12540
rect 16032 12484 16088 12540
rect 16088 12484 16092 12540
rect 16028 12480 16092 12484
rect 16108 12540 16172 12544
rect 16108 12484 16112 12540
rect 16112 12484 16168 12540
rect 16168 12484 16172 12540
rect 16108 12480 16172 12484
rect 16188 12540 16252 12544
rect 16188 12484 16192 12540
rect 16192 12484 16248 12540
rect 16248 12484 16252 12540
rect 16188 12480 16252 12484
rect 23722 12540 23786 12544
rect 23722 12484 23726 12540
rect 23726 12484 23782 12540
rect 23782 12484 23786 12540
rect 23722 12480 23786 12484
rect 23802 12540 23866 12544
rect 23802 12484 23806 12540
rect 23806 12484 23862 12540
rect 23862 12484 23866 12540
rect 23802 12480 23866 12484
rect 23882 12540 23946 12544
rect 23882 12484 23886 12540
rect 23886 12484 23942 12540
rect 23942 12484 23946 12540
rect 23882 12480 23946 12484
rect 23962 12540 24026 12544
rect 23962 12484 23966 12540
rect 23966 12484 24022 12540
rect 24022 12484 24026 12540
rect 23962 12480 24026 12484
rect 31496 12540 31560 12544
rect 31496 12484 31500 12540
rect 31500 12484 31556 12540
rect 31556 12484 31560 12540
rect 31496 12480 31560 12484
rect 31576 12540 31640 12544
rect 31576 12484 31580 12540
rect 31580 12484 31636 12540
rect 31636 12484 31640 12540
rect 31576 12480 31640 12484
rect 31656 12540 31720 12544
rect 31656 12484 31660 12540
rect 31660 12484 31716 12540
rect 31716 12484 31720 12540
rect 31656 12480 31720 12484
rect 31736 12540 31800 12544
rect 31736 12484 31740 12540
rect 31740 12484 31796 12540
rect 31796 12484 31800 12540
rect 31736 12480 31800 12484
rect 4287 11996 4351 12000
rect 4287 11940 4291 11996
rect 4291 11940 4347 11996
rect 4347 11940 4351 11996
rect 4287 11936 4351 11940
rect 4367 11996 4431 12000
rect 4367 11940 4371 11996
rect 4371 11940 4427 11996
rect 4427 11940 4431 11996
rect 4367 11936 4431 11940
rect 4447 11996 4511 12000
rect 4447 11940 4451 11996
rect 4451 11940 4507 11996
rect 4507 11940 4511 11996
rect 4447 11936 4511 11940
rect 4527 11996 4591 12000
rect 4527 11940 4531 11996
rect 4531 11940 4587 11996
rect 4587 11940 4591 11996
rect 4527 11936 4591 11940
rect 12061 11996 12125 12000
rect 12061 11940 12065 11996
rect 12065 11940 12121 11996
rect 12121 11940 12125 11996
rect 12061 11936 12125 11940
rect 12141 11996 12205 12000
rect 12141 11940 12145 11996
rect 12145 11940 12201 11996
rect 12201 11940 12205 11996
rect 12141 11936 12205 11940
rect 12221 11996 12285 12000
rect 12221 11940 12225 11996
rect 12225 11940 12281 11996
rect 12281 11940 12285 11996
rect 12221 11936 12285 11940
rect 12301 11996 12365 12000
rect 12301 11940 12305 11996
rect 12305 11940 12361 11996
rect 12361 11940 12365 11996
rect 12301 11936 12365 11940
rect 19835 11996 19899 12000
rect 19835 11940 19839 11996
rect 19839 11940 19895 11996
rect 19895 11940 19899 11996
rect 19835 11936 19899 11940
rect 19915 11996 19979 12000
rect 19915 11940 19919 11996
rect 19919 11940 19975 11996
rect 19975 11940 19979 11996
rect 19915 11936 19979 11940
rect 19995 11996 20059 12000
rect 19995 11940 19999 11996
rect 19999 11940 20055 11996
rect 20055 11940 20059 11996
rect 19995 11936 20059 11940
rect 20075 11996 20139 12000
rect 20075 11940 20079 11996
rect 20079 11940 20135 11996
rect 20135 11940 20139 11996
rect 20075 11936 20139 11940
rect 27609 11996 27673 12000
rect 27609 11940 27613 11996
rect 27613 11940 27669 11996
rect 27669 11940 27673 11996
rect 27609 11936 27673 11940
rect 27689 11996 27753 12000
rect 27689 11940 27693 11996
rect 27693 11940 27749 11996
rect 27749 11940 27753 11996
rect 27689 11936 27753 11940
rect 27769 11996 27833 12000
rect 27769 11940 27773 11996
rect 27773 11940 27829 11996
rect 27829 11940 27833 11996
rect 27769 11936 27833 11940
rect 27849 11996 27913 12000
rect 27849 11940 27853 11996
rect 27853 11940 27909 11996
rect 27909 11940 27913 11996
rect 27849 11936 27913 11940
rect 8174 11452 8238 11456
rect 8174 11396 8178 11452
rect 8178 11396 8234 11452
rect 8234 11396 8238 11452
rect 8174 11392 8238 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 15948 11452 16012 11456
rect 15948 11396 15952 11452
rect 15952 11396 16008 11452
rect 16008 11396 16012 11452
rect 15948 11392 16012 11396
rect 16028 11452 16092 11456
rect 16028 11396 16032 11452
rect 16032 11396 16088 11452
rect 16088 11396 16092 11452
rect 16028 11392 16092 11396
rect 16108 11452 16172 11456
rect 16108 11396 16112 11452
rect 16112 11396 16168 11452
rect 16168 11396 16172 11452
rect 16108 11392 16172 11396
rect 16188 11452 16252 11456
rect 16188 11396 16192 11452
rect 16192 11396 16248 11452
rect 16248 11396 16252 11452
rect 16188 11392 16252 11396
rect 23722 11452 23786 11456
rect 23722 11396 23726 11452
rect 23726 11396 23782 11452
rect 23782 11396 23786 11452
rect 23722 11392 23786 11396
rect 23802 11452 23866 11456
rect 23802 11396 23806 11452
rect 23806 11396 23862 11452
rect 23862 11396 23866 11452
rect 23802 11392 23866 11396
rect 23882 11452 23946 11456
rect 23882 11396 23886 11452
rect 23886 11396 23942 11452
rect 23942 11396 23946 11452
rect 23882 11392 23946 11396
rect 23962 11452 24026 11456
rect 23962 11396 23966 11452
rect 23966 11396 24022 11452
rect 24022 11396 24026 11452
rect 23962 11392 24026 11396
rect 31496 11452 31560 11456
rect 31496 11396 31500 11452
rect 31500 11396 31556 11452
rect 31556 11396 31560 11452
rect 31496 11392 31560 11396
rect 31576 11452 31640 11456
rect 31576 11396 31580 11452
rect 31580 11396 31636 11452
rect 31636 11396 31640 11452
rect 31576 11392 31640 11396
rect 31656 11452 31720 11456
rect 31656 11396 31660 11452
rect 31660 11396 31716 11452
rect 31716 11396 31720 11452
rect 31656 11392 31720 11396
rect 31736 11452 31800 11456
rect 31736 11396 31740 11452
rect 31740 11396 31796 11452
rect 31796 11396 31800 11452
rect 31736 11392 31800 11396
rect 4287 10908 4351 10912
rect 4287 10852 4291 10908
rect 4291 10852 4347 10908
rect 4347 10852 4351 10908
rect 4287 10848 4351 10852
rect 4367 10908 4431 10912
rect 4367 10852 4371 10908
rect 4371 10852 4427 10908
rect 4427 10852 4431 10908
rect 4367 10848 4431 10852
rect 4447 10908 4511 10912
rect 4447 10852 4451 10908
rect 4451 10852 4507 10908
rect 4507 10852 4511 10908
rect 4447 10848 4511 10852
rect 4527 10908 4591 10912
rect 4527 10852 4531 10908
rect 4531 10852 4587 10908
rect 4587 10852 4591 10908
rect 4527 10848 4591 10852
rect 12061 10908 12125 10912
rect 12061 10852 12065 10908
rect 12065 10852 12121 10908
rect 12121 10852 12125 10908
rect 12061 10848 12125 10852
rect 12141 10908 12205 10912
rect 12141 10852 12145 10908
rect 12145 10852 12201 10908
rect 12201 10852 12205 10908
rect 12141 10848 12205 10852
rect 12221 10908 12285 10912
rect 12221 10852 12225 10908
rect 12225 10852 12281 10908
rect 12281 10852 12285 10908
rect 12221 10848 12285 10852
rect 12301 10908 12365 10912
rect 12301 10852 12305 10908
rect 12305 10852 12361 10908
rect 12361 10852 12365 10908
rect 12301 10848 12365 10852
rect 19835 10908 19899 10912
rect 19835 10852 19839 10908
rect 19839 10852 19895 10908
rect 19895 10852 19899 10908
rect 19835 10848 19899 10852
rect 19915 10908 19979 10912
rect 19915 10852 19919 10908
rect 19919 10852 19975 10908
rect 19975 10852 19979 10908
rect 19915 10848 19979 10852
rect 19995 10908 20059 10912
rect 19995 10852 19999 10908
rect 19999 10852 20055 10908
rect 20055 10852 20059 10908
rect 19995 10848 20059 10852
rect 20075 10908 20139 10912
rect 20075 10852 20079 10908
rect 20079 10852 20135 10908
rect 20135 10852 20139 10908
rect 20075 10848 20139 10852
rect 27609 10908 27673 10912
rect 27609 10852 27613 10908
rect 27613 10852 27669 10908
rect 27669 10852 27673 10908
rect 27609 10848 27673 10852
rect 27689 10908 27753 10912
rect 27689 10852 27693 10908
rect 27693 10852 27749 10908
rect 27749 10852 27753 10908
rect 27689 10848 27753 10852
rect 27769 10908 27833 10912
rect 27769 10852 27773 10908
rect 27773 10852 27829 10908
rect 27829 10852 27833 10908
rect 27769 10848 27833 10852
rect 27849 10908 27913 10912
rect 27849 10852 27853 10908
rect 27853 10852 27909 10908
rect 27909 10852 27913 10908
rect 27849 10848 27913 10852
rect 8174 10364 8238 10368
rect 8174 10308 8178 10364
rect 8178 10308 8234 10364
rect 8234 10308 8238 10364
rect 8174 10304 8238 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 15948 10364 16012 10368
rect 15948 10308 15952 10364
rect 15952 10308 16008 10364
rect 16008 10308 16012 10364
rect 15948 10304 16012 10308
rect 16028 10364 16092 10368
rect 16028 10308 16032 10364
rect 16032 10308 16088 10364
rect 16088 10308 16092 10364
rect 16028 10304 16092 10308
rect 16108 10364 16172 10368
rect 16108 10308 16112 10364
rect 16112 10308 16168 10364
rect 16168 10308 16172 10364
rect 16108 10304 16172 10308
rect 16188 10364 16252 10368
rect 16188 10308 16192 10364
rect 16192 10308 16248 10364
rect 16248 10308 16252 10364
rect 16188 10304 16252 10308
rect 23722 10364 23786 10368
rect 23722 10308 23726 10364
rect 23726 10308 23782 10364
rect 23782 10308 23786 10364
rect 23722 10304 23786 10308
rect 23802 10364 23866 10368
rect 23802 10308 23806 10364
rect 23806 10308 23862 10364
rect 23862 10308 23866 10364
rect 23802 10304 23866 10308
rect 23882 10364 23946 10368
rect 23882 10308 23886 10364
rect 23886 10308 23942 10364
rect 23942 10308 23946 10364
rect 23882 10304 23946 10308
rect 23962 10364 24026 10368
rect 23962 10308 23966 10364
rect 23966 10308 24022 10364
rect 24022 10308 24026 10364
rect 23962 10304 24026 10308
rect 31496 10364 31560 10368
rect 31496 10308 31500 10364
rect 31500 10308 31556 10364
rect 31556 10308 31560 10364
rect 31496 10304 31560 10308
rect 31576 10364 31640 10368
rect 31576 10308 31580 10364
rect 31580 10308 31636 10364
rect 31636 10308 31640 10364
rect 31576 10304 31640 10308
rect 31656 10364 31720 10368
rect 31656 10308 31660 10364
rect 31660 10308 31716 10364
rect 31716 10308 31720 10364
rect 31656 10304 31720 10308
rect 31736 10364 31800 10368
rect 31736 10308 31740 10364
rect 31740 10308 31796 10364
rect 31796 10308 31800 10364
rect 31736 10304 31800 10308
rect 4287 9820 4351 9824
rect 4287 9764 4291 9820
rect 4291 9764 4347 9820
rect 4347 9764 4351 9820
rect 4287 9760 4351 9764
rect 4367 9820 4431 9824
rect 4367 9764 4371 9820
rect 4371 9764 4427 9820
rect 4427 9764 4431 9820
rect 4367 9760 4431 9764
rect 4447 9820 4511 9824
rect 4447 9764 4451 9820
rect 4451 9764 4507 9820
rect 4507 9764 4511 9820
rect 4447 9760 4511 9764
rect 4527 9820 4591 9824
rect 4527 9764 4531 9820
rect 4531 9764 4587 9820
rect 4587 9764 4591 9820
rect 4527 9760 4591 9764
rect 12061 9820 12125 9824
rect 12061 9764 12065 9820
rect 12065 9764 12121 9820
rect 12121 9764 12125 9820
rect 12061 9760 12125 9764
rect 12141 9820 12205 9824
rect 12141 9764 12145 9820
rect 12145 9764 12201 9820
rect 12201 9764 12205 9820
rect 12141 9760 12205 9764
rect 12221 9820 12285 9824
rect 12221 9764 12225 9820
rect 12225 9764 12281 9820
rect 12281 9764 12285 9820
rect 12221 9760 12285 9764
rect 12301 9820 12365 9824
rect 12301 9764 12305 9820
rect 12305 9764 12361 9820
rect 12361 9764 12365 9820
rect 12301 9760 12365 9764
rect 19835 9820 19899 9824
rect 19835 9764 19839 9820
rect 19839 9764 19895 9820
rect 19895 9764 19899 9820
rect 19835 9760 19899 9764
rect 19915 9820 19979 9824
rect 19915 9764 19919 9820
rect 19919 9764 19975 9820
rect 19975 9764 19979 9820
rect 19915 9760 19979 9764
rect 19995 9820 20059 9824
rect 19995 9764 19999 9820
rect 19999 9764 20055 9820
rect 20055 9764 20059 9820
rect 19995 9760 20059 9764
rect 20075 9820 20139 9824
rect 20075 9764 20079 9820
rect 20079 9764 20135 9820
rect 20135 9764 20139 9820
rect 20075 9760 20139 9764
rect 27609 9820 27673 9824
rect 27609 9764 27613 9820
rect 27613 9764 27669 9820
rect 27669 9764 27673 9820
rect 27609 9760 27673 9764
rect 27689 9820 27753 9824
rect 27689 9764 27693 9820
rect 27693 9764 27749 9820
rect 27749 9764 27753 9820
rect 27689 9760 27753 9764
rect 27769 9820 27833 9824
rect 27769 9764 27773 9820
rect 27773 9764 27829 9820
rect 27829 9764 27833 9820
rect 27769 9760 27833 9764
rect 27849 9820 27913 9824
rect 27849 9764 27853 9820
rect 27853 9764 27909 9820
rect 27909 9764 27913 9820
rect 27849 9760 27913 9764
rect 8174 9276 8238 9280
rect 8174 9220 8178 9276
rect 8178 9220 8234 9276
rect 8234 9220 8238 9276
rect 8174 9216 8238 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 15948 9276 16012 9280
rect 15948 9220 15952 9276
rect 15952 9220 16008 9276
rect 16008 9220 16012 9276
rect 15948 9216 16012 9220
rect 16028 9276 16092 9280
rect 16028 9220 16032 9276
rect 16032 9220 16088 9276
rect 16088 9220 16092 9276
rect 16028 9216 16092 9220
rect 16108 9276 16172 9280
rect 16108 9220 16112 9276
rect 16112 9220 16168 9276
rect 16168 9220 16172 9276
rect 16108 9216 16172 9220
rect 16188 9276 16252 9280
rect 16188 9220 16192 9276
rect 16192 9220 16248 9276
rect 16248 9220 16252 9276
rect 16188 9216 16252 9220
rect 23722 9276 23786 9280
rect 23722 9220 23726 9276
rect 23726 9220 23782 9276
rect 23782 9220 23786 9276
rect 23722 9216 23786 9220
rect 23802 9276 23866 9280
rect 23802 9220 23806 9276
rect 23806 9220 23862 9276
rect 23862 9220 23866 9276
rect 23802 9216 23866 9220
rect 23882 9276 23946 9280
rect 23882 9220 23886 9276
rect 23886 9220 23942 9276
rect 23942 9220 23946 9276
rect 23882 9216 23946 9220
rect 23962 9276 24026 9280
rect 23962 9220 23966 9276
rect 23966 9220 24022 9276
rect 24022 9220 24026 9276
rect 23962 9216 24026 9220
rect 31496 9276 31560 9280
rect 31496 9220 31500 9276
rect 31500 9220 31556 9276
rect 31556 9220 31560 9276
rect 31496 9216 31560 9220
rect 31576 9276 31640 9280
rect 31576 9220 31580 9276
rect 31580 9220 31636 9276
rect 31636 9220 31640 9276
rect 31576 9216 31640 9220
rect 31656 9276 31720 9280
rect 31656 9220 31660 9276
rect 31660 9220 31716 9276
rect 31716 9220 31720 9276
rect 31656 9216 31720 9220
rect 31736 9276 31800 9280
rect 31736 9220 31740 9276
rect 31740 9220 31796 9276
rect 31796 9220 31800 9276
rect 31736 9216 31800 9220
rect 4287 8732 4351 8736
rect 4287 8676 4291 8732
rect 4291 8676 4347 8732
rect 4347 8676 4351 8732
rect 4287 8672 4351 8676
rect 4367 8732 4431 8736
rect 4367 8676 4371 8732
rect 4371 8676 4427 8732
rect 4427 8676 4431 8732
rect 4367 8672 4431 8676
rect 4447 8732 4511 8736
rect 4447 8676 4451 8732
rect 4451 8676 4507 8732
rect 4507 8676 4511 8732
rect 4447 8672 4511 8676
rect 4527 8732 4591 8736
rect 4527 8676 4531 8732
rect 4531 8676 4587 8732
rect 4587 8676 4591 8732
rect 4527 8672 4591 8676
rect 12061 8732 12125 8736
rect 12061 8676 12065 8732
rect 12065 8676 12121 8732
rect 12121 8676 12125 8732
rect 12061 8672 12125 8676
rect 12141 8732 12205 8736
rect 12141 8676 12145 8732
rect 12145 8676 12201 8732
rect 12201 8676 12205 8732
rect 12141 8672 12205 8676
rect 12221 8732 12285 8736
rect 12221 8676 12225 8732
rect 12225 8676 12281 8732
rect 12281 8676 12285 8732
rect 12221 8672 12285 8676
rect 12301 8732 12365 8736
rect 12301 8676 12305 8732
rect 12305 8676 12361 8732
rect 12361 8676 12365 8732
rect 12301 8672 12365 8676
rect 19835 8732 19899 8736
rect 19835 8676 19839 8732
rect 19839 8676 19895 8732
rect 19895 8676 19899 8732
rect 19835 8672 19899 8676
rect 19915 8732 19979 8736
rect 19915 8676 19919 8732
rect 19919 8676 19975 8732
rect 19975 8676 19979 8732
rect 19915 8672 19979 8676
rect 19995 8732 20059 8736
rect 19995 8676 19999 8732
rect 19999 8676 20055 8732
rect 20055 8676 20059 8732
rect 19995 8672 20059 8676
rect 20075 8732 20139 8736
rect 20075 8676 20079 8732
rect 20079 8676 20135 8732
rect 20135 8676 20139 8732
rect 20075 8672 20139 8676
rect 27609 8732 27673 8736
rect 27609 8676 27613 8732
rect 27613 8676 27669 8732
rect 27669 8676 27673 8732
rect 27609 8672 27673 8676
rect 27689 8732 27753 8736
rect 27689 8676 27693 8732
rect 27693 8676 27749 8732
rect 27749 8676 27753 8732
rect 27689 8672 27753 8676
rect 27769 8732 27833 8736
rect 27769 8676 27773 8732
rect 27773 8676 27829 8732
rect 27829 8676 27833 8732
rect 27769 8672 27833 8676
rect 27849 8732 27913 8736
rect 27849 8676 27853 8732
rect 27853 8676 27909 8732
rect 27909 8676 27913 8732
rect 27849 8672 27913 8676
rect 8174 8188 8238 8192
rect 8174 8132 8178 8188
rect 8178 8132 8234 8188
rect 8234 8132 8238 8188
rect 8174 8128 8238 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 15948 8188 16012 8192
rect 15948 8132 15952 8188
rect 15952 8132 16008 8188
rect 16008 8132 16012 8188
rect 15948 8128 16012 8132
rect 16028 8188 16092 8192
rect 16028 8132 16032 8188
rect 16032 8132 16088 8188
rect 16088 8132 16092 8188
rect 16028 8128 16092 8132
rect 16108 8188 16172 8192
rect 16108 8132 16112 8188
rect 16112 8132 16168 8188
rect 16168 8132 16172 8188
rect 16108 8128 16172 8132
rect 16188 8188 16252 8192
rect 16188 8132 16192 8188
rect 16192 8132 16248 8188
rect 16248 8132 16252 8188
rect 16188 8128 16252 8132
rect 23722 8188 23786 8192
rect 23722 8132 23726 8188
rect 23726 8132 23782 8188
rect 23782 8132 23786 8188
rect 23722 8128 23786 8132
rect 23802 8188 23866 8192
rect 23802 8132 23806 8188
rect 23806 8132 23862 8188
rect 23862 8132 23866 8188
rect 23802 8128 23866 8132
rect 23882 8188 23946 8192
rect 23882 8132 23886 8188
rect 23886 8132 23942 8188
rect 23942 8132 23946 8188
rect 23882 8128 23946 8132
rect 23962 8188 24026 8192
rect 23962 8132 23966 8188
rect 23966 8132 24022 8188
rect 24022 8132 24026 8188
rect 23962 8128 24026 8132
rect 31496 8188 31560 8192
rect 31496 8132 31500 8188
rect 31500 8132 31556 8188
rect 31556 8132 31560 8188
rect 31496 8128 31560 8132
rect 31576 8188 31640 8192
rect 31576 8132 31580 8188
rect 31580 8132 31636 8188
rect 31636 8132 31640 8188
rect 31576 8128 31640 8132
rect 31656 8188 31720 8192
rect 31656 8132 31660 8188
rect 31660 8132 31716 8188
rect 31716 8132 31720 8188
rect 31656 8128 31720 8132
rect 31736 8188 31800 8192
rect 31736 8132 31740 8188
rect 31740 8132 31796 8188
rect 31796 8132 31800 8188
rect 31736 8128 31800 8132
rect 4287 7644 4351 7648
rect 4287 7588 4291 7644
rect 4291 7588 4347 7644
rect 4347 7588 4351 7644
rect 4287 7584 4351 7588
rect 4367 7644 4431 7648
rect 4367 7588 4371 7644
rect 4371 7588 4427 7644
rect 4427 7588 4431 7644
rect 4367 7584 4431 7588
rect 4447 7644 4511 7648
rect 4447 7588 4451 7644
rect 4451 7588 4507 7644
rect 4507 7588 4511 7644
rect 4447 7584 4511 7588
rect 4527 7644 4591 7648
rect 4527 7588 4531 7644
rect 4531 7588 4587 7644
rect 4587 7588 4591 7644
rect 4527 7584 4591 7588
rect 12061 7644 12125 7648
rect 12061 7588 12065 7644
rect 12065 7588 12121 7644
rect 12121 7588 12125 7644
rect 12061 7584 12125 7588
rect 12141 7644 12205 7648
rect 12141 7588 12145 7644
rect 12145 7588 12201 7644
rect 12201 7588 12205 7644
rect 12141 7584 12205 7588
rect 12221 7644 12285 7648
rect 12221 7588 12225 7644
rect 12225 7588 12281 7644
rect 12281 7588 12285 7644
rect 12221 7584 12285 7588
rect 12301 7644 12365 7648
rect 12301 7588 12305 7644
rect 12305 7588 12361 7644
rect 12361 7588 12365 7644
rect 12301 7584 12365 7588
rect 19835 7644 19899 7648
rect 19835 7588 19839 7644
rect 19839 7588 19895 7644
rect 19895 7588 19899 7644
rect 19835 7584 19899 7588
rect 19915 7644 19979 7648
rect 19915 7588 19919 7644
rect 19919 7588 19975 7644
rect 19975 7588 19979 7644
rect 19915 7584 19979 7588
rect 19995 7644 20059 7648
rect 19995 7588 19999 7644
rect 19999 7588 20055 7644
rect 20055 7588 20059 7644
rect 19995 7584 20059 7588
rect 20075 7644 20139 7648
rect 20075 7588 20079 7644
rect 20079 7588 20135 7644
rect 20135 7588 20139 7644
rect 20075 7584 20139 7588
rect 27609 7644 27673 7648
rect 27609 7588 27613 7644
rect 27613 7588 27669 7644
rect 27669 7588 27673 7644
rect 27609 7584 27673 7588
rect 27689 7644 27753 7648
rect 27689 7588 27693 7644
rect 27693 7588 27749 7644
rect 27749 7588 27753 7644
rect 27689 7584 27753 7588
rect 27769 7644 27833 7648
rect 27769 7588 27773 7644
rect 27773 7588 27829 7644
rect 27829 7588 27833 7644
rect 27769 7584 27833 7588
rect 27849 7644 27913 7648
rect 27849 7588 27853 7644
rect 27853 7588 27909 7644
rect 27909 7588 27913 7644
rect 27849 7584 27913 7588
rect 8174 7100 8238 7104
rect 8174 7044 8178 7100
rect 8178 7044 8234 7100
rect 8234 7044 8238 7100
rect 8174 7040 8238 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 15948 7100 16012 7104
rect 15948 7044 15952 7100
rect 15952 7044 16008 7100
rect 16008 7044 16012 7100
rect 15948 7040 16012 7044
rect 16028 7100 16092 7104
rect 16028 7044 16032 7100
rect 16032 7044 16088 7100
rect 16088 7044 16092 7100
rect 16028 7040 16092 7044
rect 16108 7100 16172 7104
rect 16108 7044 16112 7100
rect 16112 7044 16168 7100
rect 16168 7044 16172 7100
rect 16108 7040 16172 7044
rect 16188 7100 16252 7104
rect 16188 7044 16192 7100
rect 16192 7044 16248 7100
rect 16248 7044 16252 7100
rect 16188 7040 16252 7044
rect 23722 7100 23786 7104
rect 23722 7044 23726 7100
rect 23726 7044 23782 7100
rect 23782 7044 23786 7100
rect 23722 7040 23786 7044
rect 23802 7100 23866 7104
rect 23802 7044 23806 7100
rect 23806 7044 23862 7100
rect 23862 7044 23866 7100
rect 23802 7040 23866 7044
rect 23882 7100 23946 7104
rect 23882 7044 23886 7100
rect 23886 7044 23942 7100
rect 23942 7044 23946 7100
rect 23882 7040 23946 7044
rect 23962 7100 24026 7104
rect 23962 7044 23966 7100
rect 23966 7044 24022 7100
rect 24022 7044 24026 7100
rect 23962 7040 24026 7044
rect 31496 7100 31560 7104
rect 31496 7044 31500 7100
rect 31500 7044 31556 7100
rect 31556 7044 31560 7100
rect 31496 7040 31560 7044
rect 31576 7100 31640 7104
rect 31576 7044 31580 7100
rect 31580 7044 31636 7100
rect 31636 7044 31640 7100
rect 31576 7040 31640 7044
rect 31656 7100 31720 7104
rect 31656 7044 31660 7100
rect 31660 7044 31716 7100
rect 31716 7044 31720 7100
rect 31656 7040 31720 7044
rect 31736 7100 31800 7104
rect 31736 7044 31740 7100
rect 31740 7044 31796 7100
rect 31796 7044 31800 7100
rect 31736 7040 31800 7044
rect 4287 6556 4351 6560
rect 4287 6500 4291 6556
rect 4291 6500 4347 6556
rect 4347 6500 4351 6556
rect 4287 6496 4351 6500
rect 4367 6556 4431 6560
rect 4367 6500 4371 6556
rect 4371 6500 4427 6556
rect 4427 6500 4431 6556
rect 4367 6496 4431 6500
rect 4447 6556 4511 6560
rect 4447 6500 4451 6556
rect 4451 6500 4507 6556
rect 4507 6500 4511 6556
rect 4447 6496 4511 6500
rect 4527 6556 4591 6560
rect 4527 6500 4531 6556
rect 4531 6500 4587 6556
rect 4587 6500 4591 6556
rect 4527 6496 4591 6500
rect 12061 6556 12125 6560
rect 12061 6500 12065 6556
rect 12065 6500 12121 6556
rect 12121 6500 12125 6556
rect 12061 6496 12125 6500
rect 12141 6556 12205 6560
rect 12141 6500 12145 6556
rect 12145 6500 12201 6556
rect 12201 6500 12205 6556
rect 12141 6496 12205 6500
rect 12221 6556 12285 6560
rect 12221 6500 12225 6556
rect 12225 6500 12281 6556
rect 12281 6500 12285 6556
rect 12221 6496 12285 6500
rect 12301 6556 12365 6560
rect 12301 6500 12305 6556
rect 12305 6500 12361 6556
rect 12361 6500 12365 6556
rect 12301 6496 12365 6500
rect 19835 6556 19899 6560
rect 19835 6500 19839 6556
rect 19839 6500 19895 6556
rect 19895 6500 19899 6556
rect 19835 6496 19899 6500
rect 19915 6556 19979 6560
rect 19915 6500 19919 6556
rect 19919 6500 19975 6556
rect 19975 6500 19979 6556
rect 19915 6496 19979 6500
rect 19995 6556 20059 6560
rect 19995 6500 19999 6556
rect 19999 6500 20055 6556
rect 20055 6500 20059 6556
rect 19995 6496 20059 6500
rect 20075 6556 20139 6560
rect 20075 6500 20079 6556
rect 20079 6500 20135 6556
rect 20135 6500 20139 6556
rect 20075 6496 20139 6500
rect 27609 6556 27673 6560
rect 27609 6500 27613 6556
rect 27613 6500 27669 6556
rect 27669 6500 27673 6556
rect 27609 6496 27673 6500
rect 27689 6556 27753 6560
rect 27689 6500 27693 6556
rect 27693 6500 27749 6556
rect 27749 6500 27753 6556
rect 27689 6496 27753 6500
rect 27769 6556 27833 6560
rect 27769 6500 27773 6556
rect 27773 6500 27829 6556
rect 27829 6500 27833 6556
rect 27769 6496 27833 6500
rect 27849 6556 27913 6560
rect 27849 6500 27853 6556
rect 27853 6500 27909 6556
rect 27909 6500 27913 6556
rect 27849 6496 27913 6500
rect 8174 6012 8238 6016
rect 8174 5956 8178 6012
rect 8178 5956 8234 6012
rect 8234 5956 8238 6012
rect 8174 5952 8238 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 15948 6012 16012 6016
rect 15948 5956 15952 6012
rect 15952 5956 16008 6012
rect 16008 5956 16012 6012
rect 15948 5952 16012 5956
rect 16028 6012 16092 6016
rect 16028 5956 16032 6012
rect 16032 5956 16088 6012
rect 16088 5956 16092 6012
rect 16028 5952 16092 5956
rect 16108 6012 16172 6016
rect 16108 5956 16112 6012
rect 16112 5956 16168 6012
rect 16168 5956 16172 6012
rect 16108 5952 16172 5956
rect 16188 6012 16252 6016
rect 16188 5956 16192 6012
rect 16192 5956 16248 6012
rect 16248 5956 16252 6012
rect 16188 5952 16252 5956
rect 23722 6012 23786 6016
rect 23722 5956 23726 6012
rect 23726 5956 23782 6012
rect 23782 5956 23786 6012
rect 23722 5952 23786 5956
rect 23802 6012 23866 6016
rect 23802 5956 23806 6012
rect 23806 5956 23862 6012
rect 23862 5956 23866 6012
rect 23802 5952 23866 5956
rect 23882 6012 23946 6016
rect 23882 5956 23886 6012
rect 23886 5956 23942 6012
rect 23942 5956 23946 6012
rect 23882 5952 23946 5956
rect 23962 6012 24026 6016
rect 23962 5956 23966 6012
rect 23966 5956 24022 6012
rect 24022 5956 24026 6012
rect 23962 5952 24026 5956
rect 31496 6012 31560 6016
rect 31496 5956 31500 6012
rect 31500 5956 31556 6012
rect 31556 5956 31560 6012
rect 31496 5952 31560 5956
rect 31576 6012 31640 6016
rect 31576 5956 31580 6012
rect 31580 5956 31636 6012
rect 31636 5956 31640 6012
rect 31576 5952 31640 5956
rect 31656 6012 31720 6016
rect 31656 5956 31660 6012
rect 31660 5956 31716 6012
rect 31716 5956 31720 6012
rect 31656 5952 31720 5956
rect 31736 6012 31800 6016
rect 31736 5956 31740 6012
rect 31740 5956 31796 6012
rect 31796 5956 31800 6012
rect 31736 5952 31800 5956
rect 4287 5468 4351 5472
rect 4287 5412 4291 5468
rect 4291 5412 4347 5468
rect 4347 5412 4351 5468
rect 4287 5408 4351 5412
rect 4367 5468 4431 5472
rect 4367 5412 4371 5468
rect 4371 5412 4427 5468
rect 4427 5412 4431 5468
rect 4367 5408 4431 5412
rect 4447 5468 4511 5472
rect 4447 5412 4451 5468
rect 4451 5412 4507 5468
rect 4507 5412 4511 5468
rect 4447 5408 4511 5412
rect 4527 5468 4591 5472
rect 4527 5412 4531 5468
rect 4531 5412 4587 5468
rect 4587 5412 4591 5468
rect 4527 5408 4591 5412
rect 12061 5468 12125 5472
rect 12061 5412 12065 5468
rect 12065 5412 12121 5468
rect 12121 5412 12125 5468
rect 12061 5408 12125 5412
rect 12141 5468 12205 5472
rect 12141 5412 12145 5468
rect 12145 5412 12201 5468
rect 12201 5412 12205 5468
rect 12141 5408 12205 5412
rect 12221 5468 12285 5472
rect 12221 5412 12225 5468
rect 12225 5412 12281 5468
rect 12281 5412 12285 5468
rect 12221 5408 12285 5412
rect 12301 5468 12365 5472
rect 12301 5412 12305 5468
rect 12305 5412 12361 5468
rect 12361 5412 12365 5468
rect 12301 5408 12365 5412
rect 19835 5468 19899 5472
rect 19835 5412 19839 5468
rect 19839 5412 19895 5468
rect 19895 5412 19899 5468
rect 19835 5408 19899 5412
rect 19915 5468 19979 5472
rect 19915 5412 19919 5468
rect 19919 5412 19975 5468
rect 19975 5412 19979 5468
rect 19915 5408 19979 5412
rect 19995 5468 20059 5472
rect 19995 5412 19999 5468
rect 19999 5412 20055 5468
rect 20055 5412 20059 5468
rect 19995 5408 20059 5412
rect 20075 5468 20139 5472
rect 20075 5412 20079 5468
rect 20079 5412 20135 5468
rect 20135 5412 20139 5468
rect 20075 5408 20139 5412
rect 27609 5468 27673 5472
rect 27609 5412 27613 5468
rect 27613 5412 27669 5468
rect 27669 5412 27673 5468
rect 27609 5408 27673 5412
rect 27689 5468 27753 5472
rect 27689 5412 27693 5468
rect 27693 5412 27749 5468
rect 27749 5412 27753 5468
rect 27689 5408 27753 5412
rect 27769 5468 27833 5472
rect 27769 5412 27773 5468
rect 27773 5412 27829 5468
rect 27829 5412 27833 5468
rect 27769 5408 27833 5412
rect 27849 5468 27913 5472
rect 27849 5412 27853 5468
rect 27853 5412 27909 5468
rect 27909 5412 27913 5468
rect 27849 5408 27913 5412
rect 8174 4924 8238 4928
rect 8174 4868 8178 4924
rect 8178 4868 8234 4924
rect 8234 4868 8238 4924
rect 8174 4864 8238 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 15948 4924 16012 4928
rect 15948 4868 15952 4924
rect 15952 4868 16008 4924
rect 16008 4868 16012 4924
rect 15948 4864 16012 4868
rect 16028 4924 16092 4928
rect 16028 4868 16032 4924
rect 16032 4868 16088 4924
rect 16088 4868 16092 4924
rect 16028 4864 16092 4868
rect 16108 4924 16172 4928
rect 16108 4868 16112 4924
rect 16112 4868 16168 4924
rect 16168 4868 16172 4924
rect 16108 4864 16172 4868
rect 16188 4924 16252 4928
rect 16188 4868 16192 4924
rect 16192 4868 16248 4924
rect 16248 4868 16252 4924
rect 16188 4864 16252 4868
rect 23722 4924 23786 4928
rect 23722 4868 23726 4924
rect 23726 4868 23782 4924
rect 23782 4868 23786 4924
rect 23722 4864 23786 4868
rect 23802 4924 23866 4928
rect 23802 4868 23806 4924
rect 23806 4868 23862 4924
rect 23862 4868 23866 4924
rect 23802 4864 23866 4868
rect 23882 4924 23946 4928
rect 23882 4868 23886 4924
rect 23886 4868 23942 4924
rect 23942 4868 23946 4924
rect 23882 4864 23946 4868
rect 23962 4924 24026 4928
rect 23962 4868 23966 4924
rect 23966 4868 24022 4924
rect 24022 4868 24026 4924
rect 23962 4864 24026 4868
rect 31496 4924 31560 4928
rect 31496 4868 31500 4924
rect 31500 4868 31556 4924
rect 31556 4868 31560 4924
rect 31496 4864 31560 4868
rect 31576 4924 31640 4928
rect 31576 4868 31580 4924
rect 31580 4868 31636 4924
rect 31636 4868 31640 4924
rect 31576 4864 31640 4868
rect 31656 4924 31720 4928
rect 31656 4868 31660 4924
rect 31660 4868 31716 4924
rect 31716 4868 31720 4924
rect 31656 4864 31720 4868
rect 31736 4924 31800 4928
rect 31736 4868 31740 4924
rect 31740 4868 31796 4924
rect 31796 4868 31800 4924
rect 31736 4864 31800 4868
rect 4287 4380 4351 4384
rect 4287 4324 4291 4380
rect 4291 4324 4347 4380
rect 4347 4324 4351 4380
rect 4287 4320 4351 4324
rect 4367 4380 4431 4384
rect 4367 4324 4371 4380
rect 4371 4324 4427 4380
rect 4427 4324 4431 4380
rect 4367 4320 4431 4324
rect 4447 4380 4511 4384
rect 4447 4324 4451 4380
rect 4451 4324 4507 4380
rect 4507 4324 4511 4380
rect 4447 4320 4511 4324
rect 4527 4380 4591 4384
rect 4527 4324 4531 4380
rect 4531 4324 4587 4380
rect 4587 4324 4591 4380
rect 4527 4320 4591 4324
rect 12061 4380 12125 4384
rect 12061 4324 12065 4380
rect 12065 4324 12121 4380
rect 12121 4324 12125 4380
rect 12061 4320 12125 4324
rect 12141 4380 12205 4384
rect 12141 4324 12145 4380
rect 12145 4324 12201 4380
rect 12201 4324 12205 4380
rect 12141 4320 12205 4324
rect 12221 4380 12285 4384
rect 12221 4324 12225 4380
rect 12225 4324 12281 4380
rect 12281 4324 12285 4380
rect 12221 4320 12285 4324
rect 12301 4380 12365 4384
rect 12301 4324 12305 4380
rect 12305 4324 12361 4380
rect 12361 4324 12365 4380
rect 12301 4320 12365 4324
rect 19835 4380 19899 4384
rect 19835 4324 19839 4380
rect 19839 4324 19895 4380
rect 19895 4324 19899 4380
rect 19835 4320 19899 4324
rect 19915 4380 19979 4384
rect 19915 4324 19919 4380
rect 19919 4324 19975 4380
rect 19975 4324 19979 4380
rect 19915 4320 19979 4324
rect 19995 4380 20059 4384
rect 19995 4324 19999 4380
rect 19999 4324 20055 4380
rect 20055 4324 20059 4380
rect 19995 4320 20059 4324
rect 20075 4380 20139 4384
rect 20075 4324 20079 4380
rect 20079 4324 20135 4380
rect 20135 4324 20139 4380
rect 20075 4320 20139 4324
rect 27609 4380 27673 4384
rect 27609 4324 27613 4380
rect 27613 4324 27669 4380
rect 27669 4324 27673 4380
rect 27609 4320 27673 4324
rect 27689 4380 27753 4384
rect 27689 4324 27693 4380
rect 27693 4324 27749 4380
rect 27749 4324 27753 4380
rect 27689 4320 27753 4324
rect 27769 4380 27833 4384
rect 27769 4324 27773 4380
rect 27773 4324 27829 4380
rect 27829 4324 27833 4380
rect 27769 4320 27833 4324
rect 27849 4380 27913 4384
rect 27849 4324 27853 4380
rect 27853 4324 27909 4380
rect 27909 4324 27913 4380
rect 27849 4320 27913 4324
rect 8174 3836 8238 3840
rect 8174 3780 8178 3836
rect 8178 3780 8234 3836
rect 8234 3780 8238 3836
rect 8174 3776 8238 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 15948 3836 16012 3840
rect 15948 3780 15952 3836
rect 15952 3780 16008 3836
rect 16008 3780 16012 3836
rect 15948 3776 16012 3780
rect 16028 3836 16092 3840
rect 16028 3780 16032 3836
rect 16032 3780 16088 3836
rect 16088 3780 16092 3836
rect 16028 3776 16092 3780
rect 16108 3836 16172 3840
rect 16108 3780 16112 3836
rect 16112 3780 16168 3836
rect 16168 3780 16172 3836
rect 16108 3776 16172 3780
rect 16188 3836 16252 3840
rect 16188 3780 16192 3836
rect 16192 3780 16248 3836
rect 16248 3780 16252 3836
rect 16188 3776 16252 3780
rect 23722 3836 23786 3840
rect 23722 3780 23726 3836
rect 23726 3780 23782 3836
rect 23782 3780 23786 3836
rect 23722 3776 23786 3780
rect 23802 3836 23866 3840
rect 23802 3780 23806 3836
rect 23806 3780 23862 3836
rect 23862 3780 23866 3836
rect 23802 3776 23866 3780
rect 23882 3836 23946 3840
rect 23882 3780 23886 3836
rect 23886 3780 23942 3836
rect 23942 3780 23946 3836
rect 23882 3776 23946 3780
rect 23962 3836 24026 3840
rect 23962 3780 23966 3836
rect 23966 3780 24022 3836
rect 24022 3780 24026 3836
rect 23962 3776 24026 3780
rect 31496 3836 31560 3840
rect 31496 3780 31500 3836
rect 31500 3780 31556 3836
rect 31556 3780 31560 3836
rect 31496 3776 31560 3780
rect 31576 3836 31640 3840
rect 31576 3780 31580 3836
rect 31580 3780 31636 3836
rect 31636 3780 31640 3836
rect 31576 3776 31640 3780
rect 31656 3836 31720 3840
rect 31656 3780 31660 3836
rect 31660 3780 31716 3836
rect 31716 3780 31720 3836
rect 31656 3776 31720 3780
rect 31736 3836 31800 3840
rect 31736 3780 31740 3836
rect 31740 3780 31796 3836
rect 31796 3780 31800 3836
rect 31736 3776 31800 3780
rect 4287 3292 4351 3296
rect 4287 3236 4291 3292
rect 4291 3236 4347 3292
rect 4347 3236 4351 3292
rect 4287 3232 4351 3236
rect 4367 3292 4431 3296
rect 4367 3236 4371 3292
rect 4371 3236 4427 3292
rect 4427 3236 4431 3292
rect 4367 3232 4431 3236
rect 4447 3292 4511 3296
rect 4447 3236 4451 3292
rect 4451 3236 4507 3292
rect 4507 3236 4511 3292
rect 4447 3232 4511 3236
rect 4527 3292 4591 3296
rect 4527 3236 4531 3292
rect 4531 3236 4587 3292
rect 4587 3236 4591 3292
rect 4527 3232 4591 3236
rect 12061 3292 12125 3296
rect 12061 3236 12065 3292
rect 12065 3236 12121 3292
rect 12121 3236 12125 3292
rect 12061 3232 12125 3236
rect 12141 3292 12205 3296
rect 12141 3236 12145 3292
rect 12145 3236 12201 3292
rect 12201 3236 12205 3292
rect 12141 3232 12205 3236
rect 12221 3292 12285 3296
rect 12221 3236 12225 3292
rect 12225 3236 12281 3292
rect 12281 3236 12285 3292
rect 12221 3232 12285 3236
rect 12301 3292 12365 3296
rect 12301 3236 12305 3292
rect 12305 3236 12361 3292
rect 12361 3236 12365 3292
rect 12301 3232 12365 3236
rect 19835 3292 19899 3296
rect 19835 3236 19839 3292
rect 19839 3236 19895 3292
rect 19895 3236 19899 3292
rect 19835 3232 19899 3236
rect 19915 3292 19979 3296
rect 19915 3236 19919 3292
rect 19919 3236 19975 3292
rect 19975 3236 19979 3292
rect 19915 3232 19979 3236
rect 19995 3292 20059 3296
rect 19995 3236 19999 3292
rect 19999 3236 20055 3292
rect 20055 3236 20059 3292
rect 19995 3232 20059 3236
rect 20075 3292 20139 3296
rect 20075 3236 20079 3292
rect 20079 3236 20135 3292
rect 20135 3236 20139 3292
rect 20075 3232 20139 3236
rect 27609 3292 27673 3296
rect 27609 3236 27613 3292
rect 27613 3236 27669 3292
rect 27669 3236 27673 3292
rect 27609 3232 27673 3236
rect 27689 3292 27753 3296
rect 27689 3236 27693 3292
rect 27693 3236 27749 3292
rect 27749 3236 27753 3292
rect 27689 3232 27753 3236
rect 27769 3292 27833 3296
rect 27769 3236 27773 3292
rect 27773 3236 27829 3292
rect 27829 3236 27833 3292
rect 27769 3232 27833 3236
rect 27849 3292 27913 3296
rect 27849 3236 27853 3292
rect 27853 3236 27909 3292
rect 27909 3236 27913 3292
rect 27849 3232 27913 3236
rect 8174 2748 8238 2752
rect 8174 2692 8178 2748
rect 8178 2692 8234 2748
rect 8234 2692 8238 2748
rect 8174 2688 8238 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 15948 2748 16012 2752
rect 15948 2692 15952 2748
rect 15952 2692 16008 2748
rect 16008 2692 16012 2748
rect 15948 2688 16012 2692
rect 16028 2748 16092 2752
rect 16028 2692 16032 2748
rect 16032 2692 16088 2748
rect 16088 2692 16092 2748
rect 16028 2688 16092 2692
rect 16108 2748 16172 2752
rect 16108 2692 16112 2748
rect 16112 2692 16168 2748
rect 16168 2692 16172 2748
rect 16108 2688 16172 2692
rect 16188 2748 16252 2752
rect 16188 2692 16192 2748
rect 16192 2692 16248 2748
rect 16248 2692 16252 2748
rect 16188 2688 16252 2692
rect 23722 2748 23786 2752
rect 23722 2692 23726 2748
rect 23726 2692 23782 2748
rect 23782 2692 23786 2748
rect 23722 2688 23786 2692
rect 23802 2748 23866 2752
rect 23802 2692 23806 2748
rect 23806 2692 23862 2748
rect 23862 2692 23866 2748
rect 23802 2688 23866 2692
rect 23882 2748 23946 2752
rect 23882 2692 23886 2748
rect 23886 2692 23942 2748
rect 23942 2692 23946 2748
rect 23882 2688 23946 2692
rect 23962 2748 24026 2752
rect 23962 2692 23966 2748
rect 23966 2692 24022 2748
rect 24022 2692 24026 2748
rect 23962 2688 24026 2692
rect 31496 2748 31560 2752
rect 31496 2692 31500 2748
rect 31500 2692 31556 2748
rect 31556 2692 31560 2748
rect 31496 2688 31560 2692
rect 31576 2748 31640 2752
rect 31576 2692 31580 2748
rect 31580 2692 31636 2748
rect 31636 2692 31640 2748
rect 31576 2688 31640 2692
rect 31656 2748 31720 2752
rect 31656 2692 31660 2748
rect 31660 2692 31716 2748
rect 31716 2692 31720 2748
rect 31656 2688 31720 2692
rect 31736 2748 31800 2752
rect 31736 2692 31740 2748
rect 31740 2692 31796 2748
rect 31796 2692 31800 2748
rect 31736 2688 31800 2692
rect 4287 2204 4351 2208
rect 4287 2148 4291 2204
rect 4291 2148 4347 2204
rect 4347 2148 4351 2204
rect 4287 2144 4351 2148
rect 4367 2204 4431 2208
rect 4367 2148 4371 2204
rect 4371 2148 4427 2204
rect 4427 2148 4431 2204
rect 4367 2144 4431 2148
rect 4447 2204 4511 2208
rect 4447 2148 4451 2204
rect 4451 2148 4507 2204
rect 4507 2148 4511 2204
rect 4447 2144 4511 2148
rect 4527 2204 4591 2208
rect 4527 2148 4531 2204
rect 4531 2148 4587 2204
rect 4587 2148 4591 2204
rect 4527 2144 4591 2148
rect 12061 2204 12125 2208
rect 12061 2148 12065 2204
rect 12065 2148 12121 2204
rect 12121 2148 12125 2204
rect 12061 2144 12125 2148
rect 12141 2204 12205 2208
rect 12141 2148 12145 2204
rect 12145 2148 12201 2204
rect 12201 2148 12205 2204
rect 12141 2144 12205 2148
rect 12221 2204 12285 2208
rect 12221 2148 12225 2204
rect 12225 2148 12281 2204
rect 12281 2148 12285 2204
rect 12221 2144 12285 2148
rect 12301 2204 12365 2208
rect 12301 2148 12305 2204
rect 12305 2148 12361 2204
rect 12361 2148 12365 2204
rect 12301 2144 12365 2148
rect 19835 2204 19899 2208
rect 19835 2148 19839 2204
rect 19839 2148 19895 2204
rect 19895 2148 19899 2204
rect 19835 2144 19899 2148
rect 19915 2204 19979 2208
rect 19915 2148 19919 2204
rect 19919 2148 19975 2204
rect 19975 2148 19979 2204
rect 19915 2144 19979 2148
rect 19995 2204 20059 2208
rect 19995 2148 19999 2204
rect 19999 2148 20055 2204
rect 20055 2148 20059 2204
rect 19995 2144 20059 2148
rect 20075 2204 20139 2208
rect 20075 2148 20079 2204
rect 20079 2148 20135 2204
rect 20135 2148 20139 2204
rect 20075 2144 20139 2148
rect 27609 2204 27673 2208
rect 27609 2148 27613 2204
rect 27613 2148 27669 2204
rect 27669 2148 27673 2204
rect 27609 2144 27673 2148
rect 27689 2204 27753 2208
rect 27689 2148 27693 2204
rect 27693 2148 27749 2204
rect 27749 2148 27753 2204
rect 27689 2144 27753 2148
rect 27769 2204 27833 2208
rect 27769 2148 27773 2204
rect 27773 2148 27829 2204
rect 27829 2148 27833 2204
rect 27769 2144 27833 2148
rect 27849 2204 27913 2208
rect 27849 2148 27853 2204
rect 27853 2148 27909 2204
rect 27909 2148 27913 2204
rect 27849 2144 27913 2148
rect 8174 1660 8238 1664
rect 8174 1604 8178 1660
rect 8178 1604 8234 1660
rect 8234 1604 8238 1660
rect 8174 1600 8238 1604
rect 8254 1660 8318 1664
rect 8254 1604 8258 1660
rect 8258 1604 8314 1660
rect 8314 1604 8318 1660
rect 8254 1600 8318 1604
rect 8334 1660 8398 1664
rect 8334 1604 8338 1660
rect 8338 1604 8394 1660
rect 8394 1604 8398 1660
rect 8334 1600 8398 1604
rect 8414 1660 8478 1664
rect 8414 1604 8418 1660
rect 8418 1604 8474 1660
rect 8474 1604 8478 1660
rect 8414 1600 8478 1604
rect 15948 1660 16012 1664
rect 15948 1604 15952 1660
rect 15952 1604 16008 1660
rect 16008 1604 16012 1660
rect 15948 1600 16012 1604
rect 16028 1660 16092 1664
rect 16028 1604 16032 1660
rect 16032 1604 16088 1660
rect 16088 1604 16092 1660
rect 16028 1600 16092 1604
rect 16108 1660 16172 1664
rect 16108 1604 16112 1660
rect 16112 1604 16168 1660
rect 16168 1604 16172 1660
rect 16108 1600 16172 1604
rect 16188 1660 16252 1664
rect 16188 1604 16192 1660
rect 16192 1604 16248 1660
rect 16248 1604 16252 1660
rect 16188 1600 16252 1604
rect 23722 1660 23786 1664
rect 23722 1604 23726 1660
rect 23726 1604 23782 1660
rect 23782 1604 23786 1660
rect 23722 1600 23786 1604
rect 23802 1660 23866 1664
rect 23802 1604 23806 1660
rect 23806 1604 23862 1660
rect 23862 1604 23866 1660
rect 23802 1600 23866 1604
rect 23882 1660 23946 1664
rect 23882 1604 23886 1660
rect 23886 1604 23942 1660
rect 23942 1604 23946 1660
rect 23882 1600 23946 1604
rect 23962 1660 24026 1664
rect 23962 1604 23966 1660
rect 23966 1604 24022 1660
rect 24022 1604 24026 1660
rect 23962 1600 24026 1604
rect 31496 1660 31560 1664
rect 31496 1604 31500 1660
rect 31500 1604 31556 1660
rect 31556 1604 31560 1660
rect 31496 1600 31560 1604
rect 31576 1660 31640 1664
rect 31576 1604 31580 1660
rect 31580 1604 31636 1660
rect 31636 1604 31640 1660
rect 31576 1600 31640 1604
rect 31656 1660 31720 1664
rect 31656 1604 31660 1660
rect 31660 1604 31716 1660
rect 31716 1604 31720 1660
rect 31656 1600 31720 1604
rect 31736 1660 31800 1664
rect 31736 1604 31740 1660
rect 31740 1604 31796 1660
rect 31796 1604 31800 1660
rect 31736 1600 31800 1604
rect 4287 1116 4351 1120
rect 4287 1060 4291 1116
rect 4291 1060 4347 1116
rect 4347 1060 4351 1116
rect 4287 1056 4351 1060
rect 4367 1116 4431 1120
rect 4367 1060 4371 1116
rect 4371 1060 4427 1116
rect 4427 1060 4431 1116
rect 4367 1056 4431 1060
rect 4447 1116 4511 1120
rect 4447 1060 4451 1116
rect 4451 1060 4507 1116
rect 4507 1060 4511 1116
rect 4447 1056 4511 1060
rect 4527 1116 4591 1120
rect 4527 1060 4531 1116
rect 4531 1060 4587 1116
rect 4587 1060 4591 1116
rect 4527 1056 4591 1060
rect 12061 1116 12125 1120
rect 12061 1060 12065 1116
rect 12065 1060 12121 1116
rect 12121 1060 12125 1116
rect 12061 1056 12125 1060
rect 12141 1116 12205 1120
rect 12141 1060 12145 1116
rect 12145 1060 12201 1116
rect 12201 1060 12205 1116
rect 12141 1056 12205 1060
rect 12221 1116 12285 1120
rect 12221 1060 12225 1116
rect 12225 1060 12281 1116
rect 12281 1060 12285 1116
rect 12221 1056 12285 1060
rect 12301 1116 12365 1120
rect 12301 1060 12305 1116
rect 12305 1060 12361 1116
rect 12361 1060 12365 1116
rect 12301 1056 12365 1060
rect 19835 1116 19899 1120
rect 19835 1060 19839 1116
rect 19839 1060 19895 1116
rect 19895 1060 19899 1116
rect 19835 1056 19899 1060
rect 19915 1116 19979 1120
rect 19915 1060 19919 1116
rect 19919 1060 19975 1116
rect 19975 1060 19979 1116
rect 19915 1056 19979 1060
rect 19995 1116 20059 1120
rect 19995 1060 19999 1116
rect 19999 1060 20055 1116
rect 20055 1060 20059 1116
rect 19995 1056 20059 1060
rect 20075 1116 20139 1120
rect 20075 1060 20079 1116
rect 20079 1060 20135 1116
rect 20135 1060 20139 1116
rect 20075 1056 20139 1060
rect 27609 1116 27673 1120
rect 27609 1060 27613 1116
rect 27613 1060 27669 1116
rect 27669 1060 27673 1116
rect 27609 1056 27673 1060
rect 27689 1116 27753 1120
rect 27689 1060 27693 1116
rect 27693 1060 27749 1116
rect 27749 1060 27753 1116
rect 27689 1056 27753 1060
rect 27769 1116 27833 1120
rect 27769 1060 27773 1116
rect 27773 1060 27829 1116
rect 27829 1060 27833 1116
rect 27769 1056 27833 1060
rect 27849 1116 27913 1120
rect 27849 1060 27853 1116
rect 27853 1060 27909 1116
rect 27909 1060 27913 1116
rect 27849 1056 27913 1060
rect 8174 572 8238 576
rect 8174 516 8178 572
rect 8178 516 8234 572
rect 8234 516 8238 572
rect 8174 512 8238 516
rect 8254 572 8318 576
rect 8254 516 8258 572
rect 8258 516 8314 572
rect 8314 516 8318 572
rect 8254 512 8318 516
rect 8334 572 8398 576
rect 8334 516 8338 572
rect 8338 516 8394 572
rect 8394 516 8398 572
rect 8334 512 8398 516
rect 8414 572 8478 576
rect 8414 516 8418 572
rect 8418 516 8474 572
rect 8474 516 8478 572
rect 8414 512 8478 516
rect 15948 572 16012 576
rect 15948 516 15952 572
rect 15952 516 16008 572
rect 16008 516 16012 572
rect 15948 512 16012 516
rect 16028 572 16092 576
rect 16028 516 16032 572
rect 16032 516 16088 572
rect 16088 516 16092 572
rect 16028 512 16092 516
rect 16108 572 16172 576
rect 16108 516 16112 572
rect 16112 516 16168 572
rect 16168 516 16172 572
rect 16108 512 16172 516
rect 16188 572 16252 576
rect 16188 516 16192 572
rect 16192 516 16248 572
rect 16248 516 16252 572
rect 16188 512 16252 516
rect 23722 572 23786 576
rect 23722 516 23726 572
rect 23726 516 23782 572
rect 23782 516 23786 572
rect 23722 512 23786 516
rect 23802 572 23866 576
rect 23802 516 23806 572
rect 23806 516 23862 572
rect 23862 516 23866 572
rect 23802 512 23866 516
rect 23882 572 23946 576
rect 23882 516 23886 572
rect 23886 516 23942 572
rect 23942 516 23946 572
rect 23882 512 23946 516
rect 23962 572 24026 576
rect 23962 516 23966 572
rect 23966 516 24022 572
rect 24022 516 24026 572
rect 23962 512 24026 516
rect 31496 572 31560 576
rect 31496 516 31500 572
rect 31500 516 31556 572
rect 31556 516 31560 572
rect 31496 512 31560 516
rect 31576 572 31640 576
rect 31576 516 31580 572
rect 31580 516 31636 572
rect 31636 516 31640 572
rect 31576 512 31640 516
rect 31656 572 31720 576
rect 31656 516 31660 572
rect 31660 516 31716 572
rect 31716 516 31720 572
rect 31656 512 31720 516
rect 31736 572 31800 576
rect 31736 516 31740 572
rect 31740 516 31796 572
rect 31796 516 31800 572
rect 31736 512 31800 516
<< metal4 >>
rect 798 21861 858 22304
rect 1534 21861 1594 22304
rect 2270 21861 2330 22304
rect 3006 21861 3066 22304
rect 3742 21861 3802 22304
rect 4478 21997 4538 22304
rect 4475 21996 4541 21997
rect 4475 21932 4476 21996
rect 4540 21932 4541 21996
rect 4475 21931 4541 21932
rect 5214 21861 5274 22304
rect 5950 21861 6010 22304
rect 6686 21861 6746 22304
rect 7422 21861 7482 22304
rect 8158 21997 8218 22304
rect 8155 21996 8221 21997
rect 8155 21932 8156 21996
rect 8220 21932 8221 21996
rect 8155 21931 8221 21932
rect 8894 21861 8954 22304
rect 9630 21861 9690 22304
rect 10366 21861 10426 22304
rect 11102 21861 11162 22304
rect 795 21860 861 21861
rect 795 21796 796 21860
rect 860 21796 861 21860
rect 795 21795 861 21796
rect 1531 21860 1597 21861
rect 1531 21796 1532 21860
rect 1596 21796 1597 21860
rect 1531 21795 1597 21796
rect 2267 21860 2333 21861
rect 2267 21796 2268 21860
rect 2332 21796 2333 21860
rect 2267 21795 2333 21796
rect 3003 21860 3069 21861
rect 3003 21796 3004 21860
rect 3068 21796 3069 21860
rect 3003 21795 3069 21796
rect 3739 21860 3805 21861
rect 3739 21796 3740 21860
rect 3804 21796 3805 21860
rect 5211 21860 5277 21861
rect 3739 21795 3805 21796
rect 4279 21792 4599 21808
rect 5211 21796 5212 21860
rect 5276 21796 5277 21860
rect 5211 21795 5277 21796
rect 5947 21860 6013 21861
rect 5947 21796 5948 21860
rect 6012 21796 6013 21860
rect 5947 21795 6013 21796
rect 6683 21860 6749 21861
rect 6683 21796 6684 21860
rect 6748 21796 6749 21860
rect 6683 21795 6749 21796
rect 7419 21860 7485 21861
rect 7419 21796 7420 21860
rect 7484 21796 7485 21860
rect 8891 21860 8957 21861
rect 7419 21795 7485 21796
rect 4279 21728 4287 21792
rect 4351 21728 4367 21792
rect 4431 21728 4447 21792
rect 4511 21728 4527 21792
rect 4591 21728 4599 21792
rect 4279 20704 4599 21728
rect 4279 20640 4287 20704
rect 4351 20640 4367 20704
rect 4431 20640 4447 20704
rect 4511 20640 4527 20704
rect 4591 20640 4599 20704
rect 4279 19616 4599 20640
rect 4279 19552 4287 19616
rect 4351 19552 4367 19616
rect 4431 19552 4447 19616
rect 4511 19552 4527 19616
rect 4591 19552 4599 19616
rect 4279 18528 4599 19552
rect 4279 18464 4287 18528
rect 4351 18464 4367 18528
rect 4431 18464 4447 18528
rect 4511 18464 4527 18528
rect 4591 18464 4599 18528
rect 4279 17440 4599 18464
rect 4279 17376 4287 17440
rect 4351 17376 4367 17440
rect 4431 17376 4447 17440
rect 4511 17376 4527 17440
rect 4591 17376 4599 17440
rect 4279 16352 4599 17376
rect 4279 16288 4287 16352
rect 4351 16288 4367 16352
rect 4431 16288 4447 16352
rect 4511 16288 4527 16352
rect 4591 16288 4599 16352
rect 4279 15264 4599 16288
rect 4279 15200 4287 15264
rect 4351 15200 4367 15264
rect 4431 15200 4447 15264
rect 4511 15200 4527 15264
rect 4591 15200 4599 15264
rect 4279 14176 4599 15200
rect 4279 14112 4287 14176
rect 4351 14112 4367 14176
rect 4431 14112 4447 14176
rect 4511 14112 4527 14176
rect 4591 14112 4599 14176
rect 4279 13088 4599 14112
rect 4279 13024 4287 13088
rect 4351 13024 4367 13088
rect 4431 13024 4447 13088
rect 4511 13024 4527 13088
rect 4591 13024 4599 13088
rect 4279 12000 4599 13024
rect 4279 11936 4287 12000
rect 4351 11936 4367 12000
rect 4431 11936 4447 12000
rect 4511 11936 4527 12000
rect 4591 11936 4599 12000
rect 4279 10912 4599 11936
rect 4279 10848 4287 10912
rect 4351 10848 4367 10912
rect 4431 10848 4447 10912
rect 4511 10848 4527 10912
rect 4591 10848 4599 10912
rect 4279 9824 4599 10848
rect 4279 9760 4287 9824
rect 4351 9760 4367 9824
rect 4431 9760 4447 9824
rect 4511 9760 4527 9824
rect 4591 9760 4599 9824
rect 4279 8736 4599 9760
rect 4279 8672 4287 8736
rect 4351 8672 4367 8736
rect 4431 8672 4447 8736
rect 4511 8672 4527 8736
rect 4591 8672 4599 8736
rect 4279 7648 4599 8672
rect 4279 7584 4287 7648
rect 4351 7584 4367 7648
rect 4431 7584 4447 7648
rect 4511 7584 4527 7648
rect 4591 7584 4599 7648
rect 4279 6560 4599 7584
rect 4279 6496 4287 6560
rect 4351 6496 4367 6560
rect 4431 6496 4447 6560
rect 4511 6496 4527 6560
rect 4591 6496 4599 6560
rect 4279 5472 4599 6496
rect 4279 5408 4287 5472
rect 4351 5408 4367 5472
rect 4431 5408 4447 5472
rect 4511 5408 4527 5472
rect 4591 5408 4599 5472
rect 4279 4384 4599 5408
rect 4279 4320 4287 4384
rect 4351 4320 4367 4384
rect 4431 4320 4447 4384
rect 4511 4320 4527 4384
rect 4591 4320 4599 4384
rect 4279 3296 4599 4320
rect 4279 3232 4287 3296
rect 4351 3232 4367 3296
rect 4431 3232 4447 3296
rect 4511 3232 4527 3296
rect 4591 3232 4599 3296
rect 4279 2208 4599 3232
rect 4279 2144 4287 2208
rect 4351 2144 4367 2208
rect 4431 2144 4447 2208
rect 4511 2144 4527 2208
rect 4591 2144 4599 2208
rect 4279 1120 4599 2144
rect 4279 1056 4287 1120
rect 4351 1056 4367 1120
rect 4431 1056 4447 1120
rect 4511 1056 4527 1120
rect 4591 1056 4599 1120
rect 4279 496 4599 1056
rect 8166 21248 8486 21808
rect 8891 21796 8892 21860
rect 8956 21796 8957 21860
rect 8891 21795 8957 21796
rect 9627 21860 9693 21861
rect 9627 21796 9628 21860
rect 9692 21796 9693 21860
rect 9627 21795 9693 21796
rect 10363 21860 10429 21861
rect 10363 21796 10364 21860
rect 10428 21796 10429 21860
rect 10363 21795 10429 21796
rect 11099 21860 11165 21861
rect 11099 21796 11100 21860
rect 11164 21796 11165 21860
rect 11099 21795 11165 21796
rect 11838 21589 11898 22304
rect 12053 21792 12373 21808
rect 12053 21728 12061 21792
rect 12125 21728 12141 21792
rect 12205 21728 12221 21792
rect 12285 21728 12301 21792
rect 12365 21728 12373 21792
rect 11835 21588 11901 21589
rect 11835 21524 11836 21588
rect 11900 21524 11901 21588
rect 11835 21523 11901 21524
rect 8166 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8486 21248
rect 8166 20160 8486 21184
rect 8166 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8486 20160
rect 8166 19072 8486 20096
rect 8166 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8486 19072
rect 8166 17984 8486 19008
rect 8166 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8486 17984
rect 8166 16896 8486 17920
rect 8166 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8486 16896
rect 8166 15808 8486 16832
rect 8166 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8486 15808
rect 8166 14720 8486 15744
rect 8166 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8486 14720
rect 8166 13632 8486 14656
rect 8166 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8486 13632
rect 8166 12544 8486 13568
rect 8166 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8486 12544
rect 8166 11456 8486 12480
rect 8166 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8486 11456
rect 8166 10368 8486 11392
rect 8166 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8486 10368
rect 8166 9280 8486 10304
rect 8166 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8486 9280
rect 8166 8192 8486 9216
rect 8166 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8486 8192
rect 8166 7104 8486 8128
rect 8166 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8486 7104
rect 8166 6016 8486 7040
rect 8166 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8486 6016
rect 8166 4928 8486 5952
rect 8166 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8486 4928
rect 8166 3840 8486 4864
rect 8166 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8486 3840
rect 8166 2752 8486 3776
rect 8166 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8486 2752
rect 8166 1664 8486 2688
rect 8166 1600 8174 1664
rect 8238 1600 8254 1664
rect 8318 1600 8334 1664
rect 8398 1600 8414 1664
rect 8478 1600 8486 1664
rect 8166 576 8486 1600
rect 8166 512 8174 576
rect 8238 512 8254 576
rect 8318 512 8334 576
rect 8398 512 8414 576
rect 8478 512 8486 576
rect 8166 496 8486 512
rect 12053 20704 12373 21728
rect 12574 21450 12634 22304
rect 13310 21589 13370 22304
rect 13307 21588 13373 21589
rect 13307 21524 13308 21588
rect 13372 21524 13373 21588
rect 13307 21523 13373 21524
rect 12574 21390 13002 21450
rect 12053 20640 12061 20704
rect 12125 20640 12141 20704
rect 12205 20640 12221 20704
rect 12285 20640 12301 20704
rect 12365 20640 12373 20704
rect 12053 19616 12373 20640
rect 12942 20501 13002 21390
rect 14046 20773 14106 22304
rect 14043 20772 14109 20773
rect 14043 20708 14044 20772
rect 14108 20708 14109 20772
rect 14043 20707 14109 20708
rect 12939 20500 13005 20501
rect 12939 20436 12940 20500
rect 13004 20436 13005 20500
rect 12939 20435 13005 20436
rect 12053 19552 12061 19616
rect 12125 19552 12141 19616
rect 12205 19552 12221 19616
rect 12285 19552 12301 19616
rect 12365 19552 12373 19616
rect 12053 18528 12373 19552
rect 12053 18464 12061 18528
rect 12125 18464 12141 18528
rect 12205 18464 12221 18528
rect 12285 18464 12301 18528
rect 12365 18464 12373 18528
rect 12053 17440 12373 18464
rect 14782 17917 14842 22304
rect 15518 19141 15578 22304
rect 16254 22130 16314 22304
rect 16254 22070 16498 22130
rect 15940 21248 16260 21808
rect 15940 21184 15948 21248
rect 16012 21184 16028 21248
rect 16092 21184 16108 21248
rect 16172 21184 16188 21248
rect 16252 21184 16260 21248
rect 15940 20160 16260 21184
rect 15940 20096 15948 20160
rect 16012 20096 16028 20160
rect 16092 20096 16108 20160
rect 16172 20096 16188 20160
rect 16252 20096 16260 20160
rect 15515 19140 15581 19141
rect 15515 19076 15516 19140
rect 15580 19076 15581 19140
rect 15515 19075 15581 19076
rect 15940 19072 16260 20096
rect 15940 19008 15948 19072
rect 16012 19008 16028 19072
rect 16092 19008 16108 19072
rect 16172 19008 16188 19072
rect 16252 19008 16260 19072
rect 15940 17984 16260 19008
rect 15940 17920 15948 17984
rect 16012 17920 16028 17984
rect 16092 17920 16108 17984
rect 16172 17920 16188 17984
rect 16252 17920 16260 17984
rect 14779 17916 14845 17917
rect 14779 17852 14780 17916
rect 14844 17852 14845 17916
rect 14779 17851 14845 17852
rect 12053 17376 12061 17440
rect 12125 17376 12141 17440
rect 12205 17376 12221 17440
rect 12285 17376 12301 17440
rect 12365 17376 12373 17440
rect 12053 16352 12373 17376
rect 12053 16288 12061 16352
rect 12125 16288 12141 16352
rect 12205 16288 12221 16352
rect 12285 16288 12301 16352
rect 12365 16288 12373 16352
rect 12053 15264 12373 16288
rect 12053 15200 12061 15264
rect 12125 15200 12141 15264
rect 12205 15200 12221 15264
rect 12285 15200 12301 15264
rect 12365 15200 12373 15264
rect 12053 14176 12373 15200
rect 12053 14112 12061 14176
rect 12125 14112 12141 14176
rect 12205 14112 12221 14176
rect 12285 14112 12301 14176
rect 12365 14112 12373 14176
rect 12053 13088 12373 14112
rect 12053 13024 12061 13088
rect 12125 13024 12141 13088
rect 12205 13024 12221 13088
rect 12285 13024 12301 13088
rect 12365 13024 12373 13088
rect 12053 12000 12373 13024
rect 12053 11936 12061 12000
rect 12125 11936 12141 12000
rect 12205 11936 12221 12000
rect 12285 11936 12301 12000
rect 12365 11936 12373 12000
rect 12053 10912 12373 11936
rect 12053 10848 12061 10912
rect 12125 10848 12141 10912
rect 12205 10848 12221 10912
rect 12285 10848 12301 10912
rect 12365 10848 12373 10912
rect 12053 9824 12373 10848
rect 12053 9760 12061 9824
rect 12125 9760 12141 9824
rect 12205 9760 12221 9824
rect 12285 9760 12301 9824
rect 12365 9760 12373 9824
rect 12053 8736 12373 9760
rect 12053 8672 12061 8736
rect 12125 8672 12141 8736
rect 12205 8672 12221 8736
rect 12285 8672 12301 8736
rect 12365 8672 12373 8736
rect 12053 7648 12373 8672
rect 12053 7584 12061 7648
rect 12125 7584 12141 7648
rect 12205 7584 12221 7648
rect 12285 7584 12301 7648
rect 12365 7584 12373 7648
rect 12053 6560 12373 7584
rect 12053 6496 12061 6560
rect 12125 6496 12141 6560
rect 12205 6496 12221 6560
rect 12285 6496 12301 6560
rect 12365 6496 12373 6560
rect 12053 5472 12373 6496
rect 12053 5408 12061 5472
rect 12125 5408 12141 5472
rect 12205 5408 12221 5472
rect 12285 5408 12301 5472
rect 12365 5408 12373 5472
rect 12053 4384 12373 5408
rect 12053 4320 12061 4384
rect 12125 4320 12141 4384
rect 12205 4320 12221 4384
rect 12285 4320 12301 4384
rect 12365 4320 12373 4384
rect 12053 3296 12373 4320
rect 12053 3232 12061 3296
rect 12125 3232 12141 3296
rect 12205 3232 12221 3296
rect 12285 3232 12301 3296
rect 12365 3232 12373 3296
rect 12053 2208 12373 3232
rect 12053 2144 12061 2208
rect 12125 2144 12141 2208
rect 12205 2144 12221 2208
rect 12285 2144 12301 2208
rect 12365 2144 12373 2208
rect 12053 1120 12373 2144
rect 12053 1056 12061 1120
rect 12125 1056 12141 1120
rect 12205 1056 12221 1120
rect 12285 1056 12301 1120
rect 12365 1056 12373 1120
rect 12053 496 12373 1056
rect 15940 16896 16260 17920
rect 16438 17917 16498 22070
rect 16990 21317 17050 22304
rect 16987 21316 17053 21317
rect 16987 21252 16988 21316
rect 17052 21252 17053 21316
rect 16987 21251 17053 21252
rect 16435 17916 16501 17917
rect 16435 17852 16436 17916
rect 16500 17852 16501 17916
rect 16435 17851 16501 17852
rect 15940 16832 15948 16896
rect 16012 16832 16028 16896
rect 16092 16832 16108 16896
rect 16172 16832 16188 16896
rect 16252 16832 16260 16896
rect 15940 15808 16260 16832
rect 17726 16557 17786 22304
rect 18462 22104 18522 22304
rect 19198 22104 19258 22304
rect 19934 22104 19994 22304
rect 20670 22104 20730 22304
rect 21406 22104 21466 22304
rect 22142 22104 22202 22304
rect 22878 22104 22938 22304
rect 23614 22104 23674 22304
rect 24350 22104 24410 22304
rect 25086 22104 25146 22304
rect 25822 21861 25882 22304
rect 26558 21861 26618 22304
rect 27294 22130 27354 22304
rect 27294 22070 27538 22130
rect 27478 21997 27538 22070
rect 27475 21996 27541 21997
rect 27475 21932 27476 21996
rect 27540 21932 27541 21996
rect 27475 21931 27541 21932
rect 28030 21861 28090 22304
rect 25819 21860 25885 21861
rect 19827 21792 20147 21808
rect 19827 21728 19835 21792
rect 19899 21728 19915 21792
rect 19979 21728 19995 21792
rect 20059 21728 20075 21792
rect 20139 21728 20147 21792
rect 19827 20704 20147 21728
rect 19827 20640 19835 20704
rect 19899 20640 19915 20704
rect 19979 20640 19995 20704
rect 20059 20640 20075 20704
rect 20139 20640 20147 20704
rect 19827 19616 20147 20640
rect 19827 19552 19835 19616
rect 19899 19552 19915 19616
rect 19979 19552 19995 19616
rect 20059 19552 20075 19616
rect 20139 19552 20147 19616
rect 19827 18528 20147 19552
rect 19827 18464 19835 18528
rect 19899 18464 19915 18528
rect 19979 18464 19995 18528
rect 20059 18464 20075 18528
rect 20139 18464 20147 18528
rect 19827 17440 20147 18464
rect 19827 17376 19835 17440
rect 19899 17376 19915 17440
rect 19979 17376 19995 17440
rect 20059 17376 20075 17440
rect 20139 17376 20147 17440
rect 17723 16556 17789 16557
rect 17723 16492 17724 16556
rect 17788 16492 17789 16556
rect 17723 16491 17789 16492
rect 15940 15744 15948 15808
rect 16012 15744 16028 15808
rect 16092 15744 16108 15808
rect 16172 15744 16188 15808
rect 16252 15744 16260 15808
rect 15940 14720 16260 15744
rect 15940 14656 15948 14720
rect 16012 14656 16028 14720
rect 16092 14656 16108 14720
rect 16172 14656 16188 14720
rect 16252 14656 16260 14720
rect 15940 13632 16260 14656
rect 15940 13568 15948 13632
rect 16012 13568 16028 13632
rect 16092 13568 16108 13632
rect 16172 13568 16188 13632
rect 16252 13568 16260 13632
rect 15940 12544 16260 13568
rect 15940 12480 15948 12544
rect 16012 12480 16028 12544
rect 16092 12480 16108 12544
rect 16172 12480 16188 12544
rect 16252 12480 16260 12544
rect 15940 11456 16260 12480
rect 15940 11392 15948 11456
rect 16012 11392 16028 11456
rect 16092 11392 16108 11456
rect 16172 11392 16188 11456
rect 16252 11392 16260 11456
rect 15940 10368 16260 11392
rect 15940 10304 15948 10368
rect 16012 10304 16028 10368
rect 16092 10304 16108 10368
rect 16172 10304 16188 10368
rect 16252 10304 16260 10368
rect 15940 9280 16260 10304
rect 15940 9216 15948 9280
rect 16012 9216 16028 9280
rect 16092 9216 16108 9280
rect 16172 9216 16188 9280
rect 16252 9216 16260 9280
rect 15940 8192 16260 9216
rect 15940 8128 15948 8192
rect 16012 8128 16028 8192
rect 16092 8128 16108 8192
rect 16172 8128 16188 8192
rect 16252 8128 16260 8192
rect 15940 7104 16260 8128
rect 15940 7040 15948 7104
rect 16012 7040 16028 7104
rect 16092 7040 16108 7104
rect 16172 7040 16188 7104
rect 16252 7040 16260 7104
rect 15940 6016 16260 7040
rect 15940 5952 15948 6016
rect 16012 5952 16028 6016
rect 16092 5952 16108 6016
rect 16172 5952 16188 6016
rect 16252 5952 16260 6016
rect 15940 4928 16260 5952
rect 15940 4864 15948 4928
rect 16012 4864 16028 4928
rect 16092 4864 16108 4928
rect 16172 4864 16188 4928
rect 16252 4864 16260 4928
rect 15940 3840 16260 4864
rect 15940 3776 15948 3840
rect 16012 3776 16028 3840
rect 16092 3776 16108 3840
rect 16172 3776 16188 3840
rect 16252 3776 16260 3840
rect 15940 2752 16260 3776
rect 15940 2688 15948 2752
rect 16012 2688 16028 2752
rect 16092 2688 16108 2752
rect 16172 2688 16188 2752
rect 16252 2688 16260 2752
rect 15940 1664 16260 2688
rect 15940 1600 15948 1664
rect 16012 1600 16028 1664
rect 16092 1600 16108 1664
rect 16172 1600 16188 1664
rect 16252 1600 16260 1664
rect 15940 576 16260 1600
rect 15940 512 15948 576
rect 16012 512 16028 576
rect 16092 512 16108 576
rect 16172 512 16188 576
rect 16252 512 16260 576
rect 15940 496 16260 512
rect 19827 16352 20147 17376
rect 19827 16288 19835 16352
rect 19899 16288 19915 16352
rect 19979 16288 19995 16352
rect 20059 16288 20075 16352
rect 20139 16288 20147 16352
rect 19827 15264 20147 16288
rect 19827 15200 19835 15264
rect 19899 15200 19915 15264
rect 19979 15200 19995 15264
rect 20059 15200 20075 15264
rect 20139 15200 20147 15264
rect 19827 14176 20147 15200
rect 19827 14112 19835 14176
rect 19899 14112 19915 14176
rect 19979 14112 19995 14176
rect 20059 14112 20075 14176
rect 20139 14112 20147 14176
rect 19827 13088 20147 14112
rect 19827 13024 19835 13088
rect 19899 13024 19915 13088
rect 19979 13024 19995 13088
rect 20059 13024 20075 13088
rect 20139 13024 20147 13088
rect 19827 12000 20147 13024
rect 19827 11936 19835 12000
rect 19899 11936 19915 12000
rect 19979 11936 19995 12000
rect 20059 11936 20075 12000
rect 20139 11936 20147 12000
rect 19827 10912 20147 11936
rect 19827 10848 19835 10912
rect 19899 10848 19915 10912
rect 19979 10848 19995 10912
rect 20059 10848 20075 10912
rect 20139 10848 20147 10912
rect 19827 9824 20147 10848
rect 19827 9760 19835 9824
rect 19899 9760 19915 9824
rect 19979 9760 19995 9824
rect 20059 9760 20075 9824
rect 20139 9760 20147 9824
rect 19827 8736 20147 9760
rect 19827 8672 19835 8736
rect 19899 8672 19915 8736
rect 19979 8672 19995 8736
rect 20059 8672 20075 8736
rect 20139 8672 20147 8736
rect 19827 7648 20147 8672
rect 19827 7584 19835 7648
rect 19899 7584 19915 7648
rect 19979 7584 19995 7648
rect 20059 7584 20075 7648
rect 20139 7584 20147 7648
rect 19827 6560 20147 7584
rect 19827 6496 19835 6560
rect 19899 6496 19915 6560
rect 19979 6496 19995 6560
rect 20059 6496 20075 6560
rect 20139 6496 20147 6560
rect 19827 5472 20147 6496
rect 19827 5408 19835 5472
rect 19899 5408 19915 5472
rect 19979 5408 19995 5472
rect 20059 5408 20075 5472
rect 20139 5408 20147 5472
rect 19827 4384 20147 5408
rect 19827 4320 19835 4384
rect 19899 4320 19915 4384
rect 19979 4320 19995 4384
rect 20059 4320 20075 4384
rect 20139 4320 20147 4384
rect 19827 3296 20147 4320
rect 19827 3232 19835 3296
rect 19899 3232 19915 3296
rect 19979 3232 19995 3296
rect 20059 3232 20075 3296
rect 20139 3232 20147 3296
rect 19827 2208 20147 3232
rect 19827 2144 19835 2208
rect 19899 2144 19915 2208
rect 19979 2144 19995 2208
rect 20059 2144 20075 2208
rect 20139 2144 20147 2208
rect 19827 1120 20147 2144
rect 19827 1056 19835 1120
rect 19899 1056 19915 1120
rect 19979 1056 19995 1120
rect 20059 1056 20075 1120
rect 20139 1056 20147 1120
rect 19827 496 20147 1056
rect 23714 21248 24034 21808
rect 25819 21796 25820 21860
rect 25884 21796 25885 21860
rect 25819 21795 25885 21796
rect 26555 21860 26621 21861
rect 26555 21796 26556 21860
rect 26620 21796 26621 21860
rect 28027 21860 28093 21861
rect 26555 21795 26621 21796
rect 23714 21184 23722 21248
rect 23786 21184 23802 21248
rect 23866 21184 23882 21248
rect 23946 21184 23962 21248
rect 24026 21184 24034 21248
rect 23714 20160 24034 21184
rect 23714 20096 23722 20160
rect 23786 20096 23802 20160
rect 23866 20096 23882 20160
rect 23946 20096 23962 20160
rect 24026 20096 24034 20160
rect 23714 19072 24034 20096
rect 23714 19008 23722 19072
rect 23786 19008 23802 19072
rect 23866 19008 23882 19072
rect 23946 19008 23962 19072
rect 24026 19008 24034 19072
rect 23714 17984 24034 19008
rect 23714 17920 23722 17984
rect 23786 17920 23802 17984
rect 23866 17920 23882 17984
rect 23946 17920 23962 17984
rect 24026 17920 24034 17984
rect 23714 16896 24034 17920
rect 23714 16832 23722 16896
rect 23786 16832 23802 16896
rect 23866 16832 23882 16896
rect 23946 16832 23962 16896
rect 24026 16832 24034 16896
rect 23714 15808 24034 16832
rect 23714 15744 23722 15808
rect 23786 15744 23802 15808
rect 23866 15744 23882 15808
rect 23946 15744 23962 15808
rect 24026 15744 24034 15808
rect 23714 14720 24034 15744
rect 23714 14656 23722 14720
rect 23786 14656 23802 14720
rect 23866 14656 23882 14720
rect 23946 14656 23962 14720
rect 24026 14656 24034 14720
rect 23714 13632 24034 14656
rect 23714 13568 23722 13632
rect 23786 13568 23802 13632
rect 23866 13568 23882 13632
rect 23946 13568 23962 13632
rect 24026 13568 24034 13632
rect 23714 12544 24034 13568
rect 23714 12480 23722 12544
rect 23786 12480 23802 12544
rect 23866 12480 23882 12544
rect 23946 12480 23962 12544
rect 24026 12480 24034 12544
rect 23714 11456 24034 12480
rect 23714 11392 23722 11456
rect 23786 11392 23802 11456
rect 23866 11392 23882 11456
rect 23946 11392 23962 11456
rect 24026 11392 24034 11456
rect 23714 10368 24034 11392
rect 23714 10304 23722 10368
rect 23786 10304 23802 10368
rect 23866 10304 23882 10368
rect 23946 10304 23962 10368
rect 24026 10304 24034 10368
rect 23714 9280 24034 10304
rect 23714 9216 23722 9280
rect 23786 9216 23802 9280
rect 23866 9216 23882 9280
rect 23946 9216 23962 9280
rect 24026 9216 24034 9280
rect 23714 8192 24034 9216
rect 23714 8128 23722 8192
rect 23786 8128 23802 8192
rect 23866 8128 23882 8192
rect 23946 8128 23962 8192
rect 24026 8128 24034 8192
rect 23714 7104 24034 8128
rect 23714 7040 23722 7104
rect 23786 7040 23802 7104
rect 23866 7040 23882 7104
rect 23946 7040 23962 7104
rect 24026 7040 24034 7104
rect 23714 6016 24034 7040
rect 23714 5952 23722 6016
rect 23786 5952 23802 6016
rect 23866 5952 23882 6016
rect 23946 5952 23962 6016
rect 24026 5952 24034 6016
rect 23714 4928 24034 5952
rect 23714 4864 23722 4928
rect 23786 4864 23802 4928
rect 23866 4864 23882 4928
rect 23946 4864 23962 4928
rect 24026 4864 24034 4928
rect 23714 3840 24034 4864
rect 23714 3776 23722 3840
rect 23786 3776 23802 3840
rect 23866 3776 23882 3840
rect 23946 3776 23962 3840
rect 24026 3776 24034 3840
rect 23714 2752 24034 3776
rect 23714 2688 23722 2752
rect 23786 2688 23802 2752
rect 23866 2688 23882 2752
rect 23946 2688 23962 2752
rect 24026 2688 24034 2752
rect 23714 1664 24034 2688
rect 23714 1600 23722 1664
rect 23786 1600 23802 1664
rect 23866 1600 23882 1664
rect 23946 1600 23962 1664
rect 24026 1600 24034 1664
rect 23714 576 24034 1600
rect 23714 512 23722 576
rect 23786 512 23802 576
rect 23866 512 23882 576
rect 23946 512 23962 576
rect 24026 512 24034 576
rect 23714 496 24034 512
rect 27601 21792 27921 21808
rect 28027 21796 28028 21860
rect 28092 21796 28093 21860
rect 28027 21795 28093 21796
rect 27601 21728 27609 21792
rect 27673 21728 27689 21792
rect 27753 21728 27769 21792
rect 27833 21728 27849 21792
rect 27913 21728 27921 21792
rect 27601 20704 27921 21728
rect 28766 21725 28826 22304
rect 29502 21861 29562 22304
rect 30238 22104 30298 22304
rect 30974 22104 31034 22304
rect 31710 22104 31770 22304
rect 29499 21860 29565 21861
rect 29499 21796 29500 21860
rect 29564 21796 29565 21860
rect 29499 21795 29565 21796
rect 28763 21724 28829 21725
rect 28763 21660 28764 21724
rect 28828 21660 28829 21724
rect 28763 21659 28829 21660
rect 27601 20640 27609 20704
rect 27673 20640 27689 20704
rect 27753 20640 27769 20704
rect 27833 20640 27849 20704
rect 27913 20640 27921 20704
rect 27601 19616 27921 20640
rect 27601 19552 27609 19616
rect 27673 19552 27689 19616
rect 27753 19552 27769 19616
rect 27833 19552 27849 19616
rect 27913 19552 27921 19616
rect 27601 18528 27921 19552
rect 27601 18464 27609 18528
rect 27673 18464 27689 18528
rect 27753 18464 27769 18528
rect 27833 18464 27849 18528
rect 27913 18464 27921 18528
rect 27601 17440 27921 18464
rect 27601 17376 27609 17440
rect 27673 17376 27689 17440
rect 27753 17376 27769 17440
rect 27833 17376 27849 17440
rect 27913 17376 27921 17440
rect 27601 16352 27921 17376
rect 27601 16288 27609 16352
rect 27673 16288 27689 16352
rect 27753 16288 27769 16352
rect 27833 16288 27849 16352
rect 27913 16288 27921 16352
rect 27601 15264 27921 16288
rect 27601 15200 27609 15264
rect 27673 15200 27689 15264
rect 27753 15200 27769 15264
rect 27833 15200 27849 15264
rect 27913 15200 27921 15264
rect 27601 14176 27921 15200
rect 27601 14112 27609 14176
rect 27673 14112 27689 14176
rect 27753 14112 27769 14176
rect 27833 14112 27849 14176
rect 27913 14112 27921 14176
rect 27601 13088 27921 14112
rect 27601 13024 27609 13088
rect 27673 13024 27689 13088
rect 27753 13024 27769 13088
rect 27833 13024 27849 13088
rect 27913 13024 27921 13088
rect 27601 12000 27921 13024
rect 27601 11936 27609 12000
rect 27673 11936 27689 12000
rect 27753 11936 27769 12000
rect 27833 11936 27849 12000
rect 27913 11936 27921 12000
rect 27601 10912 27921 11936
rect 27601 10848 27609 10912
rect 27673 10848 27689 10912
rect 27753 10848 27769 10912
rect 27833 10848 27849 10912
rect 27913 10848 27921 10912
rect 27601 9824 27921 10848
rect 27601 9760 27609 9824
rect 27673 9760 27689 9824
rect 27753 9760 27769 9824
rect 27833 9760 27849 9824
rect 27913 9760 27921 9824
rect 27601 8736 27921 9760
rect 27601 8672 27609 8736
rect 27673 8672 27689 8736
rect 27753 8672 27769 8736
rect 27833 8672 27849 8736
rect 27913 8672 27921 8736
rect 27601 7648 27921 8672
rect 27601 7584 27609 7648
rect 27673 7584 27689 7648
rect 27753 7584 27769 7648
rect 27833 7584 27849 7648
rect 27913 7584 27921 7648
rect 27601 6560 27921 7584
rect 27601 6496 27609 6560
rect 27673 6496 27689 6560
rect 27753 6496 27769 6560
rect 27833 6496 27849 6560
rect 27913 6496 27921 6560
rect 27601 5472 27921 6496
rect 27601 5408 27609 5472
rect 27673 5408 27689 5472
rect 27753 5408 27769 5472
rect 27833 5408 27849 5472
rect 27913 5408 27921 5472
rect 27601 4384 27921 5408
rect 27601 4320 27609 4384
rect 27673 4320 27689 4384
rect 27753 4320 27769 4384
rect 27833 4320 27849 4384
rect 27913 4320 27921 4384
rect 27601 3296 27921 4320
rect 27601 3232 27609 3296
rect 27673 3232 27689 3296
rect 27753 3232 27769 3296
rect 27833 3232 27849 3296
rect 27913 3232 27921 3296
rect 27601 2208 27921 3232
rect 27601 2144 27609 2208
rect 27673 2144 27689 2208
rect 27753 2144 27769 2208
rect 27833 2144 27849 2208
rect 27913 2144 27921 2208
rect 27601 1120 27921 2144
rect 27601 1056 27609 1120
rect 27673 1056 27689 1120
rect 27753 1056 27769 1120
rect 27833 1056 27849 1120
rect 27913 1056 27921 1120
rect 27601 496 27921 1056
rect 31488 21248 31808 21808
rect 31488 21184 31496 21248
rect 31560 21184 31576 21248
rect 31640 21184 31656 21248
rect 31720 21184 31736 21248
rect 31800 21184 31808 21248
rect 31488 20160 31808 21184
rect 31488 20096 31496 20160
rect 31560 20096 31576 20160
rect 31640 20096 31656 20160
rect 31720 20096 31736 20160
rect 31800 20096 31808 20160
rect 31488 19072 31808 20096
rect 31488 19008 31496 19072
rect 31560 19008 31576 19072
rect 31640 19008 31656 19072
rect 31720 19008 31736 19072
rect 31800 19008 31808 19072
rect 31488 17984 31808 19008
rect 31488 17920 31496 17984
rect 31560 17920 31576 17984
rect 31640 17920 31656 17984
rect 31720 17920 31736 17984
rect 31800 17920 31808 17984
rect 31488 16896 31808 17920
rect 31488 16832 31496 16896
rect 31560 16832 31576 16896
rect 31640 16832 31656 16896
rect 31720 16832 31736 16896
rect 31800 16832 31808 16896
rect 31488 15808 31808 16832
rect 31488 15744 31496 15808
rect 31560 15744 31576 15808
rect 31640 15744 31656 15808
rect 31720 15744 31736 15808
rect 31800 15744 31808 15808
rect 31488 14720 31808 15744
rect 31488 14656 31496 14720
rect 31560 14656 31576 14720
rect 31640 14656 31656 14720
rect 31720 14656 31736 14720
rect 31800 14656 31808 14720
rect 31488 13632 31808 14656
rect 31488 13568 31496 13632
rect 31560 13568 31576 13632
rect 31640 13568 31656 13632
rect 31720 13568 31736 13632
rect 31800 13568 31808 13632
rect 31488 12544 31808 13568
rect 31488 12480 31496 12544
rect 31560 12480 31576 12544
rect 31640 12480 31656 12544
rect 31720 12480 31736 12544
rect 31800 12480 31808 12544
rect 31488 11456 31808 12480
rect 31488 11392 31496 11456
rect 31560 11392 31576 11456
rect 31640 11392 31656 11456
rect 31720 11392 31736 11456
rect 31800 11392 31808 11456
rect 31488 10368 31808 11392
rect 31488 10304 31496 10368
rect 31560 10304 31576 10368
rect 31640 10304 31656 10368
rect 31720 10304 31736 10368
rect 31800 10304 31808 10368
rect 31488 9280 31808 10304
rect 31488 9216 31496 9280
rect 31560 9216 31576 9280
rect 31640 9216 31656 9280
rect 31720 9216 31736 9280
rect 31800 9216 31808 9280
rect 31488 8192 31808 9216
rect 31488 8128 31496 8192
rect 31560 8128 31576 8192
rect 31640 8128 31656 8192
rect 31720 8128 31736 8192
rect 31800 8128 31808 8192
rect 31488 7104 31808 8128
rect 31488 7040 31496 7104
rect 31560 7040 31576 7104
rect 31640 7040 31656 7104
rect 31720 7040 31736 7104
rect 31800 7040 31808 7104
rect 31488 6016 31808 7040
rect 31488 5952 31496 6016
rect 31560 5952 31576 6016
rect 31640 5952 31656 6016
rect 31720 5952 31736 6016
rect 31800 5952 31808 6016
rect 31488 4928 31808 5952
rect 31488 4864 31496 4928
rect 31560 4864 31576 4928
rect 31640 4864 31656 4928
rect 31720 4864 31736 4928
rect 31800 4864 31808 4928
rect 31488 3840 31808 4864
rect 31488 3776 31496 3840
rect 31560 3776 31576 3840
rect 31640 3776 31656 3840
rect 31720 3776 31736 3840
rect 31800 3776 31808 3840
rect 31488 2752 31808 3776
rect 31488 2688 31496 2752
rect 31560 2688 31576 2752
rect 31640 2688 31656 2752
rect 31720 2688 31736 2752
rect 31800 2688 31808 2752
rect 31488 1664 31808 2688
rect 31488 1600 31496 1664
rect 31560 1600 31576 1664
rect 31640 1600 31656 1664
rect 31720 1600 31736 1664
rect 31800 1600 31808 1664
rect 31488 576 31808 1600
rect 31488 512 31496 576
rect 31560 512 31576 576
rect 31640 512 31656 576
rect 31720 512 31736 576
rect 31800 512 31808 576
rect 31488 496 31808 512
use sky130_fd_sc_hd__clkbuf_2  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 25944 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 27232 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 25300 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _238_
timestamp 1698431365
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 25944 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15088 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 16744 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _242_
timestamp 1698431365
transform -1 0 24932 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_2  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 24104 0 1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _244_
timestamp 1698431365
transform 1 0 12880 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _245_
timestamp 1698431365
transform -1 0 27232 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _246_
timestamp 1698431365
transform -1 0 15916 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _247_
timestamp 1698431365
transform 1 0 13708 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16744 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 15548 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _250_
timestamp 1698431365
transform -1 0 17756 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _251_
timestamp 1698431365
transform -1 0 20148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 25116 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 23000 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _254_
timestamp 1698431365
transform -1 0 16652 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 24840 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _256_
timestamp 1698431365
transform -1 0 23184 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 25852 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 26312 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21252 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21436 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21712 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 17112 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 17112 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1698431365
transform -1 0 14720 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _265_
timestamp 1698431365
transform 1 0 13524 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _266_
timestamp 1698431365
transform 1 0 13708 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _267_
timestamp 1698431365
transform 1 0 15088 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _268_
timestamp 1698431365
transform -1 0 24840 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _269_
timestamp 1698431365
transform -1 0 24840 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _270_
timestamp 1698431365
transform -1 0 25760 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _271_
timestamp 1698431365
transform -1 0 24380 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _272_
timestamp 1698431365
transform -1 0 16560 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _273_
timestamp 1698431365
transform 1 0 16560 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _274_
timestamp 1698431365
transform 1 0 13064 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _275_
timestamp 1698431365
transform 1 0 14352 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _276_
timestamp 1698431365
transform 1 0 13800 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 27324 0 -1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__a311o_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 22540 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _279_
timestamp 1698431365
transform 1 0 21620 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _280_
timestamp 1698431365
transform -1 0 22724 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _281_
timestamp 1698431365
transform 1 0 22264 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_4  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 16100 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _283_
timestamp 1698431365
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _284_
timestamp 1698431365
transform -1 0 23644 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _285_
timestamp 1698431365
transform -1 0 18492 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _286_
timestamp 1698431365
transform -1 0 18308 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _287_
timestamp 1698431365
transform 1 0 13524 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _288_
timestamp 1698431365
transform 1 0 12696 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _289_
timestamp 1698431365
transform 1 0 12696 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _290_
timestamp 1698431365
transform 1 0 13432 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1698431365
transform 1 0 14352 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _292_
timestamp 1698431365
transform -1 0 15088 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _293_
timestamp 1698431365
transform 1 0 12052 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _294_
timestamp 1698431365
transform 1 0 12696 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _295_
timestamp 1698431365
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _296_
timestamp 1698431365
transform 1 0 26404 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _297_
timestamp 1698431365
transform 1 0 27324 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _298_
timestamp 1698431365
transform -1 0 28244 0 -1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__a2111o_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 26496 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 20884 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _301_
timestamp 1698431365
transform -1 0 20700 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 14812 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _303_
timestamp 1698431365
transform -1 0 13984 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _304_
timestamp 1698431365
transform -1 0 13248 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _305_
timestamp 1698431365
transform -1 0 24748 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _306_
timestamp 1698431365
transform -1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _307_
timestamp 1698431365
transform -1 0 13248 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _308_
timestamp 1698431365
transform -1 0 19596 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _309_
timestamp 1698431365
transform -1 0 19320 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _310_
timestamp 1698431365
transform 1 0 18676 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 13248 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_1  _312_
timestamp 1698431365
transform 1 0 13524 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _313_
timestamp 1698431365
transform 1 0 12788 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _314_
timestamp 1698431365
transform 1 0 13156 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _315_
timestamp 1698431365
transform 1 0 13892 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _316_
timestamp 1698431365
transform -1 0 25484 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _317_
timestamp 1698431365
transform 1 0 24104 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _318_
timestamp 1698431365
transform 1 0 23828 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 25024 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _320_
timestamp 1698431365
transform -1 0 15088 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _321_
timestamp 1698431365
transform 1 0 14076 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_1  _322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 13524 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 13892 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 13708 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 14168 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _326_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 14168 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _327_
timestamp 1698431365
transform -1 0 12052 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _328_
timestamp 1698431365
transform -1 0 13248 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _329_
timestamp 1698431365
transform -1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _330_
timestamp 1698431365
transform 1 0 8740 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _331_
timestamp 1698431365
transform -1 0 9476 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _332_
timestamp 1698431365
transform -1 0 8188 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _333_
timestamp 1698431365
transform -1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _334_
timestamp 1698431365
transform -1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _335_
timestamp 1698431365
transform -1 0 6992 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _336_
timestamp 1698431365
transform -1 0 7728 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _337_
timestamp 1698431365
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _338_
timestamp 1698431365
transform -1 0 7360 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _339_
timestamp 1698431365
transform 1 0 5244 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _340_
timestamp 1698431365
transform -1 0 6348 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _341_
timestamp 1698431365
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _342_
timestamp 1698431365
transform 1 0 2668 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 2300 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 2576 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _345_
timestamp 1698431365
transform -1 0 3128 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _346_
timestamp 1698431365
transform -1 0 1656 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _347_
timestamp 1698431365
transform 1 0 3404 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _348_
timestamp 1698431365
transform -1 0 6440 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _349_
timestamp 1698431365
transform -1 0 5428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3772 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 6440 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _352_
timestamp 1698431365
transform 1 0 828 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _353_
timestamp 1698431365
transform 1 0 2852 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _354_
timestamp 1698431365
transform 1 0 3404 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _355_
timestamp 1698431365
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _356_
timestamp 1698431365
transform -1 0 2116 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 2576 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _358_
timestamp 1698431365
transform -1 0 1288 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _359_
timestamp 1698431365
transform 1 0 1012 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _360_
timestamp 1698431365
transform 1 0 28244 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _361_
timestamp 1698431365
transform -1 0 29072 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _362_
timestamp 1698431365
transform 1 0 28428 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _363_
timestamp 1698431365
transform 1 0 29348 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _364_
timestamp 1698431365
transform 1 0 28796 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _365_
timestamp 1698431365
transform -1 0 29808 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _366_
timestamp 1698431365
transform 1 0 29072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _367_
timestamp 1698431365
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _368_
timestamp 1698431365
transform 1 0 26404 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _369_
timestamp 1698431365
transform -1 0 25208 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _370_
timestamp 1698431365
transform 1 0 24288 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _371_
timestamp 1698431365
transform -1 0 24288 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _372_
timestamp 1698431365
transform 1 0 25208 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _373_
timestamp 1698431365
transform 1 0 24564 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _374_
timestamp 1698431365
transform -1 0 25300 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1698431365
transform -1 0 25576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _376_
timestamp 1698431365
transform -1 0 23736 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _377_
timestamp 1698431365
transform 1 0 22172 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _378_
timestamp 1698431365
transform 1 0 23184 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _379_
timestamp 1698431365
transform 1 0 24472 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _380_
timestamp 1698431365
transform 1 0 23368 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _381_
timestamp 1698431365
transform 1 0 25208 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _382_
timestamp 1698431365
transform 1 0 25576 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _383_
timestamp 1698431365
transform -1 0 21712 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _384_
timestamp 1698431365
transform 1 0 21068 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _385_
timestamp 1698431365
transform -1 0 21896 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _386_
timestamp 1698431365
transform 1 0 20792 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _387_
timestamp 1698431365
transform -1 0 22172 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _388_
timestamp 1698431365
transform 1 0 19872 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _389_
timestamp 1698431365
transform -1 0 23276 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _390_
timestamp 1698431365
transform -1 0 17388 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _391_
timestamp 1698431365
transform -1 0 18308 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _392_
timestamp 1698431365
transform -1 0 17940 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _393_
timestamp 1698431365
transform 1 0 17480 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _394_
timestamp 1698431365
transform 1 0 17664 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _395_
timestamp 1698431365
transform -1 0 18400 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _396_
timestamp 1698431365
transform 1 0 18308 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _397_
timestamp 1698431365
transform 1 0 19320 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1698431365
transform -1 0 12144 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1698431365
transform -1 0 26956 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _400_
timestamp 1698431365
transform 1 0 12420 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _401_
timestamp 1698431365
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _402_
timestamp 1698431365
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _403_
timestamp 1698431365
transform 1 0 20608 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _404_
timestamp 1698431365
transform 1 0 20884 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _405_
timestamp 1698431365
transform -1 0 23184 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _406_
timestamp 1698431365
transform 1 0 21252 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _407_
timestamp 1698431365
transform -1 0 18860 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_4  _408_
timestamp 1698431365
transform 1 0 5060 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1698431365
transform 1 0 12236 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1698431365
transform 1 0 15548 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1698431365
transform -1 0 14996 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1698431365
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1698431365
transform 1 0 10396 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1698431365
transform -1 0 10764 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1698431365
transform -1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1698431365
transform 1 0 6072 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1698431365
transform -1 0 5520 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1698431365
transform -1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1698431365
transform -1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1698431365
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1698431365
transform -1 0 3312 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1698431365
transform 1 0 4324 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1698431365
transform -1 0 2760 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1698431365
transform -1 0 2484 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _425_
timestamp 1698431365
transform 1 0 28888 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1698431365
transform -1 0 28704 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1698431365
transform 1 0 29992 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1698431365
transform 1 0 30176 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1698431365
transform 1 0 30912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1698431365
transform -1 0 28612 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1698431365
transform -1 0 25760 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1698431365
transform 1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1698431365
transform -1 0 25668 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1698431365
transform -1 0 26128 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1698431365
transform -1 0 27600 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1698431365
transform 1 0 22816 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1698431365
transform 1 0 19688 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1698431365
transform -1 0 18584 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1698431365
transform -1 0 18952 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1698431365
transform -1 0 17112 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1698431365
transform -1 0 21528 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 11960 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1698431365
transform 1 0 14536 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _444_
timestamp 1698431365
transform 1 0 12696 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _445_
timestamp 1698431365
transform 1 0 13064 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1698431365
transform 1 0 10488 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1698431365
transform 1 0 10948 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1698431365
transform 1 0 8832 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _449_
timestamp 1698431365
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp 1698431365
transform 1 0 6532 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1698431365
transform 1 0 8004 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp 1698431365
transform 1 0 5612 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1698431365
transform 1 0 5796 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1698431365
transform 1 0 3496 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1698431365
transform 1 0 4968 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp 1698431365
transform 1 0 3312 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1698431365
transform 1 0 3220 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1698431365
transform 1 0 15548 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1698431365
transform 1 0 14536 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1698431365
transform 1 0 14260 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1698431365
transform 1 0 10212 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1698431365
transform 1 0 13524 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1698431365
transform 1 0 11408 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1698431365
transform 1 0 8740 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _465_
timestamp 1698431365
transform 1 0 11500 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _466_
timestamp 1698431365
transform 1 0 16100 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _467_
timestamp 1698431365
transform 1 0 14628 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _468_
timestamp 1698431365
transform 1 0 9384 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _469_
timestamp 1698431365
transform 1 0 8096 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _470_
timestamp 1698431365
transform 1 0 7452 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _471_
timestamp 1698431365
transform 1 0 7084 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _472_
timestamp 1698431365
transform 1 0 6716 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _473_
timestamp 1698431365
transform 1 0 4876 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1698431365
transform 1 0 5428 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _475_
timestamp 1698431365
transform 1 0 5060 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _476_
timestamp 1698431365
transform 1 0 10948 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _477_
timestamp 1698431365
transform 1 0 10948 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _478_
timestamp 1698431365
transform 1 0 10856 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _479_
timestamp 1698431365
transform 1 0 8740 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _480_
timestamp 1698431365
transform 1 0 9936 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _481_
timestamp 1698431365
transform 1 0 11316 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1698431365
transform 1 0 11316 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1698431365
transform 1 0 14168 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1698431365
transform 1 0 10856 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1698431365
transform 1 0 7544 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1698431365
transform 1 0 8372 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1698431365
transform 1 0 6532 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1698431365
transform 1 0 16100 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1698431365
transform 1 0 6532 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 11224 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 13616 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15640 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1698431365
transform 1 0 11132 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1698431365
transform 1 0 9384 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1698431365
transform 1 0 8648 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1698431365
transform 1 0 6440 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _497_
timestamp 1698431365
transform 1 0 5796 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _498_
timestamp 1698431365
transform 1 0 3312 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _499_
timestamp 1698431365
transform 1 0 3404 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1698431365
transform 1 0 1104 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1698431365
transform 1 0 3404 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _502_
timestamp 1698431365
transform 1 0 1104 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _503_
timestamp 1698431365
transform 1 0 3312 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp 1698431365
transform 1 0 1288 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _505_
timestamp 1698431365
transform 1 0 1196 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1698431365
transform -1 0 28704 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1698431365
transform -1 0 29440 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1698431365
transform 1 0 29900 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1698431365
transform 1 0 29900 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1698431365
transform -1 0 25760 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1698431365
transform 1 0 25760 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1698431365
transform -1 0 23368 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _513_
timestamp 1698431365
transform 1 0 23828 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _514_
timestamp 1698431365
transform 1 0 19136 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _515_
timestamp 1698431365
transform 1 0 21436 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _516_
timestamp 1698431365
transform 1 0 22908 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _517_
timestamp 1698431365
transform 1 0 21252 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _518_
timestamp 1698431365
transform 1 0 16836 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _519_
timestamp 1698431365
transform 1 0 18676 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _520_
timestamp 1698431365
transform 1 0 17480 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _521_
timestamp 1698431365
transform 1 0 22172 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _522_
timestamp 1698431365
transform 1 0 18860 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _523_
timestamp 1698431365
transform -1 0 20148 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _524_
timestamp 1698431365
transform 1 0 14536 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _525_
timestamp 1698431365
transform 1 0 21712 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _526_
timestamp 1698431365
transform -1 0 16560 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _527_
timestamp 1698431365
transform 1 0 18768 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _528_
timestamp 1698431365
transform 1 0 17664 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _529_
timestamp 1698431365
transform -1 0 18124 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _530_
timestamp 1698431365
transform 1 0 20332 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _531_
timestamp 1698431365
transform 1 0 21252 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _532_
timestamp 1698431365
transform 1 0 22264 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _533_
timestamp 1698431365
transform -1 0 28888 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _534_
timestamp 1698431365
transform -1 0 30452 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _535_
timestamp 1698431365
transform 1 0 29532 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _536_
timestamp 1698431365
transform -1 0 30452 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _537_
timestamp 1698431365
transform -1 0 29348 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _538_
timestamp 1698431365
transform -1 0 26312 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _539_
timestamp 1698431365
transform 1 0 21712 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _540_
timestamp 1698431365
transform 1 0 23000 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _541_
timestamp 1698431365
transform 1 0 20240 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _542_
timestamp 1698431365
transform 1 0 16376 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _543_
timestamp 1698431365
transform 1 0 21252 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _544_
timestamp 1698431365
transform 1 0 16928 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _545_
timestamp 1698431365
transform 1 0 22724 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _546_
timestamp 1698431365
transform 1 0 19228 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _547_
timestamp 1698431365
transform 1 0 22908 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _548_
timestamp 1698431365
transform 1 0 24104 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _549_
timestamp 1698431365
transform -1 0 28152 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _550_
timestamp 1698431365
transform 1 0 29900 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _551_
timestamp 1698431365
transform -1 0 31188 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _552_
timestamp 1698431365
transform 1 0 29624 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _553_
timestamp 1698431365
transform -1 0 28152 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _554_
timestamp 1698431365
transform 1 0 26956 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _555_
timestamp 1698431365
transform 1 0 28980 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _556_
timestamp 1698431365
transform 1 0 29164 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _557_
timestamp 1698431365
transform 1 0 29072 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _558_
timestamp 1698431365
transform -1 0 28336 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _559_
timestamp 1698431365
transform 1 0 24288 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _560_
timestamp 1698431365
transform -1 0 28244 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _561_
timestamp 1698431365
transform 1 0 24288 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _562_
timestamp 1698431365
transform 1 0 23920 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _563_
timestamp 1698431365
transform -1 0 28244 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _564_
timestamp 1698431365
transform 1 0 21712 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _565_
timestamp 1698431365
transform 1 0 18768 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _566_
timestamp 1698431365
transform 1 0 16376 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _567_
timestamp 1698431365
transform 1 0 16744 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _568_
timestamp 1698431365
transform 1 0 15824 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _569_
timestamp 1698431365
transform 1 0 20056 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _624_
timestamp 1698431365
transform -1 0 16192 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _625_
timestamp 1698431365
transform 1 0 16192 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _626_
timestamp 1698431365
transform -1 0 2944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _627_
timestamp 1698431365
transform 1 0 29440 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout7
timestamp 1698431365
transform -1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout8
timestamp 1698431365
transform 1 0 9476 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout9
timestamp 1698431365
transform -1 0 26220 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout10
timestamp 1698431365
transform 1 0 26588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1698431365
transform 1 0 18216 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1698431365
transform 1 0 19872 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 1698431365
transform -1 0 18032 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1698431365
transform -1 0 28060 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1698431365
transform -1 0 27416 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1698431365
transform -1 0 4692 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1698431365
transform 1 0 4416 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1698431365
transform -1 0 9292 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1698431365
transform -1 0 7084 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1698431365
transform 1 0 7084 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1698431365
transform -1 0 9936 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1698431365
transform -1 0 9200 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1698431365
transform -1 0 9568 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1698431365
transform -1 0 15088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16100 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1698431365
transform -1 0 16468 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1698431365
transform -1 0 16008 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1698431365
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1698431365
transform -1 0 23552 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 1698431365
transform -1 0 24196 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout36
timestamp 1698431365
transform -1 0 28888 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1698431365
transform 1 0 29072 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1698431365
transform -1 0 29716 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1698431365
transform -1 0 10304 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout40
timestamp 1698431365
transform 1 0 9936 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1698431365
transform -1 0 26496 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 1698431365
transform -1 0 27968 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1698431365
transform -1 0 28336 0 1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1698431365
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1698431365
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1698431365
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1698431365
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1698431365
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1698431365
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1698431365
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1698431365
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1698431365
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1698431365
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1698431365
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1698431365
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1698431365
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1698431365
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1698431365
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1698431365
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1698431365
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1698431365
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1698431365
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1698431365
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1698431365
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1698431365
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1698431365
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1698431365
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1698431365
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1698431365
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1698431365
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1698431365
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1698431365
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1698431365
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1698431365
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1698431365
transform 1 0 30084 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1698431365
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1698431365
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1698431365
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1698431365
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1698431365
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1698431365
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1698431365
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1698431365
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1698431365
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1698431365
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1698431365
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1698431365
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1698431365
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1698431365
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1698431365
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1698431365
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1698431365
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1698431365
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1698431365
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1698431365
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1698431365
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1698431365
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1698431365
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1698431365
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1698431365
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1698431365
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1698431365
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1698431365
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1698431365
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1698431365
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1698431365
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1698431365
transform 1 0 30820 0 -1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1698431365
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1698431365
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1698431365
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1698431365
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1698431365
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1698431365
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1698431365
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1698431365
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1698431365
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1698431365
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1698431365
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1698431365
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1698431365
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1698431365
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1698431365
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1698431365
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1698431365
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1698431365
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1698431365
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1698431365
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1698431365
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1698431365
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1698431365
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1698431365
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1698431365
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1698431365
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1698431365
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1698431365
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1698431365
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1698431365
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1698431365
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1698431365
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1698431365
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1698431365
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1698431365
transform 1 0 30084 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 1698431365
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1698431365
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1698431365
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1698431365
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1698431365
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1698431365
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1698431365
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1698431365
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1698431365
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1698431365
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1698431365
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1698431365
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1698431365
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1698431365
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1698431365
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1698431365
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1698431365
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1698431365
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1698431365
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1698431365
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1698431365
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1698431365
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1698431365
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1698431365
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1698431365
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1698431365
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1698431365
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1698431365
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1698431365
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1698431365
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1698431365
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1698431365
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1698431365
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1698431365
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1698431365
transform 1 0 30820 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1698431365
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1698431365
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1698431365
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1698431365
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1698431365
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1698431365
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1698431365
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1698431365
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1698431365
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1698431365
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1698431365
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1698431365
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1698431365
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1698431365
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1698431365
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1698431365
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1698431365
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1698431365
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1698431365
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1698431365
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1698431365
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1698431365
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1698431365
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1698431365
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1698431365
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1698431365
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1698431365
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1698431365
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1698431365
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1698431365
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1698431365
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1698431365
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1698431365
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1698431365
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1698431365
transform 1 0 30084 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_333
timestamp 1698431365
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1698431365
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1698431365
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1698431365
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1698431365
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1698431365
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1698431365
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1698431365
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1698431365
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1698431365
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1698431365
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1698431365
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1698431365
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1698431365
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1698431365
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1698431365
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1698431365
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1698431365
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1698431365
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1698431365
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1698431365
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1698431365
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1698431365
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1698431365
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1698431365
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1698431365
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1698431365
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1698431365
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1698431365
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1698431365
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1698431365
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1698431365
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1698431365
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1698431365
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1698431365
transform 1 0 30820 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1698431365
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1698431365
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1698431365
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1698431365
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1698431365
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1698431365
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1698431365
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1698431365
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1698431365
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1698431365
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1698431365
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1698431365
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1698431365
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1698431365
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1698431365
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1698431365
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1698431365
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1698431365
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1698431365
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1698431365
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1698431365
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1698431365
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1698431365
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1698431365
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1698431365
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1698431365
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1698431365
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1698431365
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1698431365
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1698431365
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1698431365
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1698431365
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1698431365
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1698431365
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1698431365
transform 1 0 30084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 1698431365
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1698431365
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1698431365
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1698431365
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1698431365
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1698431365
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1698431365
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1698431365
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1698431365
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1698431365
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1698431365
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1698431365
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1698431365
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1698431365
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1698431365
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1698431365
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1698431365
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1698431365
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1698431365
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1698431365
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1698431365
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1698431365
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1698431365
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1698431365
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1698431365
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1698431365
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1698431365
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1698431365
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1698431365
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1698431365
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1698431365
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1698431365
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1698431365
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1698431365
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1698431365
transform 1 0 30820 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1698431365
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1698431365
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1698431365
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1698431365
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1698431365
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1698431365
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1698431365
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1698431365
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1698431365
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1698431365
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1698431365
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1698431365
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1698431365
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1698431365
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1698431365
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1698431365
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1698431365
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1698431365
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1698431365
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1698431365
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1698431365
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1698431365
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1698431365
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1698431365
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1698431365
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1698431365
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1698431365
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1698431365
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1698431365
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1698431365
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1698431365
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1698431365
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1698431365
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1698431365
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1698431365
transform 1 0 30084 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_333
timestamp 1698431365
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1698431365
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1698431365
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1698431365
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1698431365
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1698431365
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1698431365
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1698431365
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1698431365
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1698431365
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1698431365
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1698431365
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1698431365
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1698431365
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1698431365
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1698431365
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1698431365
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1698431365
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1698431365
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1698431365
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1698431365
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1698431365
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1698431365
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1698431365
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1698431365
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1698431365
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1698431365
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1698431365
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1698431365
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1698431365
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1698431365
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1698431365
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1698431365
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1698431365
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1698431365
transform 1 0 30820 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1698431365
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1698431365
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1698431365
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1698431365
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1698431365
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1698431365
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1698431365
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1698431365
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1698431365
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1698431365
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1698431365
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1698431365
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1698431365
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1698431365
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1698431365
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1698431365
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1698431365
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1698431365
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1698431365
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1698431365
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1698431365
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1698431365
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1698431365
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1698431365
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1698431365
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1698431365
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1698431365
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1698431365
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1698431365
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1698431365
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1698431365
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1698431365
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1698431365
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1698431365
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1698431365
transform 1 0 30084 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_333
timestamp 1698431365
transform 1 0 31188 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1698431365
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1698431365
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1698431365
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1698431365
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1698431365
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1698431365
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1698431365
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1698431365
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1698431365
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1698431365
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1698431365
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1698431365
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1698431365
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1698431365
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1698431365
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1698431365
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1698431365
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1698431365
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1698431365
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1698431365
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1698431365
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1698431365
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1698431365
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1698431365
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1698431365
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1698431365
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1698431365
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1698431365
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1698431365
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1698431365
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1698431365
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1698431365
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1698431365
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1698431365
transform 1 0 30820 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1698431365
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1698431365
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1698431365
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1698431365
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1698431365
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1698431365
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1698431365
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1698431365
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1698431365
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1698431365
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1698431365
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1698431365
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1698431365
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1698431365
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1698431365
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1698431365
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1698431365
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1698431365
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1698431365
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1698431365
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1698431365
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1698431365
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1698431365
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1698431365
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1698431365
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1698431365
transform 1 0 23092 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1698431365
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1698431365
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1698431365
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1698431365
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1698431365
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1698431365
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1698431365
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1698431365
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1698431365
transform 1 0 30084 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 1698431365
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1698431365
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1698431365
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1698431365
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1698431365
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1698431365
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1698431365
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1698431365
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1698431365
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1698431365
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1698431365
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1698431365
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1698431365
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1698431365
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1698431365
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1698431365
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1698431365
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1698431365
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1698431365
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1698431365
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1698431365
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1698431365
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1698431365
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1698431365
transform 1 0 20516 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1698431365
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1698431365
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1698431365
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1698431365
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1698431365
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1698431365
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1698431365
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1698431365
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1698431365
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1698431365
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1698431365
transform 1 0 30820 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1698431365
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1698431365
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1698431365
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1698431365
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1698431365
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1698431365
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1698431365
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1698431365
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1698431365
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1698431365
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1698431365
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1698431365
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1698431365
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1698431365
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1698431365
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1698431365
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1698431365
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1698431365
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1698431365
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1698431365
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1698431365
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1698431365
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1698431365
transform 1 0 19780 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1698431365
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1698431365
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1698431365
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1698431365
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1698431365
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1698431365
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1698431365
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1698431365
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1698431365
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1698431365
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1698431365
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1698431365
transform 1 0 30084 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_333
timestamp 1698431365
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1698431365
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1698431365
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1698431365
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1698431365
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1698431365
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1698431365
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1698431365
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1698431365
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1698431365
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1698431365
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1698431365
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1698431365
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1698431365
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1698431365
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1698431365
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1698431365
transform 1 0 14260 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1698431365
transform 1 0 15364 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1698431365
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1698431365
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1698431365
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1698431365
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1698431365
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1698431365
transform 1 0 20516 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1698431365
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1698431365
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1698431365
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1698431365
transform 1 0 23460 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1698431365
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1698431365
transform 1 0 25668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1698431365
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1698431365
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1698431365
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1698431365
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1698431365
transform 1 0 30820 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1698431365
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1698431365
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1698431365
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1698431365
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1698431365
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1698431365
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1698431365
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1698431365
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1698431365
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1698431365
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1698431365
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1698431365
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_121
timestamp 1698431365
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_126
timestamp 1698431365
transform 1 0 12144 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 12512 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1698431365
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_148
timestamp 1698431365
transform 1 0 14168 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_160
timestamp 1698431365
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_172
timestamp 1698431365
transform 1 0 16376 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_184
timestamp 1698431365
transform 1 0 17480 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1698431365
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1698431365
transform 1 0 19780 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1698431365
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1698431365
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1698431365
transform 1 0 23092 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1698431365
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1698431365
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1698431365
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1698431365
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1698431365
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1698431365
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1698431365
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1698431365
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1698431365
transform 1 0 30084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_333
timestamp 1698431365
transform 1 0 31188 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1698431365
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1698431365
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1698431365
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1698431365
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1698431365
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1698431365
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1698431365
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1698431365
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1698431365
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1698431365
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_105
timestamp 1698431365
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1698431365
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp 1698431365
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_139
timestamp 1698431365
transform 1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1698431365
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_169
timestamp 1698431365
transform 1 0 16100 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_175
timestamp 1698431365
transform 1 0 16652 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_183
timestamp 1698431365
transform 1 0 17388 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_190
timestamp 1698431365
transform 1 0 18032 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_202
timestamp 1698431365
transform 1 0 19136 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_211
timestamp 1698431365
transform 1 0 19964 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1698431365
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_230
timestamp 1698431365
transform 1 0 21712 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_245
timestamp 1698431365
transform 1 0 23092 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_255
timestamp 1698431365
transform 1 0 24012 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_267
timestamp 1698431365
transform 1 0 25116 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1698431365
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1698431365
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1698431365
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1698431365
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1698431365
transform 1 0 30820 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1698431365
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1698431365
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1698431365
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1698431365
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1698431365
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_53
timestamp 1698431365
transform 1 0 5428 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_59
timestamp 1698431365
transform 1 0 5980 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_63
timestamp 1698431365
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_88
timestamp 1698431365
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_116
timestamp 1698431365
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_121
timestamp 1698431365
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_128
timestamp 1698431365
transform 1 0 12328 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_148
timestamp 1698431365
transform 1 0 14168 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_157
timestamp 1698431365
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_169
timestamp 1698431365
transform 1 0 16100 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_197
timestamp 1698431365
transform 1 0 18676 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_218
timestamp 1698431365
transform 1 0 20608 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_222
timestamp 1698431365
transform 1 0 20976 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1698431365
transform 1 0 23552 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_253
timestamp 1698431365
transform 1 0 23828 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_278
timestamp 1698431365
transform 1 0 26128 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_290
timestamp 1698431365
transform 1 0 27232 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_294
timestamp 1698431365
transform 1 0 27600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_306
timestamp 1698431365
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1698431365
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1698431365
transform 1 0 30084 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_333
timestamp 1698431365
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1698431365
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_15
timestamp 1698431365
transform 1 0 1932 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1698431365
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_80
timestamp 1698431365
transform 1 0 7912 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_88
timestamp 1698431365
transform 1 0 8648 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1698431365
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1698431365
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1698431365
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1698431365
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_143
timestamp 1698431365
transform 1 0 13708 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_164
timestamp 1698431365
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1698431365
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_178
timestamp 1698431365
transform 1 0 16928 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1698431365
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_205
timestamp 1698431365
transform 1 0 19412 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 19780 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_216
timestamp 1698431365
transform 1 0 20424 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_235
timestamp 1698431365
transform 1 0 22172 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_259
timestamp 1698431365
transform 1 0 24380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_267
timestamp 1698431365
transform 1 0 25116 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_271
timestamp 1698431365
transform 1 0 25484 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_301
timestamp 1698431365
transform 1 0 28244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_306
timestamp 1698431365
transform 1 0 28704 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_314
timestamp 1698431365
transform 1 0 29440 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_326
timestamp 1698431365
transform 1 0 30544 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_334
timestamp 1698431365
transform 1 0 31280 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1698431365
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1698431365
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1698431365
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1698431365
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_41
timestamp 1698431365
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_46
timestamp 1698431365
transform 1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_55
timestamp 1698431365
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_70
timestamp 1698431365
transform 1 0 6992 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_74
timestamp 1698431365
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1698431365
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_111
timestamp 1698431365
transform 1 0 10764 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_119
timestamp 1698431365
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_125
timestamp 1698431365
transform 1 0 12052 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1698431365
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_148
timestamp 1698431365
transform 1 0 14168 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_158
timestamp 1698431365
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_174
timestamp 1698431365
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_200
timestamp 1698431365
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_218
timestamp 1698431365
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_243
timestamp 1698431365
transform 1 0 22908 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1698431365
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_253
timestamp 1698431365
transform 1 0 23828 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_259
timestamp 1698431365
transform 1 0 24380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_268
timestamp 1698431365
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_273
timestamp 1698431365
transform 1 0 25668 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_281
timestamp 1698431365
transform 1 0 26404 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_309
timestamp 1698431365
transform 1 0 28980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_317
timestamp 1698431365
transform 1 0 29716 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_323
timestamp 1698431365
transform 1 0 30268 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1698431365
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_15
timestamp 1698431365
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_29
timestamp 1698431365
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 1698431365
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_63
timestamp 1698431365
transform 1 0 6348 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_74
timestamp 1698431365
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_86
timestamp 1698431365
transform 1 0 8464 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_101
timestamp 1698431365
transform 1 0 9844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1698431365
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_129
timestamp 1698431365
transform 1 0 12420 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_135
timestamp 1698431365
transform 1 0 12972 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1698431365
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_180
timestamp 1698431365
transform 1 0 17112 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_194
timestamp 1698431365
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_213
timestamp 1698431365
transform 1 0 20148 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 1698431365
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_241
timestamp 1698431365
transform 1 0 22724 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_245
timestamp 1698431365
transform 1 0 23092 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_250
timestamp 1698431365
transform 1 0 23552 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_278
timestamp 1698431365
transform 1 0 26128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_308
timestamp 1698431365
transform 1 0 28888 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_330
timestamp 1698431365
transform 1 0 30912 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_334
timestamp 1698431365
transform 1 0 31280 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1698431365
transform 1 0 828 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_12
timestamp 1698431365
transform 1 0 1656 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_20
timestamp 1698431365
transform 1 0 2392 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1698431365
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_38
timestamp 1698431365
transform 1 0 4048 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_44
timestamp 1698431365
transform 1 0 4600 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_53
timestamp 1698431365
transform 1 0 5428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_64
timestamp 1698431365
transform 1 0 6440 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1698431365
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_89
timestamp 1698431365
transform 1 0 8740 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_106
timestamp 1698431365
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1698431365
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1698431365
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_165
timestamp 1698431365
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1698431365
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_209
timestamp 1698431365
transform 1 0 19780 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_232
timestamp 1698431365
transform 1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_253
timestamp 1698431365
transform 1 0 23828 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_272
timestamp 1698431365
transform 1 0 25576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_279
timestamp 1698431365
transform 1 0 26220 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_285
timestamp 1698431365
transform 1 0 26772 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1698431365
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_301
timestamp 1698431365
transform 1 0 28244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_309
timestamp 1698431365
transform 1 0 28980 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_333
timestamp 1698431365
transform 1 0 31188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_3
timestamp 1698431365
transform 1 0 828 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_29
timestamp 1698431365
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1698431365
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1698431365
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_64
timestamp 1698431365
transform 1 0 6440 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_97
timestamp 1698431365
transform 1 0 9476 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1698431365
transform 1 0 10580 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp 1698431365
transform 1 0 10948 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_117
timestamp 1698431365
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_129
timestamp 1698431365
transform 1 0 12420 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_164
timestamp 1698431365
transform 1 0 15640 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1698431365
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_181
timestamp 1698431365
transform 1 0 17204 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_200
timestamp 1698431365
transform 1 0 18952 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_211
timestamp 1698431365
transform 1 0 19964 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1698431365
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_228
timestamp 1698431365
transform 1 0 21528 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_248
timestamp 1698431365
transform 1 0 23368 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_256
timestamp 1698431365
transform 1 0 24104 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_274
timestamp 1698431365
transform 1 0 25760 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_281
timestamp 1698431365
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_305
timestamp 1698431365
transform 1 0 28612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_316
timestamp 1698431365
transform 1 0 29624 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_325
timestamp 1698431365
transform 1 0 30452 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_333
timestamp 1698431365
transform 1 0 31188 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_10
timestamp 1698431365
transform 1 0 1472 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_22
timestamp 1698431365
transform 1 0 2576 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_29
timestamp 1698431365
transform 1 0 3220 0 1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1698431365
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_53
timestamp 1698431365
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_71
timestamp 1698431365
transform 1 0 7084 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1698431365
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_88
timestamp 1698431365
transform 1 0 8648 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_96
timestamp 1698431365
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_115
timestamp 1698431365
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1698431365
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1698431365
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 1698431365
transform 1 0 13524 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_147
timestamp 1698431365
transform 1 0 14076 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_151
timestamp 1698431365
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_169
timestamp 1698431365
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1698431365
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1698431365
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_209
timestamp 1698431365
transform 1 0 19780 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_217
timestamp 1698431365
transform 1 0 20516 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_225
timestamp 1698431365
transform 1 0 21252 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_233
timestamp 1698431365
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1698431365
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_253
timestamp 1698431365
transform 1 0 23828 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_278
timestamp 1698431365
transform 1 0 26128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_282
timestamp 1698431365
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_287
timestamp 1698431365
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_299
timestamp 1698431365
transform 1 0 28060 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_309
timestamp 1698431365
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_331
timestamp 1698431365
transform 1 0 31004 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_3
timestamp 1698431365
transform 1 0 828 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_30
timestamp 1698431365
transform 1 0 3312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_37
timestamp 1698431365
transform 1 0 3956 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_44
timestamp 1698431365
transform 1 0 4600 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_73
timestamp 1698431365
transform 1 0 7268 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_92
timestamp 1698431365
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1698431365
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 1698431365
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_121
timestamp 1698431365
transform 1 0 11684 0 -1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_150
timestamp 1698431365
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 1698431365
transform 1 0 15732 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_185
timestamp 1698431365
transform 1 0 17572 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_197
timestamp 1698431365
transform 1 0 18676 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_219
timestamp 1698431365
transform 1 0 20700 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1698431365
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_241
timestamp 1698431365
transform 1 0 22724 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_253
timestamp 1698431365
transform 1 0 23828 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_257
timestamp 1698431365
transform 1 0 24196 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_274
timestamp 1698431365
transform 1 0 25760 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_288
timestamp 1698431365
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_300
timestamp 1698431365
transform 1 0 28152 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_306
timestamp 1698431365
transform 1 0 28704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_318
timestamp 1698431365
transform 1 0 29808 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1698431365
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_15
timestamp 1698431365
transform 1 0 1932 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_23
timestamp 1698431365
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1698431365
transform 1 0 3220 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_50
timestamp 1698431365
transform 1 0 5152 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_69
timestamp 1698431365
transform 1 0 6900 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1698431365
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_92
timestamp 1698431365
transform 1 0 9016 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_128
timestamp 1698431365
transform 1 0 12328 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_149
timestamp 1698431365
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_187
timestamp 1698431365
transform 1 0 17756 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1698431365
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_205
timestamp 1698431365
transform 1 0 19412 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_211
timestamp 1698431365
transform 1 0 19964 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_231
timestamp 1698431365
transform 1 0 21804 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_250
timestamp 1698431365
transform 1 0 23552 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_269
timestamp 1698431365
transform 1 0 25300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_273
timestamp 1698431365
transform 1 0 25668 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_306
timestamp 1698431365
transform 1 0 28704 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1698431365
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1698431365
transform 1 0 30084 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_333
timestamp 1698431365
transform 1 0 31188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_3
timestamp 1698431365
transform 1 0 828 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_9
timestamp 1698431365
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_22
timestamp 1698431365
transform 1 0 2576 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_30
timestamp 1698431365
transform 1 0 3312 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_37
timestamp 1698431365
transform 1 0 3956 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1698431365
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1698431365
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_69
timestamp 1698431365
transform 1 0 6900 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_102
timestamp 1698431365
transform 1 0 9936 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1698431365
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_129
timestamp 1698431365
transform 1 0 12420 0 -1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_154
timestamp 1698431365
transform 1 0 14720 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1698431365
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_179
timestamp 1698431365
transform 1 0 17020 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_215
timestamp 1698431365
transform 1 0 20332 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1698431365
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_230
timestamp 1698431365
transform 1 0 21712 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_241
timestamp 1698431365
transform 1 0 22724 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_260
timestamp 1698431365
transform 1 0 24472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_281
timestamp 1698431365
transform 1 0 26404 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_290
timestamp 1698431365
transform 1 0 27232 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_318
timestamp 1698431365
transform 1 0 29808 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_3
timestamp 1698431365
transform 1 0 828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1698431365
transform 1 0 3220 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_46
timestamp 1698431365
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_64
timestamp 1698431365
transform 1 0 6440 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1698431365
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_121
timestamp 1698431365
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_141
timestamp 1698431365
transform 1 0 13524 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_152
timestamp 1698431365
transform 1 0 14536 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_156
timestamp 1698431365
transform 1 0 14904 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_182
timestamp 1698431365
transform 1 0 17296 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_187
timestamp 1698431365
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1698431365
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1698431365
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_226
timestamp 1698431365
transform 1 0 21344 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_233
timestamp 1698431365
transform 1 0 21988 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1698431365
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_253
timestamp 1698431365
transform 1 0 23828 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_272
timestamp 1698431365
transform 1 0 25576 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_300
timestamp 1698431365
transform 1 0 28152 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_325
timestamp 1698431365
transform 1 0 30452 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_333
timestamp 1698431365
transform 1 0 31188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_3
timestamp 1698431365
transform 1 0 828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_12
timestamp 1698431365
transform 1 0 1656 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_24
timestamp 1698431365
transform 1 0 2760 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_48
timestamp 1698431365
transform 1 0 4968 0 -1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1698431365
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_69
timestamp 1698431365
transform 1 0 6900 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_80
timestamp 1698431365
transform 1 0 7912 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_92
timestamp 1698431365
transform 1 0 9016 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 1698431365
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_116
timestamp 1698431365
transform 1 0 11224 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_128
timestamp 1698431365
transform 1 0 12328 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_146
timestamp 1698431365
transform 1 0 13984 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_158
timestamp 1698431365
transform 1 0 15088 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_162
timestamp 1698431365
transform 1 0 15456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_169
timestamp 1698431365
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_195
timestamp 1698431365
transform 1 0 18492 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_214
timestamp 1698431365
transform 1 0 20240 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1698431365
transform 1 0 20976 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_225
timestamp 1698431365
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_236
timestamp 1698431365
transform 1 0 22264 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_247
timestamp 1698431365
transform 1 0 23276 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_264
timestamp 1698431365
transform 1 0 24840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 26128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_302
timestamp 1698431365
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_318
timestamp 1698431365
transform 1 0 29808 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_3
timestamp 1698431365
transform 1 0 828 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1698431365
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_45
timestamp 1698431365
transform 1 0 4692 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_65
timestamp 1698431365
transform 1 0 6532 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_74
timestamp 1698431365
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_79
timestamp 1698431365
transform 1 0 7820 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1698431365
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_101
timestamp 1698431365
transform 1 0 9844 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_129
timestamp 1698431365
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1698431365
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 1698431365
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_207
timestamp 1698431365
transform 1 0 19596 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_246
timestamp 1698431365
transform 1 0 23184 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_253
timestamp 1698431365
transform 1 0 23828 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_265
timestamp 1698431365
transform 1 0 24932 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_273
timestamp 1698431365
transform 1 0 25668 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_282
timestamp 1698431365
transform 1 0 26496 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_313
timestamp 1698431365
transform 1 0 29348 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_320
timestamp 1698431365
transform 1 0 29992 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_332
timestamp 1698431365
transform 1 0 31096 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_3
timestamp 1698431365
transform 1 0 828 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_7
timestamp 1698431365
transform 1 0 1196 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_12
timestamp 1698431365
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_24
timestamp 1698431365
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_36
timestamp 1698431365
transform 1 0 3864 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1698431365
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_60
timestamp 1698431365
transform 1 0 6072 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1698431365
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_120
timestamp 1698431365
transform 1 0 11592 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_132
timestamp 1698431365
transform 1 0 12696 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_145
timestamp 1698431365
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_149
timestamp 1698431365
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_159
timestamp 1698431365
transform 1 0 15180 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_163
timestamp 1698431365
transform 1 0 15548 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1698431365
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_169
timestamp 1698431365
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_177
timestamp 1698431365
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_194
timestamp 1698431365
transform 1 0 18400 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_200
timestamp 1698431365
transform 1 0 18952 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_220
timestamp 1698431365
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1698431365
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_237
timestamp 1698431365
transform 1 0 22356 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_267
timestamp 1698431365
transform 1 0 25116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 1698431365
transform 1 0 25852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_301
timestamp 1698431365
transform 1 0 28244 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_312
timestamp 1698431365
transform 1 0 29256 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_332
timestamp 1698431365
transform 1 0 31096 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1698431365
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1698431365
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1698431365
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1698431365
transform 1 0 3220 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_49
timestamp 1698431365
transform 1 0 5060 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_56
timestamp 1698431365
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_65
timestamp 1698431365
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_78
timestamp 1698431365
transform 1 0 7728 0 1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1698431365
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_97
timestamp 1698431365
transform 1 0 9476 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_111
timestamp 1698431365
transform 1 0 10764 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_131
timestamp 1698431365
transform 1 0 12604 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1698431365
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_157
timestamp 1698431365
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_169
timestamp 1698431365
transform 1 0 16100 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_181
timestamp 1698431365
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_189
timestamp 1698431365
transform 1 0 17940 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_208
timestamp 1698431365
transform 1 0 19688 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_219
timestamp 1698431365
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_224
timestamp 1698431365
transform 1 0 21160 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_232
timestamp 1698431365
transform 1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_249
timestamp 1698431365
transform 1 0 23460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_253
timestamp 1698431365
transform 1 0 23828 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_266
timestamp 1698431365
transform 1 0 25024 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_274
timestamp 1698431365
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_280
timestamp 1698431365
transform 1 0 26312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_295
timestamp 1698431365
transform 1 0 27692 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_303
timestamp 1698431365
transform 1 0 28428 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 29348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_331
timestamp 1698431365
transform 1 0 31004 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1698431365
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_15
timestamp 1698431365
transform 1 0 1932 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_21
timestamp 1698431365
transform 1 0 2484 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_26
timestamp 1698431365
transform 1 0 2944 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1698431365
transform 1 0 5796 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_70
timestamp 1698431365
transform 1 0 6992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_87
timestamp 1698431365
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1698431365
transform 1 0 10948 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_117
timestamp 1698431365
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_129
timestamp 1698431365
transform 1 0 12420 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_155
timestamp 1698431365
transform 1 0 14812 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1698431365
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_188
timestamp 1698431365
transform 1 0 17848 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_200
timestamp 1698431365
transform 1 0 18952 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_204
timestamp 1698431365
transform 1 0 19320 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1698431365
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_247
timestamp 1698431365
transform 1 0 23276 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_263
timestamp 1698431365
transform 1 0 24748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_267
timestamp 1698431365
transform 1 0 25116 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_299
timestamp 1698431365
transform 1 0 28060 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_305
timestamp 1698431365
transform 1 0 28612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_312
timestamp 1698431365
transform 1 0 29256 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_316
timestamp 1698431365
transform 1 0 29624 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_333
timestamp 1698431365
transform 1 0 31188 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1698431365
transform 1 0 828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1698431365
transform 1 0 1932 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1698431365
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_45
timestamp 1698431365
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_75
timestamp 1698431365
transform 1 0 7452 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1698431365
transform 1 0 8188 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_85
timestamp 1698431365
transform 1 0 8372 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_97
timestamp 1698431365
transform 1 0 9476 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_105
timestamp 1698431365
transform 1 0 10212 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_117
timestamp 1698431365
transform 1 0 11316 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_134
timestamp 1698431365
transform 1 0 12880 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_146
timestamp 1698431365
transform 1 0 13984 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_174
timestamp 1698431365
transform 1 0 16560 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_182
timestamp 1698431365
transform 1 0 17296 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1698431365
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_200
timestamp 1698431365
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_222
timestamp 1698431365
transform 1 0 20976 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_230
timestamp 1698431365
transform 1 0 21712 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_235
timestamp 1698431365
transform 1 0 22172 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_253
timestamp 1698431365
transform 1 0 23828 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_269
timestamp 1698431365
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_281
timestamp 1698431365
transform 1 0 26404 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_294
timestamp 1698431365
transform 1 0 27600 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_306
timestamp 1698431365
transform 1 0 28704 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_326
timestamp 1698431365
transform 1 0 30544 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_334
timestamp 1698431365
transform 1 0 31280 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1698431365
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_15
timestamp 1698431365
transform 1 0 1932 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_23
timestamp 1698431365
transform 1 0 2668 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_32
timestamp 1698431365
transform 1 0 3496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_37
timestamp 1698431365
transform 1 0 3956 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1698431365
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_61
timestamp 1698431365
transform 1 0 6164 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_81
timestamp 1698431365
transform 1 0 8004 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_96
timestamp 1698431365
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1698431365
transform 1 0 10304 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_113
timestamp 1698431365
transform 1 0 10948 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_133
timestamp 1698431365
transform 1 0 12788 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_150
timestamp 1698431365
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_205
timestamp 1698431365
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 1698431365
transform 1 0 20792 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_281
timestamp 1698431365
transform 1 0 26404 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_300
timestamp 1698431365
transform 1 0 28152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_308
timestamp 1698431365
transform 1 0 28888 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_320
timestamp 1698431365
transform 1 0 29992 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_332
timestamp 1698431365
transform 1 0 31096 0 -1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1698431365
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1698431365
transform 1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1698431365
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1698431365
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_41
timestamp 1698431365
transform 1 0 4324 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_50
timestamp 1698431365
transform 1 0 5152 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_58
timestamp 1698431365
transform 1 0 5888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_62
timestamp 1698431365
transform 1 0 6256 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_66
timestamp 1698431365
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1698431365
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_85
timestamp 1698431365
transform 1 0 8372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_95
timestamp 1698431365
transform 1 0 9292 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_124
timestamp 1698431365
transform 1 0 11960 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_132
timestamp 1698431365
transform 1 0 12696 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1698431365
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_146
timestamp 1698431365
transform 1 0 13984 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_167
timestamp 1698431365
transform 1 0 15916 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_194
timestamp 1698431365
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_197
timestamp 1698431365
transform 1 0 18676 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_207
timestamp 1698431365
transform 1 0 19596 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_211
timestamp 1698431365
transform 1 0 19964 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_218
timestamp 1698431365
transform 1 0 20608 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_222
timestamp 1698431365
transform 1 0 20976 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_246
timestamp 1698431365
transform 1 0 23184 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_253
timestamp 1698431365
transform 1 0 23828 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_259
timestamp 1698431365
transform 1 0 24380 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_271
timestamp 1698431365
transform 1 0 25484 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_282
timestamp 1698431365
transform 1 0 26496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_293
timestamp 1698431365
transform 1 0 27508 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_297
timestamp 1698431365
transform 1 0 27876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1698431365
transform 1 0 28796 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_325
timestamp 1698431365
transform 1 0 30452 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_333
timestamp 1698431365
transform 1 0 31188 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1698431365
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1698431365
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1698431365
transform 1 0 3036 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1698431365
transform 1 0 4140 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1698431365
transform 1 0 5244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1698431365
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1698431365
transform 1 0 5796 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1698431365
transform 1 0 6900 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_81
timestamp 1698431365
transform 1 0 8004 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 1698431365
transform 1 0 10488 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_119
timestamp 1698431365
transform 1 0 11500 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_126
timestamp 1698431365
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_172
timestamp 1698431365
transform 1 0 16376 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_197
timestamp 1698431365
transform 1 0 18676 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_202
timestamp 1698431365
transform 1 0 19136 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_238
timestamp 1698431365
transform 1 0 22448 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_260
timestamp 1698431365
transform 1 0 24472 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_266
timestamp 1698431365
transform 1 0 25024 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_270
timestamp 1698431365
transform 1 0 25392 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_296
timestamp 1698431365
transform 1 0 27784 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_320
timestamp 1698431365
transform 1 0 29992 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_332
timestamp 1698431365
transform 1 0 31096 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_6
timestamp 1698431365
transform 1 0 1104 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_10
timestamp 1698431365
transform 1 0 1472 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_14
timestamp 1698431365
transform 1 0 1840 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_18
timestamp 1698431365
transform 1 0 2208 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_22
timestamp 1698431365
transform 1 0 2576 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_32
timestamp 1698431365
transform 1 0 3496 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_38
timestamp 1698431365
transform 1 0 4048 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_42
timestamp 1698431365
transform 1 0 4416 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_46
timestamp 1698431365
transform 1 0 4784 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_50
timestamp 1698431365
transform 1 0 5152 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_54
timestamp 1698431365
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 1698431365
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_62
timestamp 1698431365
transform 1 0 6256 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_66
timestamp 1698431365
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_70
timestamp 1698431365
transform 1 0 6992 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_74
timestamp 1698431365
transform 1 0 7360 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_78
timestamp 1698431365
transform 1 0 7728 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 1698431365
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_98
timestamp 1698431365
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_102
timestamp 1698431365
transform 1 0 9936 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_106
timestamp 1698431365
transform 1 0 10304 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_110
timestamp 1698431365
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_113
timestamp 1698431365
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_118
timestamp 1698431365
transform 1 0 11408 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_135
timestamp 1698431365
transform 1 0 12972 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1698431365
transform 1 0 13340 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_141
timestamp 1698431365
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_158
timestamp 1698431365
transform 1 0 15088 0 1 21216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_173
timestamp 1698431365
transform 1 0 16468 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_185
timestamp 1698431365
transform 1 0 17572 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1698431365
transform 1 0 18308 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_213
timestamp 1698431365
transform 1 0 20148 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_221
timestamp 1698431365
transform 1 0 20884 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_228
timestamp 1698431365
transform 1 0 21528 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1698431365
transform 1 0 23552 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_257
timestamp 1698431365
transform 1 0 24196 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_265
timestamp 1698431365
transform 1 0 24932 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_271
timestamp 1698431365
transform 1 0 25484 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_278
timestamp 1698431365
transform 1 0 26128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_281
timestamp 1698431365
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_287
timestamp 1698431365
transform 1 0 26956 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_293
timestamp 1698431365
transform 1 0 27508 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1698431365
transform 1 0 28704 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1698431365
transform 1 0 30084 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_333
timestamp 1698431365
transform 1 0 31188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 29808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1698431365
transform -1 0 29808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1698431365
transform -1 0 28704 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 29256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1698431365
transform -1 0 26956 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1698431365
transform 1 0 25852 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap11
timestamp 1698431365
transform 1 0 11408 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap12
timestamp 1698431365
transform 1 0 5428 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap13
timestamp 1698431365
transform 1 0 5060 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap24
timestamp 1698431365
transform -1 0 27692 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap25
timestamp 1698431365
transform -1 0 26128 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1698431365
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1698431365
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1698431365
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1698431365
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1698431365
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1698431365
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1698431365
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1698431365
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1698431365
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1698431365
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1698431365
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1698431365
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1698431365
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1698431365
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1698431365
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1698431365
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1698431365
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1698431365
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1698431365
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1698431365
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1698431365
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1698431365
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1698431365
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1698431365
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1698431365
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1698431365
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1698431365
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1698431365
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1698431365
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1698431365
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1698431365
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1698431365
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1698431365
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1698431365
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1698431365
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1698431365
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1698431365
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1698431365
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1698431365
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1698431365
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1698431365
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1698431365
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1698431365
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1698431365
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1698431365
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1698431365
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1698431365
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1698431365
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1698431365
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1698431365
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1698431365
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1698431365
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1698431365
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1698431365
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1698431365
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1698431365
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1698431365
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1698431365
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1698431365
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1698431365
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1698431365
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1698431365
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1698431365
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1698431365
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1698431365
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1698431365
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1698431365
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1698431365
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1698431365
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1698431365
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1698431365
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1698431365
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1698431365
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1698431365
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1698431365
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1698431365
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1698431365
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1698431365
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1698431365
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1698431365
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1698431365
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1698431365
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1698431365
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1698431365
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1698431365
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1698431365
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1698431365
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1698431365
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1698431365
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1698431365
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1698431365
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1698431365
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1698431365
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1698431365
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1698431365
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1698431365
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1698431365
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1698431365
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1698431365
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1698431365
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1698431365
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1698431365
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1698431365
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1698431365
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1698431365
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1698431365
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1698431365
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1698431365
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1698431365
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1698431365
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1698431365
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1698431365
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1698431365
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1698431365
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1698431365
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1698431365
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1698431365
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1698431365
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1698431365
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1698431365
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1698431365
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1698431365
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1698431365
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1698431365
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1698431365
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1698431365
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1698431365
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1698431365
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1698431365
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1698431365
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1698431365
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1698431365
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1698431365
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1698431365
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1698431365
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1698431365
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1698431365
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1698431365
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1698431365
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1698431365
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1698431365
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1698431365
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1698431365
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1698431365
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1698431365
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1698431365
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1698431365
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1698431365
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1698431365
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1698431365
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1698431365
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1698431365
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1698431365
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1698431365
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1698431365
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1698431365
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1698431365
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1698431365
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1698431365
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1698431365
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1698431365
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1698431365
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1698431365
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1698431365
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1698431365
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1698431365
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1698431365
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1698431365
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1698431365
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1698431365
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1698431365
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1698431365
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1698431365
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1698431365
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1698431365
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1698431365
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1698431365
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1698431365
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1698431365
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1698431365
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1698431365
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1698431365
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1698431365
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1698431365
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1698431365
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1698431365
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1698431365
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1698431365
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1698431365
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1698431365
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1698431365
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1698431365
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1698431365
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1698431365
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1698431365
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1698431365
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1698431365
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1698431365
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1698431365
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1698431365
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1698431365
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1698431365
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1698431365
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1698431365
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1698431365
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1698431365
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1698431365
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1698431365
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1698431365
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1698431365
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1698431365
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1698431365
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1698431365
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1698431365
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1698431365
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1698431365
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1698431365
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1698431365
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1698431365
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1698431365
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1698431365
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1698431365
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1698431365
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1698431365
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1698431365
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1698431365
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1698431365
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1698431365
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1698431365
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1698431365
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1698431365
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1698431365
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1698431365
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1698431365
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1698431365
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1698431365
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1698431365
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1698431365
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1698431365
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1698431365
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1698431365
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1698431365
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1698431365
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1698431365
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1698431365
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1698431365
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1698431365
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1698431365
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1698431365
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1698431365
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1698431365
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1698431365
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1698431365
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1698431365
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1698431365
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1698431365
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1698431365
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1698431365
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1698431365
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1698431365
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1698431365
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1698431365
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1698431365
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  tdc0.g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 4784 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[0\].dly_stp
timestamp 1698431365
transform 1 0 3220 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[1\].dly_stp
timestamp 1698431365
transform -1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[2\].dly_stp
timestamp 1698431365
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_dly_stp\[3\].dly_stp
timestamp 1698431365
transform -1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  tdc0.g_dly_stp\[4\].dly_stp
timestamp 1698431365
transform 1 0 3680 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[1\].g_buf1.ctr_buf
timestamp 1698431365
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[1\].stg01
timestamp 1698431365
transform -1 0 5060 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[1\].stg02 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 5152 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[2\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 11316 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[2\].stg01
timestamp 1698431365
transform 1 0 11316 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[2\].stg02
timestamp 1698431365
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[3\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 10396 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[3\].stg01
timestamp 1698431365
transform -1 0 10764 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[3\].stg02
timestamp 1698431365
transform 1 0 10304 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[4\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 12604 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[4\].stg01
timestamp 1698431365
transform 1 0 9476 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[4\].stg02
timestamp 1698431365
transform -1 0 10120 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[5\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 10580 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[5\].stg01
timestamp 1698431365
transform 1 0 10028 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[5\].stg02
timestamp 1698431365
transform 1 0 9292 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[6\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 8924 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[6\].stg01
timestamp 1698431365
transform 1 0 9200 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[6\].stg02
timestamp 1698431365
transform 1 0 9016 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[7\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 11500 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[7\].stg01
timestamp 1698431365
transform 1 0 8648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[7\].stg02
timestamp 1698431365
transform -1 0 10212 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[8\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 15732 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[8\].stg01
timestamp 1698431365
transform 1 0 10948 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[8\].stg02
timestamp 1698431365
transform 1 0 10580 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[9\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 14444 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[9\].stg01
timestamp 1698431365
transform 1 0 11408 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[9\].stg02
timestamp 1698431365
transform 1 0 10764 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[10\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 9384 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[10\].stg01
timestamp 1698431365
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[10\].stg02
timestamp 1698431365
transform 1 0 9844 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[11\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 8096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[11\].stg01
timestamp 1698431365
transform 1 0 8740 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[11\].stg02
timestamp 1698431365
transform 1 0 7820 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[12\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 7728 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[12\].stg01
timestamp 1698431365
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[12\].stg02
timestamp 1698431365
transform 1 0 7544 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[13\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 7176 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[13\].stg01
timestamp 1698431365
transform 1 0 6164 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[13\].stg02
timestamp 1698431365
transform -1 0 7452 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[14\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 6532 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[14\].stg01
timestamp 1698431365
transform 1 0 5980 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[14\].stg02
timestamp 1698431365
transform 1 0 6624 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[15\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 5152 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[15\].stg01
timestamp 1698431365
transform -1 0 7452 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[15\].stg02
timestamp 1698431365
transform 1 0 5336 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring1\[16\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 5336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring1\[16\].stg01
timestamp 1698431365
transform -1 0 5060 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring1\[16\].stg02
timestamp 1698431365
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring1\[16\].stg02_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[16\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 5612 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[16\].stg01_45
timestamp 1698431365
transform -1 0 4784 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[16\].stg01
timestamp 1698431365
transform -1 0 4048 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[16\].stg02
timestamp 1698431365
transform -1 0 4784 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[17\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 5060 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[17\].stg01_46
timestamp 1698431365
transform 1 0 4140 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[17\].stg01
timestamp 1698431365
transform -1 0 4508 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[17\].stg02
timestamp 1698431365
transform -1 0 5520 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[18\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 10948 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[18\].stg01_47
timestamp 1698431365
transform 1 0 5152 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[18\].stg01
timestamp 1698431365
transform -1 0 6072 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[18\].stg02
timestamp 1698431365
transform -1 0 10672 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[19\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 10764 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[19\].stg01_48
timestamp 1698431365
transform -1 0 11224 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[19\].stg01
timestamp 1698431365
transform -1 0 10672 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[19\].stg02
timestamp 1698431365
transform 1 0 9936 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[20\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[20\].stg01_49
timestamp 1698431365
transform 1 0 8924 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[20\].stg01
timestamp 1698431365
transform 1 0 9200 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[20\].stg02
timestamp 1698431365
transform -1 0 10488 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[21\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 9016 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[21\].stg01
timestamp 1698431365
transform 1 0 9568 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[21\].stg01_50
timestamp 1698431365
transform 1 0 9016 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[21\].stg02
timestamp 1698431365
transform -1 0 10028 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[22\].g_buf1.ctr_buf
timestamp 1698431365
transform 1 0 10212 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[22\].stg01_51
timestamp 1698431365
transform 1 0 8372 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[22\].stg01
timestamp 1698431365
transform 1 0 8924 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[22\].stg02
timestamp 1698431365
transform -1 0 9016 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[23\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 11316 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[23\].stg01_52
timestamp 1698431365
transform 1 0 9384 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[23\].stg01
timestamp 1698431365
transform 1 0 9660 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[23\].stg02
timestamp 1698431365
transform -1 0 9936 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[24\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 11408 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[24\].stg01_53
timestamp 1698431365
transform -1 0 11960 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[24\].stg01
timestamp 1698431365
transform -1 0 10856 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[24\].stg02
timestamp 1698431365
transform -1 0 11316 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[25\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 11316 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[25\].stg01_54
timestamp 1698431365
transform 1 0 9844 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[25\].stg01
timestamp 1698431365
transform 1 0 10120 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[25\].stg02
timestamp 1698431365
transform -1 0 10764 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[26\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[26\].stg01_55
timestamp 1698431365
transform -1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[26\].stg01
timestamp 1698431365
transform -1 0 9844 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[26\].stg02
timestamp 1698431365
transform 1 0 9476 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[27\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 7544 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[27\].stg01
timestamp 1698431365
transform -1 0 7820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[27\].stg01_56
timestamp 1698431365
transform -1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[27\].stg02
timestamp 1698431365
transform -1 0 8740 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[28\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 7820 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[28\].stg01
timestamp 1698431365
transform -1 0 7544 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[28\].stg01_57
timestamp 1698431365
transform -1 0 7820 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[28\].stg02
timestamp 1698431365
transform 1 0 7176 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[29\].g_buf1.ctr_buf
timestamp 1698431365
transform 1 0 7084 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[29\].stg01_58
timestamp 1698431365
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[29\].stg01
timestamp 1698431365
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[29\].stg02
timestamp 1698431365
transform -1 0 7084 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[30\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 6900 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[30\].stg01_59
timestamp 1698431365
transform 1 0 5980 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[30\].stg01
timestamp 1698431365
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[30\].stg02
timestamp 1698431365
transform -1 0 6624 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc0.g_ring3\[31\].g_buf1.ctr_buf
timestamp 1698431365
transform -1 0 6256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc0.g_ring3\[31\].stg01_60
timestamp 1698431365
transform 1 0 5888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.g_ring3\[31\].stg01
timestamp 1698431365
transform 1 0 6348 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.g_ring3\[31\].stg02
timestamp 1698431365
transform 1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tdc0.stg01_61
timestamp 1698431365
transform -1 0 4324 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc0.stg01
timestamp 1698431365
transform -1 0 4048 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc0.stg02
timestamp 1698431365
transform -1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  tdc1.g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 26496 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[0\].dly_stp
timestamp 1698431365
transform -1 0 15548 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[1\].dly_stp
timestamp 1698431365
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[2\].dly_stp
timestamp 1698431365
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_dly_stp\[3\].dly_stp
timestamp 1698431365
transform -1 0 16560 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  tdc1.g_dly_stp\[4\].dly_stp
timestamp 1698431365
transform 1 0 16560 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[1\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 19136 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[1\].stg01
timestamp 1698431365
transform 1 0 25484 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[1\].stg02
timestamp 1698431365
transform 1 0 24656 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[2\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 20056 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[2\].stg01
timestamp 1698431365
transform -1 0 20976 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[2\].stg02
timestamp 1698431365
transform 1 0 20516 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[3\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 21160 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[3\].stg01
timestamp 1698431365
transform 1 0 20332 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[3\].stg02
timestamp 1698431365
transform 1 0 20056 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[4\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 15640 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[4\].stg01
timestamp 1698431365
transform 1 0 20240 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[4\].stg02
timestamp 1698431365
transform 1 0 19596 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[5\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 19320 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[5\].stg01
timestamp 1698431365
transform 1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[5\].stg02
timestamp 1698431365
transform 1 0 19044 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[6\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 19136 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[6\].stg01
timestamp 1698431365
transform 1 0 18124 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[6\].stg02
timestamp 1698431365
transform 1 0 17664 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[7\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 16928 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[7\].stg01
timestamp 1698431365
transform 1 0 18400 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[7\].stg02
timestamp 1698431365
transform -1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[8\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 20332 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[8\].stg01
timestamp 1698431365
transform -1 0 19412 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[8\].stg02
timestamp 1698431365
transform -1 0 19780 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[9\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 20976 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[9\].stg01
timestamp 1698431365
transform -1 0 20424 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[9\].stg02
timestamp 1698431365
transform -1 0 20976 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[10\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 23000 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[10\].stg01
timestamp 1698431365
transform -1 0 21160 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[10\].stg02
timestamp 1698431365
transform -1 0 22816 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[11\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 28060 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[11\].stg01
timestamp 1698431365
transform -1 0 27048 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[11\].stg02
timestamp 1698431365
transform -1 0 27692 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[12\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 28520 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[12\].stg01
timestamp 1698431365
transform 1 0 29532 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[12\].stg02
timestamp 1698431365
transform 1 0 28980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[13\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 29624 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[13\].stg01
timestamp 1698431365
transform -1 0 29256 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[13\].stg02
timestamp 1698431365
transform -1 0 29348 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[14\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 29992 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[14\].stg01
timestamp 1698431365
transform 1 0 28980 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[14\].stg02
timestamp 1698431365
transform -1 0 29348 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[15\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 29716 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[15\].stg01
timestamp 1698431365
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[15\].stg02
timestamp 1698431365
transform 1 0 28428 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring1\[16\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 26036 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring1\[16\].stg01
timestamp 1698431365
transform 1 0 27600 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring1\[16\].stg02_62
timestamp 1698431365
transform 1 0 25576 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring1\[16\].stg02
timestamp 1698431365
transform 1 0 27140 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[16\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 26036 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[16\].stg01_63
timestamp 1698431365
transform -1 0 29532 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[16\].stg01
timestamp 1698431365
transform -1 0 26956 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[16\].stg02
timestamp 1698431365
transform -1 0 27140 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[17\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 22172 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[17\].stg01_64
timestamp 1698431365
transform -1 0 25484 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[17\].stg01
timestamp 1698431365
transform 1 0 25116 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[17\].stg02
timestamp 1698431365
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[18\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 21896 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[18\].stg01_65
timestamp 1698431365
transform 1 0 21252 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[18\].stg01
timestamp 1698431365
transform 1 0 21896 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[18\].stg02
timestamp 1698431365
transform 1 0 21252 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[19\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 20240 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[19\].stg01
timestamp 1698431365
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[19\].stg01_66
timestamp 1698431365
transform 1 0 20240 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[19\].stg02
timestamp 1698431365
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[20\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 18308 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[20\].stg01_67
timestamp 1698431365
transform -1 0 20792 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[20\].stg01
timestamp 1698431365
transform -1 0 20240 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[20\].stg02
timestamp 1698431365
transform 1 0 19228 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[21\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 19320 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[21\].stg01_68
timestamp 1698431365
transform 1 0 18676 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[21\].stg01
timestamp 1698431365
transform -1 0 18952 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[21\].stg02
timestamp 1698431365
transform -1 0 19044 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[22\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 17572 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[22\].stg01_69
timestamp 1698431365
transform -1 0 18952 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[22\].stg01
timestamp 1698431365
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[22\].stg02
timestamp 1698431365
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[23\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 22172 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[23\].stg01_70
timestamp 1698431365
transform -1 0 18400 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[23\].stg01
timestamp 1698431365
transform -1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[23\].stg02
timestamp 1698431365
transform 1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[24\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 19228 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[24\].stg01_71
timestamp 1698431365
transform 1 0 19780 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[24\].stg01
timestamp 1698431365
transform 1 0 20424 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[24\].stg02
timestamp 1698431365
transform 1 0 19780 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[25\].g_buf2.ctr_buf
timestamp 1698431365
transform 1 0 23184 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[25\].stg01
timestamp 1698431365
transform -1 0 19872 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[25\].stg01_72
timestamp 1698431365
transform -1 0 20240 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[25\].stg02
timestamp 1698431365
transform -1 0 20608 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[26\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 23920 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[26\].stg01_73
timestamp 1698431365
transform -1 0 23000 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[26\].stg01
timestamp 1698431365
transform -1 0 22448 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[26\].stg02
timestamp 1698431365
transform -1 0 23184 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[27\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 27232 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[27\].stg01_74
timestamp 1698431365
transform 1 0 26404 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[27\].stg01
timestamp 1698431365
transform -1 0 26956 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[27\].stg02
timestamp 1698431365
transform -1 0 27324 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[28\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 29992 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[28\].stg01
timestamp 1698431365
transform 1 0 29256 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[28\].stg01_75
timestamp 1698431365
transform 1 0 28612 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[28\].stg02
timestamp 1698431365
transform 1 0 28888 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[29\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 30544 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[29\].stg01
timestamp 1698431365
transform -1 0 29624 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[29\].stg01_76
timestamp 1698431365
transform -1 0 29716 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[29\].stg02
timestamp 1698431365
transform 1 0 28520 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[30\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 29992 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[30\].stg01_77
timestamp 1698431365
transform -1 0 30268 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[30\].stg01
timestamp 1698431365
transform -1 0 28980 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[30\].stg02
timestamp 1698431365
transform -1 0 29716 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  tdc1.g_ring3\[31\].g_buf2.ctr_buf
timestamp 1698431365
transform -1 0 27232 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.g_ring3\[31\].stg01_78
timestamp 1698431365
transform -1 0 29716 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  tdc1.g_ring3\[31\].stg01
timestamp 1698431365
transform 1 0 28612 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.g_ring3\[31\].stg02
timestamp 1698431365
transform 1 0 28060 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  tdc1.stg01
timestamp 1698431365
transform 1 0 27508 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tdc1.stg01_79
timestamp 1698431365
transform 1 0 27232 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  tdc1.stg02
timestamp 1698431365
transform 1 0 26404 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_80
timestamp 1698431365
transform -1 0 6256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_81
timestamp 1698431365
transform -1 0 5520 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_82
timestamp 1698431365
transform -1 0 4784 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_83
timestamp 1698431365
transform -1 0 4048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_84
timestamp 1698431365
transform -1 0 3496 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_85
timestamp 1698431365
transform -1 0 2576 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_86
timestamp 1698431365
transform -1 0 1840 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_87
timestamp 1698431365
transform -1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_88
timestamp 1698431365
transform -1 0 12144 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_89
timestamp 1698431365
transform -1 0 11408 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_90
timestamp 1698431365
transform -1 0 10672 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_91
timestamp 1698431365
transform -1 0 9936 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_92
timestamp 1698431365
transform 1 0 8556 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_93
timestamp 1698431365
transform 1 0 8004 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_94
timestamp 1698431365
transform -1 0 7728 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_hpretl_tt06_tdc_v2_95
timestamp 1698431365
transform -1 0 6992 0 1 21216
box -38 -48 314 592
<< labels >>
flabel metal4 s 8166 496 8486 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15940 496 16260 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23714 496 24034 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31488 496 31808 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4279 496 4599 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12053 496 12373 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19827 496 20147 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27601 496 27921 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 30974 22104 31034 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 31710 22104 31770 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 30238 22104 30298 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 29502 22104 29562 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 28030 22104 28090 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 27294 22104 27354 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 25086 22104 25146 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 22878 22104 22938 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 20670 22104 20730 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 18462 22104 18522 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal4 s 5214 22104 5274 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal4 s 4478 22104 4538 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal4 s 3742 22104 3802 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal4 s 3006 22104 3066 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal4 s 2270 22104 2330 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal4 s 1534 22104 1594 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal4 s 798 22104 858 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal4 s 11838 22104 11898 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal4 s 9630 22104 9690 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal4 s 7422 22104 7482 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal4 s 16254 22104 16314 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal4 s 14046 22104 14106 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 16180 21216 16180 21216 0 VGND
rlabel metal1 16100 21760 16100 21760 0 VPWR
rlabel metal1 11776 9690 11776 9690 0 _000_
rlabel metal1 1242 12886 1242 12886 0 _001_
rlabel metal1 3772 13430 3772 13430 0 _002_
rlabel metal2 1426 14212 1426 14212 0 _003_
rlabel metal1 3542 14586 3542 14586 0 _004_
rlabel metal1 1380 15946 1380 15946 0 _005_
rlabel metal1 1564 16694 1564 16694 0 _006_
rlabel metal1 14030 9690 14030 9690 0 _007_
rlabel metal2 14122 10880 14122 10880 0 _008_
rlabel metal1 11546 10778 11546 10778 0 _009_
rlabel metal1 9522 10642 9522 10642 0 _010_
rlabel metal1 8740 11594 8740 11594 0 _011_
rlabel metal2 7774 10812 7774 10812 0 _012_
rlabel metal1 5980 11254 5980 11254 0 _013_
rlabel metal1 3358 11050 3358 11050 0 _014_
rlabel metal1 3450 12410 3450 12410 0 _015_
rlabel metal1 27048 11594 27048 11594 0 _016_
rlabel metal1 21850 10642 21850 10642 0 _017_
rlabel metal1 19274 10642 19274 10642 0 _018_
rlabel metal1 16744 10030 16744 10030 0 _019_
rlabel metal1 17296 11322 17296 11322 0 _020_
rlabel metal1 18078 12886 18078 12886 0 _021_
rlabel metal1 20286 12818 20286 12818 0 _022_
rlabel metal1 28980 12138 28980 12138 0 _023_
rlabel metal2 29486 13634 29486 13634 0 _024_
rlabel metal1 29072 12682 29072 12682 0 _025_
rlabel metal1 27508 14246 27508 14246 0 _026_
rlabel metal1 25300 13498 25300 13498 0 _027_
rlabel metal1 27554 12206 27554 12206 0 _028_
rlabel metal1 24564 11866 24564 11866 0 _029_
rlabel metal1 24104 10030 24104 10030 0 _030_
rlabel metal1 26910 11084 26910 11084 0 _031_
rlabel metal2 12558 9894 12558 9894 0 _032_
rlabel metal1 15417 10166 15417 10166 0 _033_
rlabel metal2 14858 11016 14858 11016 0 _034_
rlabel metal2 12466 11016 12466 11016 0 _035_
rlabel metal1 10488 10234 10488 10234 0 _036_
rlabel metal1 10403 11594 10403 11594 0 _037_
rlabel metal1 8241 10506 8241 10506 0 _038_
rlabel metal2 7130 11016 7130 11016 0 _039_
rlabel metal1 5113 11254 5113 11254 0 _040_
rlabel metal1 4692 11866 4692 11866 0 _041_
rlabel metal1 2859 13430 2859 13430 0 _042_
rlabel metal1 4600 12954 4600 12954 0 _043_
rlabel metal1 2905 14518 2905 14518 0 _044_
rlabel metal1 4416 14586 4416 14586 0 _045_
rlabel metal2 2622 16184 2622 16184 0 _046_
rlabel metal1 2300 16762 2300 16762 0 _047_
rlabel metal2 28566 11458 28566 11458 0 _048_
rlabel metal1 30084 11866 30084 11866 0 _049_
rlabel metal1 30268 13498 30268 13498 0 _050_
rlabel metal1 30827 12682 30827 12682 0 _051_
rlabel metal1 28106 13498 28106 13498 0 _052_
rlabel metal2 25622 13634 25622 13634 0 _053_
rlabel metal2 26910 12381 26910 12381 0 _054_
rlabel metal1 25576 11866 25576 11866 0 _055_
rlabel metal1 25721 10506 25721 10506 0 _056_
rlabel metal2 27462 11016 27462 11016 0 _057_
rlabel metal1 23000 10234 23000 10234 0 _058_
rlabel metal2 19826 10370 19826 10370 0 _059_
rlabel metal1 18177 10506 18177 10506 0 _060_
rlabel metal1 18545 11594 18545 11594 0 _061_
rlabel metal1 16928 12410 16928 12410 0 _062_
rlabel metal1 21429 12750 21429 12750 0 _063_
rlabel metal1 27646 17578 27646 17578 0 _064_
rlabel metal1 27554 18938 27554 18938 0 _065_
rlabel via1 25251 16626 25251 16626 0 _066_
rlabel metal1 25024 17646 25024 17646 0 _067_
rlabel metal1 15042 16626 15042 16626 0 _068_
rlabel metal1 21896 16626 21896 16626 0 _069_
rlabel metal1 15962 16218 15962 16218 0 _070_
rlabel metal1 23230 15606 23230 15606 0 _071_
rlabel metal2 16514 19635 16514 19635 0 _072_
rlabel metal1 15686 16456 15686 16456 0 _073_
rlabel metal1 27232 18190 27232 18190 0 _074_
rlabel metal1 16790 20570 16790 20570 0 _075_
rlabel via1 15778 19346 15778 19346 0 _076_
rlabel metal2 16790 16456 16790 16456 0 _077_
rlabel metal1 16836 16762 16836 16762 0 _078_
rlabel metal1 21528 14926 21528 14926 0 _079_
rlabel metal1 22540 14450 22540 14450 0 _080_
rlabel metal1 22954 16116 22954 16116 0 _081_
rlabel metal1 22356 16218 22356 16218 0 _082_
rlabel metal1 15870 20026 15870 20026 0 _083_
rlabel metal3 24472 16524 24472 16524 0 _084_
rlabel metal1 22218 20400 22218 20400 0 _085_
rlabel metal2 22862 17272 22862 17272 0 _086_
rlabel metal1 21482 15572 21482 15572 0 _087_
rlabel metal1 21574 15674 21574 15674 0 _088_
rlabel metal1 21896 20366 21896 20366 0 _089_
rlabel metal1 20102 20502 20102 20502 0 _090_
rlabel metal1 17802 20434 17802 20434 0 _091_
rlabel metal1 15318 14994 15318 14994 0 _092_
rlabel metal2 15226 15266 15226 15266 0 _093_
rlabel metal1 14720 14586 14720 14586 0 _094_
rlabel metal1 16008 15130 16008 15130 0 _095_
rlabel metal1 24242 16660 24242 16660 0 _096_
rlabel metal2 24242 18054 24242 18054 0 _097_
rlabel metal1 24426 16626 24426 16626 0 _098_
rlabel metal1 19918 17170 19918 17170 0 _099_
rlabel metal1 17204 17102 17204 17102 0 _100_
rlabel metal1 13938 14586 13938 14586 0 _101_
rlabel metal1 15180 15062 15180 15062 0 _102_
rlabel metal1 15226 15946 15226 15946 0 _103_
rlabel metal1 23138 16660 23138 16660 0 _104_
rlabel metal1 22540 15538 22540 15538 0 _105_
rlabel metal1 22264 15334 22264 15334 0 _106_
rlabel metal1 22218 14586 22218 14586 0 _107_
rlabel metal1 21022 15538 21022 15538 0 _108_
rlabel metal1 18032 16218 18032 16218 0 _109_
rlabel metal2 21574 16252 21574 16252 0 _110_
rlabel metal1 17756 16490 17756 16490 0 _111_
rlabel metal1 14030 17068 14030 17068 0 _112_
rlabel metal1 13754 16762 13754 16762 0 _113_
rlabel metal1 13386 17306 13386 17306 0 _114_
rlabel metal1 13432 17714 13432 17714 0 _115_
rlabel metal1 13846 17204 13846 17204 0 _116_
rlabel metal1 14398 17204 14398 17204 0 _117_
rlabel metal1 12696 16014 12696 16014 0 _118_
rlabel metal1 13800 16218 13800 16218 0 _119_
rlabel metal1 14214 18666 14214 18666 0 _120_
rlabel metal1 27140 18394 27140 18394 0 _121_
rlabel metal1 27186 18258 27186 18258 0 _122_
rlabel metal1 27094 17850 27094 17850 0 _123_
rlabel metal1 23598 18394 23598 18394 0 _124_
rlabel metal2 20838 17204 20838 17204 0 _125_
rlabel metal1 19274 18326 19274 18326 0 _126_
rlabel metal2 13570 20706 13570 20706 0 _127_
rlabel metal2 12834 20672 12834 20672 0 _128_
rlabel metal2 13478 15827 13478 15827 0 _129_
rlabel metal1 12834 15402 12834 15402 0 _130_
rlabel metal1 14306 21012 14306 21012 0 _131_
rlabel metal1 18446 20570 18446 20570 0 _132_
rlabel metal2 18722 15946 18722 15946 0 _133_
rlabel metal1 18216 15062 18216 15062 0 _134_
rlabel metal1 13984 19482 13984 19482 0 _135_
rlabel metal1 13570 17578 13570 17578 0 _136_
rlabel metal1 13886 19890 13886 19890 0 _137_
rlabel metal1 14720 20026 14720 20026 0 _138_
rlabel metal1 25024 20570 25024 20570 0 _139_
rlabel metal2 24702 19992 24702 19992 0 _140_
rlabel metal2 24426 15759 24426 15759 0 _141_
rlabel metal2 15318 20417 15318 20417 0 _142_
rlabel metal1 14904 20366 14904 20366 0 _143_
rlabel metal1 13892 10574 13892 10574 0 _144_
rlabel metal1 13662 11050 13662 11050 0 _145_
rlabel metal1 12742 11594 12742 11594 0 _146_
rlabel metal1 5842 12206 5842 12206 0 _147_
rlabel metal1 11638 10540 11638 10540 0 _148_
rlabel metal1 5474 12104 5474 12104 0 _149_
rlabel metal1 8096 11594 8096 11594 0 _150_
rlabel metal1 8782 11322 8782 11322 0 _151_
rlabel metal2 6578 11322 6578 11322 0 _152_
rlabel metal1 7636 11186 7636 11186 0 _153_
rlabel metal1 5530 12342 5530 12342 0 _154_
rlabel metal1 6118 12342 6118 12342 0 _155_
rlabel metal1 2346 12206 2346 12206 0 _156_
rlabel metal1 2576 12206 2576 12206 0 _157_
rlabel metal1 1518 12852 1518 12852 0 _158_
rlabel metal1 4094 12954 4094 12954 0 _159_
rlabel metal1 5934 12750 5934 12750 0 _160_
rlabel metal1 4002 13872 4002 13872 0 _161_
rlabel metal1 3910 15572 3910 15572 0 _162_
rlabel metal1 3818 14484 3818 14484 0 _163_
rlabel metal1 3542 14450 3542 14450 0 _164_
rlabel metal1 1058 15946 1058 15946 0 _165_
rlabel metal1 1978 15674 1978 15674 0 _166_
rlabel metal1 29578 13328 29578 13328 0 _167_
rlabel metal1 29118 13396 29118 13396 0 _168_
rlabel metal1 29532 14450 29532 14450 0 _169_
rlabel metal2 28658 13498 28658 13498 0 _170_
rlabel metal1 28842 12784 28842 12784 0 _171_
rlabel metal1 23046 12648 23046 12648 0 _172_
rlabel metal1 25438 13396 25438 13396 0 _173_
rlabel metal1 25162 13362 25162 13362 0 _174_
rlabel metal1 25346 12716 25346 12716 0 _175_
rlabel metal1 25530 12784 25530 12784 0 _176_
rlabel metal1 23138 12750 23138 12750 0 _177_
rlabel metal1 22954 12342 22954 12342 0 _178_
rlabel metal1 24702 11696 24702 11696 0 _179_
rlabel metal1 25530 11118 25530 11118 0 _180_
rlabel metal1 21252 10234 21252 10234 0 _181_
rlabel metal1 20792 11050 20792 11050 0 _182_
rlabel metal1 22448 11186 22448 11186 0 _183_
rlabel metal1 20102 11220 20102 11220 0 _184_
rlabel metal1 18262 12614 18262 12614 0 _185_
rlabel metal1 18032 11050 18032 11050 0 _186_
rlabel metal1 17710 11254 17710 11254 0 _187_
rlabel metal1 18998 12750 18998 12750 0 _188_
rlabel metal1 18216 12410 18216 12410 0 _189_
rlabel metal1 13294 14586 13294 14586 0 _190_
rlabel metal1 14720 14790 14720 14790 0 _191_
rlabel metal1 17756 15130 17756 15130 0 _192_
rlabel metal1 21482 14042 21482 14042 0 _193_
rlabel metal1 21482 14450 21482 14450 0 _194_
rlabel metal1 21712 14382 21712 14382 0 _195_
rlabel metal1 21022 14586 21022 14586 0 _196_
rlabel metal1 6118 10540 6118 10540 0 _197_
rlabel metal1 25668 11662 25668 11662 0 _198_
rlabel metal1 29026 21386 29026 21386 0 net1
rlabel metal1 24150 10642 24150 10642 0 net10
rlabel metal1 14214 14008 14214 14008 0 net11
rlabel metal1 11546 17680 11546 17680 0 net12
rlabel metal2 5290 19176 5290 19176 0 net13
rlabel metal1 17296 19890 17296 19890 0 net14
rlabel metal2 20424 19890 20424 19890 0 net15
rlabel metal1 21482 13396 21482 13396 0 net16
rlabel metal1 27140 20978 27140 20978 0 net17
rlabel metal1 27462 17170 27462 17170 0 net18
rlabel metal1 2668 18802 2668 18802 0 net19
rlabel metal1 29578 21080 29578 21080 0 net2
rlabel metal1 2714 16660 2714 16660 0 net20
rlabel metal1 10810 17714 10810 17714 0 net21
rlabel via1 7406 16626 7406 16626 0 net22
rlabel metal1 10718 13872 10718 13872 0 net23
rlabel metal1 17388 20298 17388 20298 0 net24
rlabel metal1 19734 16456 19734 16456 0 net25
rlabel metal1 4186 16014 4186 16014 0 net26
rlabel metal2 8786 21114 8786 21114 0 net27
rlabel metal1 9200 21454 9200 21454 0 net28
rlabel metal1 14628 12274 14628 12274 0 net29
rlabel metal2 13202 19822 13202 19822 0 net3
rlabel metal1 16192 14450 16192 14450 0 net30
rlabel metal1 10948 17102 10948 17102 0 net31
rlabel metal1 15962 15470 15962 15470 0 net32
rlabel metal1 22402 11832 22402 11832 0 net33
rlabel metal1 17710 19788 17710 19788 0 net34
rlabel metal1 23506 21420 23506 21420 0 net35
rlabel metal1 26082 15538 26082 15538 0 net36
rlabel metal1 28704 19686 28704 19686 0 net37
rlabel metal1 16100 21454 16100 21454 0 net38
rlabel metal1 5474 19958 5474 19958 0 net39
rlabel metal1 27324 19278 27324 19278 0 net4
rlabel metal1 5290 18326 5290 18326 0 net40
rlabel metal1 27002 17136 27002 17136 0 net41
rlabel metal2 29026 18734 29026 18734 0 net42
rlabel metal1 10304 17714 10304 17714 0 net43
rlabel metal1 3956 18666 3956 18666 0 net44
rlabel metal1 4002 19244 4002 19244 0 net45
rlabel metal1 4416 17714 4416 17714 0 net46
rlabel metal1 5980 17714 5980 17714 0 net47
rlabel metal1 10810 16626 10810 16626 0 net48
rlabel metal1 9200 17714 9200 17714 0 net49
rlabel metal1 25990 19924 25990 19924 0 net5
rlabel metal2 9246 18819 9246 18819 0 net50
rlabel metal1 8970 19244 8970 19244 0 net51
rlabel metal1 9660 20366 9660 20366 0 net52
rlabel metal1 10810 18768 10810 18768 0 net53
rlabel metal1 10120 13838 10120 13838 0 net54
rlabel metal1 9798 13906 9798 13906 0 net55
rlabel metal1 8096 14042 8096 14042 0 net56
rlabel metal1 7544 15538 7544 15538 0 net57
rlabel metal1 6854 17136 6854 17136 0 net58
rlabel metal1 6256 18190 6256 18190 0 net59
rlabel metal1 26128 19890 26128 19890 0 net6
rlabel metal1 6256 19278 6256 19278 0 net60
rlabel metal1 3864 19414 3864 19414 0 net61
rlabel metal2 27278 21182 27278 21182 0 net62
rlabel metal2 26910 20944 26910 20944 0 net63
rlabel metal1 25208 20978 25208 20978 0 net64
rlabel metal1 21942 21012 21942 21012 0 net65
rlabel metal1 20562 20910 20562 20910 0 net66
rlabel metal1 20562 17748 20562 17748 0 net67
rlabel metal2 18906 18156 18906 18156 0 net68
rlabel metal1 18492 18802 18492 18802 0 net69
rlabel metal2 1242 17306 1242 17306 0 net7
rlabel metal1 17618 19244 17618 19244 0 net70
rlabel metal1 20516 19278 20516 19278 0 net71
rlabel metal1 19872 18394 19872 18394 0 net72
rlabel metal1 22494 18190 22494 18190 0 net73
rlabel metal1 26634 16660 26634 16660 0 net74
rlabel metal1 28934 16558 28934 16558 0 net75
rlabel metal1 29532 17306 29532 17306 0 net76
rlabel metal2 28934 19091 28934 19091 0 net77
rlabel metal1 29072 19822 29072 19822 0 net78
rlabel metal1 27508 20570 27508 20570 0 net79
rlabel metal1 11270 10166 11270 10166 0 net8
rlabel metal2 6026 21743 6026 21743 0 net80
rlabel metal2 5290 21743 5290 21743 0 net81
rlabel metal1 4600 21658 4600 21658 0 net82
rlabel metal2 3818 21743 3818 21743 0 net83
rlabel metal2 3266 21743 3266 21743 0 net84
rlabel metal2 2346 21743 2346 21743 0 net85
rlabel metal2 1610 21743 1610 21743 0 net86
rlabel metal2 874 21743 874 21743 0 net87
rlabel metal2 11914 21267 11914 21267 0 net88
rlabel metal2 11178 21743 11178 21743 0 net89
rlabel metal1 26910 11730 26910 11730 0 net9
rlabel metal2 10442 21743 10442 21743 0 net90
rlabel metal2 9706 21743 9706 21743 0 net91
rlabel metal2 8786 21743 8786 21743 0 net92
rlabel metal2 8234 21811 8234 21811 0 net93
rlabel metal2 7498 21743 7498 21743 0 net94
rlabel metal2 6762 21743 6762 21743 0 net95
rlabel metal1 13662 12954 13662 12954 0 tdc0.r_dly_store_ctr\[0\]
rlabel metal2 13754 14620 13754 14620 0 tdc0.r_dly_store_ctr\[10\]
rlabel via2 7222 14331 7222 14331 0 tdc0.r_dly_store_ctr\[11\]
rlabel metal1 13570 16660 13570 16660 0 tdc0.r_dly_store_ctr\[12\]
rlabel metal1 10902 15946 10902 15946 0 tdc0.r_dly_store_ctr\[13\]
rlabel metal2 13294 15980 13294 15980 0 tdc0.r_dly_store_ctr\[14\]
rlabel metal1 4876 17238 4876 17238 0 tdc0.r_dly_store_ctr\[15\]
rlabel metal1 16192 12410 16192 12410 0 tdc0.r_dly_store_ctr\[1\]
rlabel metal1 14076 13498 14076 13498 0 tdc0.r_dly_store_ctr\[2\]
rlabel metal1 14628 12410 14628 12410 0 tdc0.r_dly_store_ctr\[3\]
rlabel metal1 13018 17136 13018 17136 0 tdc0.r_dly_store_ctr\[4\]
rlabel metal1 12742 12410 12742 12410 0 tdc0.r_dly_store_ctr\[5\]
rlabel metal1 10948 12614 10948 12614 0 tdc0.r_dly_store_ctr\[6\]
rlabel metal2 12926 15300 12926 15300 0 tdc0.r_dly_store_ctr\[7\]
rlabel metal2 12466 13838 12466 13838 0 tdc0.r_dly_store_ctr\[8\]
rlabel metal2 13018 14858 13018 14858 0 tdc0.r_dly_store_ctr\[9\]
rlabel viali 17158 14926 17158 14926 0 tdc0.r_dly_store_ring\[0\]
rlabel metal1 11500 15130 11500 15130 0 tdc0.r_dly_store_ring\[10\]
rlabel metal2 14214 15810 14214 15810 0 tdc0.r_dly_store_ring\[11\]
rlabel metal2 12834 18326 12834 18326 0 tdc0.r_dly_store_ring\[12\]
rlabel metal1 13846 18734 13846 18734 0 tdc0.r_dly_store_ring\[13\]
rlabel metal1 13846 20332 13846 20332 0 tdc0.r_dly_store_ring\[14\]
rlabel metal1 6348 19142 6348 19142 0 tdc0.r_dly_store_ring\[15\]
rlabel via2 13662 14909 13662 14909 0 tdc0.r_dly_store_ring\[16\]
rlabel metal1 11250 16592 11250 16592 0 tdc0.r_dly_store_ring\[17\]
rlabel metal2 14306 16116 14306 16116 0 tdc0.r_dly_store_ring\[18\]
rlabel metal1 14491 14892 14491 14892 0 tdc0.r_dly_store_ring\[19\]
rlabel metal1 16652 20366 16652 20366 0 tdc0.r_dly_store_ring\[1\]
rlabel metal2 13110 18598 13110 18598 0 tdc0.r_dly_store_ring\[20\]
rlabel metal1 12834 16116 12834 16116 0 tdc0.r_dly_store_ring\[21\]
rlabel metal1 12811 20434 12811 20434 0 tdc0.r_dly_store_ring\[22\]
rlabel metal1 13156 19346 13156 19346 0 tdc0.r_dly_store_ring\[23\]
rlabel metal2 12742 14246 12742 14246 0 tdc0.r_dly_store_ring\[24\]
rlabel metal1 16698 15980 16698 15980 0 tdc0.r_dly_store_ring\[25\]
rlabel metal2 13846 15334 13846 15334 0 tdc0.r_dly_store_ring\[26\]
rlabel metal1 8970 14552 8970 14552 0 tdc0.r_dly_store_ring\[27\]
rlabel metal1 11086 17136 11086 17136 0 tdc0.r_dly_store_ring\[28\]
rlabel metal1 7958 16048 7958 16048 0 tdc0.r_dly_store_ring\[29\]
rlabel metal1 15916 19142 15916 19142 0 tdc0.r_dly_store_ring\[2\]
rlabel via2 19550 18683 19550 18683 0 tdc0.r_dly_store_ring\[30\]
rlabel metal1 7958 19992 7958 19992 0 tdc0.r_dly_store_ring\[31\]
rlabel metal1 13294 15912 13294 15912 0 tdc0.r_dly_store_ring\[3\]
rlabel metal1 14858 17850 14858 17850 0 tdc0.r_dly_store_ring\[4\]
rlabel metal1 13202 19142 13202 19142 0 tdc0.r_dly_store_ring\[5\]
rlabel metal1 12489 21114 12489 21114 0 tdc0.r_dly_store_ring\[6\]
rlabel metal1 13800 21454 13800 21454 0 tdc0.r_dly_store_ring\[7\]
rlabel metal1 17480 14586 17480 14586 0 tdc0.r_dly_store_ring\[8\]
rlabel metal1 16606 14042 16606 14042 0 tdc0.r_dly_store_ring\[9\]
rlabel metal1 12098 9520 12098 9520 0 tdc0.r_ring_ctr\[0\]
rlabel metal1 6026 13362 6026 13362 0 tdc0.r_ring_ctr\[10\]
rlabel metal1 6072 13498 6072 13498 0 tdc0.r_ring_ctr\[11\]
rlabel metal1 1978 14246 1978 14246 0 tdc0.r_ring_ctr\[12\]
rlabel metal2 5106 15538 5106 15538 0 tdc0.r_ring_ctr\[13\]
rlabel metal1 2162 15572 2162 15572 0 tdc0.r_ring_ctr\[14\]
rlabel metal2 1426 16796 1426 16796 0 tdc0.r_ring_ctr\[15\]
rlabel metal1 14674 11798 14674 11798 0 tdc0.r_ring_ctr\[1\]
rlabel metal1 13197 13362 13197 13362 0 tdc0.r_ring_ctr\[2\]
rlabel metal2 13754 11934 13754 11934 0 tdc0.r_ring_ctr\[3\]
rlabel metal1 8970 10506 8970 10506 0 tdc0.r_ring_ctr\[4\]
rlabel metal2 10442 12070 10442 12070 0 tdc0.r_ring_ctr\[5\]
rlabel metal2 7498 11713 7498 11713 0 tdc0.r_ring_ctr\[6\]
rlabel metal1 6486 11696 6486 11696 0 tdc0.r_ring_ctr\[7\]
rlabel metal1 5704 11322 5704 11322 0 tdc0.r_ring_ctr\[8\]
rlabel metal1 5290 12410 5290 12410 0 tdc0.r_ring_ctr\[9\]
rlabel metal1 3128 19482 3128 19482 0 tdc0.w_dly_stop\[1\]
rlabel metal2 3726 19482 3726 19482 0 tdc0.w_dly_stop\[2\]
rlabel metal1 3450 19482 3450 19482 0 tdc0.w_dly_stop\[3\]
rlabel metal1 3588 19890 3588 19890 0 tdc0.w_dly_stop\[4\]
rlabel metal1 4876 18802 4876 18802 0 tdc0.w_dly_stop\[5\]
rlabel metal1 5520 17510 5520 17510 0 tdc0.w_ring_buf\[0\]
rlabel metal1 9506 14858 9506 14858 0 tdc0.w_ring_buf\[10\]
rlabel metal1 8218 15606 8218 15606 0 tdc0.w_ring_buf\[11\]
rlabel via1 7769 17782 7769 17782 0 tdc0.w_ring_buf\[12\]
rlabel metal1 7252 18870 7252 18870 0 tdc0.w_ring_buf\[13\]
rlabel metal2 6486 20162 6486 20162 0 tdc0.w_ring_buf\[14\]
rlabel via1 5193 19278 5193 19278 0 tdc0.w_ring_buf\[15\]
rlabel metal1 5428 15334 5428 15334 0 tdc0.w_ring_buf\[16\]
rlabel metal1 5182 17034 5182 17034 0 tdc0.w_ring_buf\[17\]
rlabel metal1 11070 17034 11070 17034 0 tdc0.w_ring_buf\[18\]
rlabel metal1 10978 15606 10978 15606 0 tdc0.w_ring_buf\[19\]
rlabel metal1 15497 21046 15497 21046 0 tdc0.w_ring_buf\[1\]
rlabel metal1 11076 18190 11076 18190 0 tdc0.w_ring_buf\[20\]
rlabel via1 9057 16014 9057 16014 0 tdc0.w_ring_buf\[21\]
rlabel via1 10253 20366 10253 20366 0 tdc0.w_ring_buf\[22\]
rlabel metal1 11438 19958 11438 19958 0 tdc0.w_ring_buf\[23\]
rlabel metal1 11536 13838 11536 13838 0 tdc0.w_ring_buf\[24\]
rlabel metal1 13439 13430 13439 13430 0 tdc0.w_ring_buf\[25\]
rlabel metal1 9844 14586 9844 14586 0 tdc0.w_ring_buf\[26\]
rlabel metal1 7666 14518 7666 14518 0 tdc0.w_ring_buf\[27\]
rlabel metal1 8218 17034 8218 17034 0 tdc0.w_ring_buf\[28\]
rlabel metal1 6987 16014 6987 16014 0 tdc0.w_ring_buf\[29\]
rlabel metal1 12558 18938 12558 18938 0 tdc0.w_ring_buf\[2\]
rlabel via2 15226 18853 15226 18853 0 tdc0.w_ring_buf\[30\]
rlabel metal1 6516 19958 6516 19958 0 tdc0.w_ring_buf\[31\]
rlabel metal1 10432 16014 10432 16014 0 tdc0.w_ring_buf\[3\]
rlabel metal1 13186 18122 13186 18122 0 tdc0.w_ring_buf\[4\]
rlabel metal1 11116 19142 11116 19142 0 tdc0.w_ring_buf\[5\]
rlabel metal2 8878 20774 8878 20774 0 tdc0.w_ring_buf\[6\]
rlabel metal2 11454 21250 11454 21250 0 tdc0.w_ring_buf\[7\]
rlabel metal1 16268 14518 16268 14518 0 tdc0.w_ring_buf\[8\]
rlabel metal1 14848 13838 14848 13838 0 tdc0.w_ring_buf\[9\]
rlabel metal1 4646 18870 4646 18870 0 tdc0.w_ring_int_norsz\[0\]
rlabel metal1 10396 14382 10396 14382 0 tdc0.w_ring_int_norsz\[10\]
rlabel metal1 8372 14994 8372 14994 0 tdc0.w_ring_int_norsz\[11\]
rlabel metal1 7958 16218 7958 16218 0 tdc0.w_ring_int_norsz\[12\]
rlabel metal1 6716 17782 6716 17782 0 tdc0.w_ring_int_norsz\[13\]
rlabel metal1 6532 18938 6532 18938 0 tdc0.w_ring_int_norsz\[14\]
rlabel metal1 6532 19482 6532 19482 0 tdc0.w_ring_int_norsz\[15\]
rlabel metal1 4324 19482 4324 19482 0 tdc0.w_ring_int_norsz\[16\]
rlabel metal1 4830 17646 4830 17646 0 tdc0.w_ring_int_norsz\[17\]
rlabel metal1 9430 17646 9430 17646 0 tdc0.w_ring_int_norsz\[18\]
rlabel metal1 10580 16762 10580 16762 0 tdc0.w_ring_int_norsz\[19\]
rlabel metal1 4830 17816 4830 17816 0 tdc0.w_ring_int_norsz\[1\]
rlabel metal1 9752 17782 9752 17782 0 tdc0.w_ring_int_norsz\[20\]
rlabel metal2 9706 19040 9706 19040 0 tdc0.w_ring_int_norsz\[21\]
rlabel metal1 8832 19482 8832 19482 0 tdc0.w_ring_int_norsz\[22\]
rlabel metal1 9706 19958 9706 19958 0 tdc0.w_ring_int_norsz\[23\]
rlabel metal1 10856 18938 10856 18938 0 tdc0.w_ring_int_norsz\[24\]
rlabel metal1 10350 13906 10350 13906 0 tdc0.w_ring_int_norsz\[25\]
rlabel metal2 9798 14212 9798 14212 0 tdc0.w_ring_int_norsz\[26\]
rlabel metal1 8050 14858 8050 14858 0 tdc0.w_ring_int_norsz\[27\]
rlabel metal1 7452 15674 7452 15674 0 tdc0.w_ring_int_norsz\[28\]
rlabel metal1 6808 17306 6808 17306 0 tdc0.w_ring_int_norsz\[29\]
rlabel metal1 11362 17646 11362 17646 0 tdc0.w_ring_int_norsz\[2\]
rlabel metal1 6348 18054 6348 18054 0 tdc0.w_ring_int_norsz\[30\]
rlabel metal2 5658 18921 5658 18921 0 tdc0.w_ring_int_norsz\[31\]
rlabel metal1 10626 17204 10626 17204 0 tdc0.w_ring_int_norsz\[3\]
rlabel metal1 9706 17850 9706 17850 0 tdc0.w_ring_int_norsz\[4\]
rlabel metal1 9614 18802 9614 18802 0 tdc0.w_ring_int_norsz\[5\]
rlabel metal1 9292 19482 9292 19482 0 tdc0.w_ring_int_norsz\[6\]
rlabel via2 9890 19261 9890 19261 0 tdc0.w_ring_int_norsz\[7\]
rlabel metal1 10948 20774 10948 20774 0 tdc0.w_ring_int_norsz\[8\]
rlabel metal1 11086 13974 11086 13974 0 tdc0.w_ring_int_norsz\[9\]
rlabel metal1 4876 18190 4876 18190 0 tdc0.w_ring_norsz\[0\]
rlabel metal1 9752 14314 9752 14314 0 tdc0.w_ring_norsz\[10\]
rlabel metal1 8234 15062 8234 15062 0 tdc0.w_ring_norsz\[11\]
rlabel metal1 7452 16490 7452 16490 0 tdc0.w_ring_norsz\[12\]
rlabel metal1 6946 17544 6946 17544 0 tdc0.w_ring_norsz\[13\]
rlabel metal1 6348 19890 6348 19890 0 tdc0.w_ring_norsz\[14\]
rlabel metal1 5106 19856 5106 19856 0 tdc0.w_ring_norsz\[15\]
rlabel metal1 5244 15538 5244 15538 0 tdc0.w_ring_norsz\[16\]
rlabel metal1 5658 17850 5658 17850 0 tdc0.w_ring_norsz\[17\]
rlabel metal1 10856 17578 10856 17578 0 tdc0.w_ring_norsz\[18\]
rlabel metal2 10442 16320 10442 16320 0 tdc0.w_ring_norsz\[19\]
rlabel metal1 5428 17578 5428 17578 0 tdc0.w_ring_norsz\[1\]
rlabel metal1 10028 18394 10028 18394 0 tdc0.w_ring_norsz\[20\]
rlabel via1 9545 18666 9545 18666 0 tdc0.w_ring_norsz\[21\]
rlabel metal2 9890 20672 9890 20672 0 tdc0.w_ring_norsz\[22\]
rlabel metal1 10488 20026 10488 20026 0 tdc0.w_ring_norsz\[23\]
rlabel metal1 11040 14450 11040 14450 0 tdc0.w_ring_norsz\[24\]
rlabel metal1 10212 13702 10212 13702 0 tdc0.w_ring_norsz\[25\]
rlabel metal1 9982 14280 9982 14280 0 tdc0.w_ring_norsz\[26\]
rlabel metal1 8234 14926 8234 14926 0 tdc0.w_ring_norsz\[27\]
rlabel metal1 7130 16762 7130 16762 0 tdc0.w_ring_norsz\[28\]
rlabel via1 6849 17510 6849 17510 0 tdc0.w_ring_norsz\[29\]
rlabel metal1 11040 17850 11040 17850 0 tdc0.w_ring_norsz\[2\]
rlabel metal1 6670 18666 6670 18666 0 tdc0.w_ring_norsz\[30\]
rlabel metal1 5750 20366 5750 20366 0 tdc0.w_ring_norsz\[31\]
rlabel metal1 10028 17238 10028 17238 0 tdc0.w_ring_norsz\[3\]
rlabel metal1 10580 18326 10580 18326 0 tdc0.w_ring_norsz\[4\]
rlabel metal1 9430 19312 9430 19312 0 tdc0.w_ring_norsz\[5\]
rlabel metal2 8878 20128 8878 20128 0 tdc0.w_ring_norsz\[6\]
rlabel metal2 9798 19618 9798 19618 0 tdc0.w_ring_norsz\[7\]
rlabel metal1 11316 19414 11316 19414 0 tdc0.w_ring_norsz\[8\]
rlabel metal1 11270 13702 11270 13702 0 tdc0.w_ring_norsz\[9\]
rlabel metal1 22862 15028 22862 15028 0 tdc1.r_dly_store_ctr\[0\]
rlabel metal1 24564 11322 24564 11322 0 tdc1.r_dly_store_ctr\[10\]
rlabel metal2 22678 13430 22678 13430 0 tdc1.r_dly_store_ctr\[11\]
rlabel metal1 18308 14042 18308 14042 0 tdc1.r_dly_store_ctr\[12\]
rlabel metal2 20424 14212 20424 14212 0 tdc1.r_dly_store_ctr\[13\]
rlabel metal2 18906 14212 18906 14212 0 tdc1.r_dly_store_ctr\[14\]
rlabel metal2 23598 14790 23598 14790 0 tdc1.r_dly_store_ctr\[15\]
rlabel metal1 28014 15640 28014 15640 0 tdc1.r_dly_store_ctr\[1\]
rlabel metal1 30866 15674 30866 15674 0 tdc1.r_dly_store_ctr\[2\]
rlabel metal1 26073 14552 26073 14552 0 tdc1.r_dly_store_ctr\[3\]
rlabel metal1 24242 14586 24242 14586 0 tdc1.r_dly_store_ctr\[4\]
rlabel metal1 27370 15062 27370 15062 0 tdc1.r_dly_store_ctr\[5\]
rlabel metal1 20838 13498 20838 13498 0 tdc1.r_dly_store_ctr\[6\]
rlabel metal2 25254 15368 25254 15368 0 tdc1.r_dly_store_ctr\[7\]
rlabel metal1 20608 11866 20608 11866 0 tdc1.r_dly_store_ctr\[8\]
rlabel via1 22861 16014 22861 16014 0 tdc1.r_dly_store_ctr\[9\]
rlabel metal1 20608 15674 20608 15674 0 tdc1.r_dly_store_ring\[0\]
rlabel metal1 24794 19822 24794 19822 0 tdc1.r_dly_store_ring\[10\]
rlabel metal1 27048 17306 27048 17306 0 tdc1.r_dly_store_ring\[11\]
rlabel metal2 26358 16167 26358 16167 0 tdc1.r_dly_store_ring\[12\]
rlabel metal1 27186 18088 27186 18088 0 tdc1.r_dly_store_ring\[13\]
rlabel metal1 29026 20468 29026 20468 0 tdc1.r_dly_store_ring\[14\]
rlabel metal1 25438 20468 25438 20468 0 tdc1.r_dly_store_ring\[15\]
rlabel metal1 23138 14960 23138 14960 0 tdc1.r_dly_store_ring\[16\]
rlabel metal2 22770 20842 22770 20842 0 tdc1.r_dly_store_ring\[17\]
rlabel metal1 24472 19958 24472 19958 0 tdc1.r_dly_store_ring\[18\]
rlabel metal2 21666 16796 21666 16796 0 tdc1.r_dly_store_ring\[19\]
rlabel metal1 17664 20230 17664 20230 0 tdc1.r_dly_store_ring\[1\]
rlabel metal1 18446 16660 18446 16660 0 tdc1.r_dly_store_ring\[20\]
rlabel metal1 25944 18734 25944 18734 0 tdc1.r_dly_store_ring\[21\]
rlabel metal2 19274 17221 19274 17221 0 tdc1.r_dly_store_ring\[22\]
rlabel metal2 24150 19482 24150 19482 0 tdc1.r_dly_store_ring\[23\]
rlabel metal1 20930 13872 20930 13872 0 tdc1.r_dly_store_ring\[24\]
rlabel metal1 24459 17646 24459 17646 0 tdc1.r_dly_store_ring\[25\]
rlabel metal2 25530 16422 25530 16422 0 tdc1.r_dly_store_ring\[26\]
rlabel metal2 26726 16694 26726 16694 0 tdc1.r_dly_store_ring\[27\]
rlabel via2 18170 16643 18170 16643 0 tdc1.r_dly_store_ring\[28\]
rlabel metal1 28808 18734 28808 18734 0 tdc1.r_dly_store_ring\[29\]
rlabel metal1 16008 19346 16008 19346 0 tdc1.r_dly_store_ring\[2\]
rlabel via2 18998 17051 18998 17051 0 tdc1.r_dly_store_ring\[30\]
rlabel metal1 25576 19210 25576 19210 0 tdc1.r_dly_store_ring\[31\]
rlabel metal1 22954 16728 22954 16728 0 tdc1.r_dly_store_ring\[3\]
rlabel metal1 14996 17306 14996 17306 0 tdc1.r_dly_store_ring\[4\]
rlabel metal2 20470 16184 20470 16184 0 tdc1.r_dly_store_ring\[5\]
rlabel metal1 19228 20026 19228 20026 0 tdc1.r_dly_store_ring\[6\]
rlabel metal2 16698 21318 16698 21318 0 tdc1.r_dly_store_ring\[7\]
rlabel metal1 21850 14586 21850 14586 0 tdc1.r_dly_store_ring\[8\]
rlabel metal1 22816 20026 22816 20026 0 tdc1.r_dly_store_ring\[9\]
rlabel metal1 27738 11526 27738 11526 0 tdc1.r_ring_ctr\[0\]
rlabel metal1 23363 11186 23363 11186 0 tdc1.r_ring_ctr\[10\]
rlabel metal1 21390 11594 21390 11594 0 tdc1.r_ring_ctr\[11\]
rlabel metal2 17710 13328 17710 13328 0 tdc1.r_ring_ctr\[12\]
rlabel metal1 17802 12274 17802 12274 0 tdc1.r_ring_ctr\[13\]
rlabel metal1 17618 12648 17618 12648 0 tdc1.r_ring_ctr\[14\]
rlabel metal1 20838 13328 20838 13328 0 tdc1.r_ring_ctr\[15\]
rlabel metal1 28474 12342 28474 12342 0 tdc1.r_ring_ctr\[1\]
rlabel metal2 29118 15096 29118 15096 0 tdc1.r_ring_ctr\[2\]
rlabel metal1 29256 13362 29256 13362 0 tdc1.r_ring_ctr\[3\]
rlabel metal1 26588 13498 26588 13498 0 tdc1.r_ring_ctr\[4\]
rlabel metal2 26082 14450 26082 14450 0 tdc1.r_ring_ctr\[5\]
rlabel metal1 25070 12852 25070 12852 0 tdc1.r_ring_ctr\[6\]
rlabel metal1 25162 11730 25162 11730 0 tdc1.r_ring_ctr\[7\]
rlabel metal1 23598 10132 23598 10132 0 tdc1.r_ring_ctr\[8\]
rlabel metal1 25806 11152 25806 11152 0 tdc1.r_ring_ctr\[9\]
rlabel metal1 15548 11662 15548 11662 0 tdc1.w_dly_stop\[1\]
rlabel metal1 15778 11254 15778 11254 0 tdc1.w_dly_stop\[2\]
rlabel metal1 16146 11186 16146 11186 0 tdc1.w_dly_stop\[3\]
rlabel metal1 16698 11288 16698 11288 0 tdc1.w_dly_stop\[4\]
rlabel metal1 28842 11186 28842 11186 0 tdc1.w_dly_stop\[5\]
rlabel metal1 26496 13838 26496 13838 0 tdc1.w_ring_buf\[0\]
rlabel metal2 23046 19074 23046 19074 0 tdc1.w_ring_buf\[10\]
rlabel metal2 28106 16898 28106 16898 0 tdc1.w_ring_buf\[11\]
rlabel metal1 29306 16014 29306 16014 0 tdc1.w_ring_buf\[12\]
rlabel metal1 29752 18190 29752 18190 0 tdc1.w_ring_buf\[13\]
rlabel metal2 29946 20162 29946 20162 0 tdc1.w_ring_buf\[14\]
rlabel metal1 29404 20978 29404 20978 0 tdc1.w_ring_buf\[15\]
rlabel metal2 25990 18190 25990 18190 0 tdc1.w_ring_buf\[16\]
rlabel metal2 22218 21250 22218 21250 0 tdc1.w_ring_buf\[17\]
rlabel metal1 21965 21114 21965 21114 0 tdc1.w_ring_buf\[18\]
rlabel metal1 20362 17034 20362 17034 0 tdc1.w_ring_buf\[19\]
rlabel metal2 19090 21250 19090 21250 0 tdc1.w_ring_buf\[1\]
rlabel metal1 17337 16626 17337 16626 0 tdc1.w_ring_buf\[20\]
rlabel metal1 21022 18904 21022 18904 0 tdc1.w_ring_buf\[21\]
rlabel metal1 17429 17782 17429 17782 0 tdc1.w_ring_buf\[22\]
rlabel metal2 22126 19686 22126 19686 0 tdc1.w_ring_buf\[23\]
rlabel metal1 19350 14518 19350 14518 0 tdc1.w_ring_buf\[24\]
rlabel via1 23225 17782 23225 17782 0 tdc1.w_ring_buf\[25\]
rlabel metal1 24370 15946 24370 15946 0 tdc1.w_ring_buf\[26\]
rlabel metal2 27186 15810 27186 15810 0 tdc1.w_ring_buf\[27\]
rlabel metal1 30068 16694 30068 16694 0 tdc1.w_ring_buf\[28\]
rlabel metal1 30686 18870 30686 18870 0 tdc1.w_ring_buf\[29\]
rlabel metal1 14991 19890 14991 19890 0 tdc1.w_ring_buf\[2\]
rlabel via1 29941 17782 29941 17782 0 tdc1.w_ring_buf\[30\]
rlabel metal1 27512 19958 27512 19958 0 tdc1.w_ring_buf\[31\]
rlabel metal1 21558 17034 21558 17034 0 tdc1.w_ring_buf\[3\]
rlabel metal1 15966 17102 15966 17102 0 tdc1.w_ring_buf\[4\]
rlabel metal1 19223 16694 19223 16694 0 tdc1.w_ring_buf\[5\]
rlabel metal1 18717 19958 18717 19958 0 tdc1.w_ring_buf\[6\]
rlabel metal2 16882 20502 16882 20502 0 tdc1.w_ring_buf\[7\]
rlabel metal1 20454 14858 20454 14858 0 tdc1.w_ring_buf\[8\]
rlabel metal2 20930 19686 20930 19686 0 tdc1.w_ring_buf\[9\]
rlabel metal1 27186 21046 27186 21046 0 tdc1.w_ring_int_norsz\[0\]
rlabel metal1 21758 18122 21758 18122 0 tdc1.w_ring_int_norsz\[10\]
rlabel metal1 27370 16728 27370 16728 0 tdc1.w_ring_int_norsz\[11\]
rlabel metal1 29486 16762 29486 16762 0 tdc1.w_ring_int_norsz\[12\]
rlabel metal1 29072 17850 29072 17850 0 tdc1.w_ring_int_norsz\[13\]
rlabel metal1 29072 18938 29072 18938 0 tdc1.w_ring_int_norsz\[14\]
rlabel metal1 28658 19958 28658 19958 0 tdc1.w_ring_int_norsz\[15\]
rlabel metal2 27462 20672 27462 20672 0 tdc1.w_ring_int_norsz\[16\]
rlabel metal1 25024 20842 25024 20842 0 tdc1.w_ring_int_norsz\[17\]
rlabel metal1 21804 20910 21804 20910 0 tdc1.w_ring_int_norsz\[18\]
rlabel metal1 20746 19788 20746 19788 0 tdc1.w_ring_int_norsz\[19\]
rlabel metal1 25300 20910 25300 20910 0 tdc1.w_ring_int_norsz\[1\]
rlabel metal1 19826 17782 19826 17782 0 tdc1.w_ring_int_norsz\[20\]
rlabel metal1 18768 17850 18768 17850 0 tdc1.w_ring_int_norsz\[21\]
rlabel metal1 18446 18938 18446 18938 0 tdc1.w_ring_int_norsz\[22\]
rlabel metal2 17618 19652 17618 19652 0 tdc1.w_ring_int_norsz\[23\]
rlabel metal1 20237 19210 20237 19210 0 tdc1.w_ring_int_norsz\[24\]
rlabel metal1 20010 18734 20010 18734 0 tdc1.w_ring_int_norsz\[25\]
rlabel metal1 22586 18258 22586 18258 0 tdc1.w_ring_int_norsz\[26\]
rlabel metal1 26910 16558 26910 16558 0 tdc1.w_ring_int_norsz\[27\]
rlabel metal1 29302 16558 29302 16558 0 tdc1.w_ring_int_norsz\[28\]
rlabel metal2 29486 18054 29486 18054 0 tdc1.w_ring_int_norsz\[29\]
rlabel metal1 20884 20570 20884 20570 0 tdc1.w_ring_int_norsz\[2\]
rlabel metal1 29394 18904 29394 18904 0 tdc1.w_ring_int_norsz\[30\]
rlabel metal1 28566 20026 28566 20026 0 tdc1.w_ring_int_norsz\[31\]
rlabel metal1 20424 19958 20424 19958 0 tdc1.w_ring_int_norsz\[3\]
rlabel metal1 20148 17646 20148 17646 0 tdc1.w_ring_int_norsz\[4\]
rlabel metal1 19458 18122 19458 18122 0 tdc1.w_ring_int_norsz\[5\]
rlabel metal1 18124 18938 18124 18938 0 tdc1.w_ring_int_norsz\[6\]
rlabel metal2 16974 20366 16974 20366 0 tdc1.w_ring_int_norsz\[7\]
rlabel metal1 19366 19210 19366 19210 0 tdc1.w_ring_int_norsz\[8\]
rlabel metal1 20378 18870 20378 18870 0 tdc1.w_ring_int_norsz\[9\]
rlabel metal1 26082 20842 26082 20842 0 tdc1.w_ring_norsz\[0\]
rlabel metal1 23230 18734 23230 18734 0 tdc1.w_ring_norsz\[10\]
rlabel metal1 29762 16660 29762 16660 0 tdc1.w_ring_norsz\[11\]
rlabel metal2 29026 16286 29026 16286 0 tdc1.w_ring_norsz\[12\]
rlabel metal1 28980 18326 28980 18326 0 tdc1.w_ring_norsz\[13\]
rlabel metal1 29762 19822 29762 19822 0 tdc1.w_ring_norsz\[14\]
rlabel metal2 30038 20774 30038 20774 0 tdc1.w_ring_norsz\[15\]
rlabel metal1 27140 20842 27140 20842 0 tdc1.w_ring_norsz\[16\]
rlabel metal1 24794 21012 24794 21012 0 tdc1.w_ring_norsz\[17\]
rlabel metal1 20976 20842 20976 20842 0 tdc1.w_ring_norsz\[18\]
rlabel metal1 20332 19754 20332 19754 0 tdc1.w_ring_norsz\[19\]
rlabel metal2 20746 20689 20746 20689 0 tdc1.w_ring_norsz\[1\]
rlabel metal1 18722 17680 18722 17680 0 tdc1.w_ring_norsz\[20\]
rlabel metal1 18860 18802 18860 18802 0 tdc1.w_ring_norsz\[21\]
rlabel metal1 18009 19414 18009 19414 0 tdc1.w_ring_norsz\[22\]
rlabel metal1 20654 19312 20654 19312 0 tdc1.w_ring_norsz\[23\]
rlabel metal1 19090 14450 19090 14450 0 tdc1.w_ring_norsz\[24\]
rlabel metal1 22218 18258 22218 18258 0 tdc1.w_ring_norsz\[25\]
rlabel metal1 23690 16592 23690 16592 0 tdc1.w_ring_norsz\[26\]
rlabel metal1 27554 16456 27554 16456 0 tdc1.w_ring_norsz\[27\]
rlabel metal2 29118 16932 29118 16932 0 tdc1.w_ring_norsz\[28\]
rlabel metal2 28750 18598 28750 18598 0 tdc1.w_ring_norsz\[29\]
rlabel metal1 21068 20774 21068 20774 0 tdc1.w_ring_norsz\[2\]
rlabel metal1 29164 19414 29164 19414 0 tdc1.w_ring_norsz\[30\]
rlabel metal1 27830 20230 27830 20230 0 tdc1.w_ring_norsz\[31\]
rlabel metal1 20562 19720 20562 19720 0 tdc1.w_ring_norsz\[3\]
rlabel metal1 19366 17748 19366 17748 0 tdc1.w_ring_norsz\[4\]
rlabel metal1 19274 18054 19274 18054 0 tdc1.w_ring_norsz\[5\]
rlabel metal1 18170 19448 18170 19448 0 tdc1.w_ring_norsz\[6\]
rlabel metal1 17342 19754 17342 19754 0 tdc1.w_ring_norsz\[7\]
rlabel metal1 20148 14926 20148 14926 0 tdc1.w_ring_norsz\[8\]
rlabel metal2 20930 18394 20930 18394 0 tdc1.w_ring_norsz\[9\]
rlabel metal4 29532 22001 29532 22001 0 ui_in[0]
rlabel metal4 28796 21933 28796 21933 0 ui_in[1]
rlabel metal4 28060 22001 28060 22001 0 ui_in[2]
rlabel metal4 27324 22137 27324 22137 0 ui_in[3]
rlabel metal4 26588 22001 26588 22001 0 ui_in[4]
rlabel metal4 25852 22001 25852 22001 0 ui_in[5]
rlabel metal4 17756 19349 17756 19349 0 uo_out[0]
rlabel metal4 17020 21729 17020 21729 0 uo_out[1]
rlabel metal4 16284 22137 16284 22137 0 uo_out[2]
rlabel metal1 15824 16082 15824 16082 0 uo_out[3]
rlabel metal4 14812 20029 14812 20029 0 uo_out[4]
rlabel metal2 14674 19839 14674 19839 0 uo_out[5]
rlabel metal4 13340 21865 13340 21865 0 uo_out[6]
rlabel metal4 12604 21797 12604 21797 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
