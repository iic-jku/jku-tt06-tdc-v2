magic
tech sky130A
magscale 1 2
timestamp 1710691957
<< viali >>
rect 13829 18785 13863 18819
rect 13645 18581 13679 18615
rect 16497 12393 16531 12427
rect 16834 12325 16868 12359
rect 19441 12325 19475 12359
rect 11989 12257 12023 12291
rect 12148 12249 12182 12283
rect 12357 12257 12391 12291
rect 13134 12257 13168 12291
rect 13645 12257 13679 12291
rect 13829 12257 13863 12291
rect 14105 12257 14139 12291
rect 14372 12257 14406 12291
rect 16313 12257 16347 12291
rect 16589 12257 16623 12291
rect 19809 12257 19843 12291
rect 13047 12189 13081 12223
rect 12449 12121 12483 12155
rect 11897 12053 11931 12087
rect 12219 12053 12253 12087
rect 13553 12053 13587 12087
rect 13921 12053 13955 12087
rect 15485 12053 15519 12087
rect 17969 12053 18003 12087
rect 14657 11849 14691 11883
rect 16957 11849 16991 11883
rect 17325 11849 17359 11883
rect 20085 11849 20119 11883
rect 14105 11781 14139 11815
rect 15209 11781 15243 11815
rect 17141 11781 17175 11815
rect 14013 11713 14047 11747
rect 10885 11645 10919 11679
rect 10977 11645 11011 11679
rect 11253 11645 11287 11679
rect 11529 11645 11563 11679
rect 11796 11645 11830 11679
rect 13001 11645 13035 11679
rect 13737 11645 13771 11679
rect 14841 11645 14875 11679
rect 15485 11645 15519 11679
rect 16129 11645 16163 11679
rect 16221 11645 16255 11679
rect 16405 11645 16439 11679
rect 16497 11645 16531 11679
rect 16589 11645 16623 11679
rect 16773 11645 16807 11679
rect 17601 11645 17635 11679
rect 18705 11645 18739 11679
rect 18961 11645 18995 11679
rect 14473 11577 14507 11611
rect 15209 11577 15243 11611
rect 17293 11577 17327 11611
rect 17509 11577 17543 11611
rect 17693 11577 17727 11611
rect 10793 11509 10827 11543
rect 11069 11509 11103 11543
rect 11345 11509 11379 11543
rect 12909 11509 12943 11543
rect 13093 11509 13127 11543
rect 13921 11509 13955 11543
rect 15393 11509 15427 11543
rect 16313 11509 16347 11543
rect 11437 11305 11471 11339
rect 12173 11305 12207 11339
rect 13001 11305 13035 11339
rect 13737 11305 13771 11339
rect 15945 11305 15979 11339
rect 19809 11305 19843 11339
rect 20085 11305 20119 11339
rect 13369 11237 13403 11271
rect 14832 11237 14866 11271
rect 18674 11237 18708 11271
rect 19993 11237 20027 11271
rect 10517 11169 10551 11203
rect 10793 11169 10827 11203
rect 11161 11169 11195 11203
rect 11345 11169 11379 11203
rect 12081 11169 12115 11203
rect 12357 11169 12391 11203
rect 12561 11169 12595 11203
rect 12909 11169 12943 11203
rect 13553 11169 13587 11203
rect 14013 11169 14047 11203
rect 14105 11169 14139 11203
rect 14565 11169 14599 11203
rect 16129 11169 16163 11203
rect 16589 11169 16623 11203
rect 16865 11169 16899 11203
rect 17121 11169 17155 11203
rect 18429 11169 18463 11203
rect 10425 11033 10459 11067
rect 11069 11033 11103 11067
rect 16497 11033 16531 11067
rect 10701 10965 10735 10999
rect 12725 10965 12759 10999
rect 13921 10965 13955 10999
rect 14197 10965 14231 10999
rect 16221 10965 16255 10999
rect 18245 10965 18279 10999
rect 13737 10761 13771 10795
rect 14013 10761 14047 10795
rect 15393 10761 15427 10795
rect 15485 10761 15519 10795
rect 18889 10761 18923 10795
rect 14841 10625 14875 10659
rect 15301 10625 15335 10659
rect 9413 10557 9447 10591
rect 9873 10557 9907 10591
rect 9965 10557 9999 10591
rect 10241 10557 10275 10591
rect 12357 10557 12391 10591
rect 12817 10557 12851 10591
rect 12909 10557 12943 10591
rect 13185 10557 13219 10591
rect 13369 10557 13403 10591
rect 13829 10557 13863 10591
rect 13921 10557 13955 10591
rect 14381 10557 14415 10591
rect 14590 10557 14624 10591
rect 14749 10557 14783 10591
rect 15577 10557 15611 10591
rect 15761 10557 15795 10591
rect 15945 10557 15979 10591
rect 16129 10557 16163 10591
rect 16221 10557 16255 10591
rect 16589 10557 16623 10591
rect 16865 10557 16899 10591
rect 16957 10557 16991 10591
rect 17233 10557 17267 10591
rect 17509 10557 17543 10591
rect 17785 10557 17819 10591
rect 18061 10557 18095 10591
rect 18337 10557 18371 10591
rect 18797 10557 18831 10591
rect 19257 10557 19291 10591
rect 19349 10557 19383 10591
rect 19533 10557 19567 10591
rect 19809 10557 19843 10591
rect 9781 10489 9815 10523
rect 10486 10489 10520 10523
rect 11805 10489 11839 10523
rect 12449 10489 12483 10523
rect 13001 10489 13035 10523
rect 15853 10489 15887 10523
rect 16773 10489 16807 10523
rect 17877 10489 17911 10523
rect 9505 10421 9539 10455
rect 10057 10421 10091 10455
rect 11621 10421 11655 10455
rect 11897 10421 11931 10455
rect 12725 10421 12759 10455
rect 13277 10421 13311 10455
rect 14289 10421 14323 10455
rect 14519 10421 14553 10455
rect 16497 10421 16531 10455
rect 17049 10421 17083 10455
rect 17325 10421 17359 10455
rect 17601 10421 17635 10455
rect 18153 10421 18187 10455
rect 18429 10421 18463 10455
rect 19625 10421 19659 10455
rect 19901 10421 19935 10455
rect 9045 10217 9079 10251
rect 9413 10217 9447 10251
rect 10149 10217 10183 10251
rect 10701 10217 10735 10251
rect 11345 10217 11379 10251
rect 12495 10217 12529 10251
rect 12725 10217 12759 10251
rect 13185 10217 13219 10251
rect 13737 10217 13771 10251
rect 15301 10217 15335 10251
rect 19717 10217 19751 10251
rect 11897 10149 11931 10183
rect 14188 10149 14222 10183
rect 15485 10149 15519 10183
rect 18604 10149 18638 10183
rect 19901 10149 19935 10183
rect 20269 10149 20303 10183
rect 8861 10081 8895 10115
rect 9137 10081 9171 10115
rect 9229 10081 9263 10115
rect 9413 10081 9447 10115
rect 9505 10081 9539 10115
rect 9597 10081 9631 10115
rect 9781 10081 9815 10115
rect 10241 10081 10275 10115
rect 10333 10081 10367 10115
rect 10609 10081 10643 10115
rect 10793 10081 10827 10115
rect 10977 10081 11011 10115
rect 11253 10081 11287 10115
rect 11529 10081 11563 10115
rect 11805 10081 11839 10115
rect 12081 10081 12115 10115
rect 12424 10081 12458 10115
rect 12817 10081 12851 10115
rect 13001 10081 13035 10115
rect 13093 10081 13127 10115
rect 13369 10081 13403 10115
rect 13645 10081 13679 10115
rect 16313 10081 16347 10115
rect 16589 10081 16623 10115
rect 16856 10081 16890 10115
rect 18245 10081 18279 10115
rect 18337 10081 18371 10115
rect 20361 10081 20395 10115
rect 12173 10013 12207 10047
rect 13921 10013 13955 10047
rect 18153 9945 18187 9979
rect 8769 9877 8803 9911
rect 9873 9877 9907 9911
rect 10425 9877 10459 9911
rect 11069 9877 11103 9911
rect 11621 9877 11655 9911
rect 15577 9877 15611 9911
rect 16405 9877 16439 9911
rect 17969 9877 18003 9911
rect 20453 9877 20487 9911
rect 11345 9673 11379 9707
rect 16405 9673 16439 9707
rect 18061 9673 18095 9707
rect 8677 9605 8711 9639
rect 10885 9605 10919 9639
rect 13921 9605 13955 9639
rect 18981 9605 19015 9639
rect 19901 9605 19935 9639
rect 8953 9537 8987 9571
rect 8217 9469 8251 9503
rect 8769 9469 8803 9503
rect 8861 9469 8895 9503
rect 9137 9469 9171 9503
rect 9404 9469 9438 9503
rect 11437 9469 11471 9503
rect 13588 9469 13622 9503
rect 13691 9469 13725 9503
rect 13829 9469 13863 9503
rect 14105 9469 14139 9503
rect 16221 9469 16255 9503
rect 16497 9469 16531 9503
rect 19257 9469 19291 9503
rect 19441 9469 19475 9503
rect 19533 9469 19567 9503
rect 19625 9469 19659 9503
rect 19809 9469 19843 9503
rect 20269 9469 20303 9503
rect 20453 9469 20487 9503
rect 20545 9469 20579 9503
rect 20637 9469 20671 9503
rect 8125 9401 8159 9435
rect 10701 9401 10735 9435
rect 13277 9401 13311 9435
rect 16589 9401 16623 9435
rect 18797 9401 18831 9435
rect 10517 9333 10551 9367
rect 11989 9333 12023 9367
rect 15393 9333 15427 9367
rect 16129 9333 16163 9367
rect 19257 9333 19291 9367
rect 20177 9333 20211 9367
rect 20729 9333 20763 9367
rect 8401 9129 8435 9163
rect 15209 9129 15243 9163
rect 15853 9129 15887 9163
rect 16221 9129 16255 9163
rect 19625 9129 19659 9163
rect 20085 9129 20119 9163
rect 11989 9061 12023 9095
rect 13645 9061 13679 9095
rect 16405 9061 16439 9095
rect 18512 9061 18546 9095
rect 19809 9061 19843 9095
rect 7849 8993 7883 9027
rect 7941 8993 7975 9027
rect 8217 8993 8251 9027
rect 8401 8993 8435 9027
rect 8677 8993 8711 9027
rect 8861 8993 8895 9027
rect 8953 8993 8987 9027
rect 9045 8993 9079 9027
rect 9312 8993 9346 9027
rect 10609 8993 10643 9027
rect 11069 8993 11103 9027
rect 11621 8993 11655 9027
rect 13921 8993 13955 9027
rect 15945 8993 15979 9027
rect 16129 8993 16163 9027
rect 18245 8993 18279 9027
rect 20361 8993 20395 9027
rect 20821 8993 20855 9027
rect 21281 8993 21315 9027
rect 21557 8993 21591 9027
rect 21649 8925 21683 8959
rect 7757 8857 7791 8891
rect 10425 8857 10459 8891
rect 10701 8857 10735 8891
rect 20637 8857 20671 8891
rect 8033 8789 8067 8823
rect 8585 8789 8619 8823
rect 11161 8789 11195 8823
rect 11713 8789 11747 8823
rect 17693 8789 17727 8823
rect 20913 8789 20947 8823
rect 21373 8789 21407 8823
rect 10241 8585 10275 8619
rect 10517 8585 10551 8619
rect 11345 8585 11379 8619
rect 17141 8585 17175 8619
rect 17417 8585 17451 8619
rect 20085 8585 20119 8619
rect 11069 8517 11103 8551
rect 12173 8517 12207 8551
rect 13277 8517 13311 8551
rect 17693 8517 17727 8551
rect 17969 8517 18003 8551
rect 18245 8517 18279 8551
rect 8125 8449 8159 8483
rect 9137 8449 9171 8483
rect 13553 8449 13587 8483
rect 18705 8449 18739 8483
rect 8217 8381 8251 8415
rect 8493 8381 8527 8415
rect 8677 8381 8711 8415
rect 8953 8381 8987 8415
rect 9045 8381 9079 8415
rect 9321 8381 9355 8415
rect 9781 8381 9815 8415
rect 9965 8381 9999 8415
rect 10057 8381 10091 8415
rect 10333 8381 10367 8415
rect 10425 8381 10459 8415
rect 10701 8381 10735 8415
rect 11161 8381 11195 8415
rect 11253 8381 11287 8415
rect 11713 8381 11747 8415
rect 11989 8381 12023 8415
rect 12081 8381 12115 8415
rect 12541 8381 12575 8415
rect 12633 8381 12667 8415
rect 13001 8381 13035 8415
rect 13093 8381 13127 8415
rect 13369 8381 13403 8415
rect 13809 8381 13843 8415
rect 15853 8381 15887 8415
rect 16129 8381 16163 8415
rect 16405 8381 16439 8415
rect 16681 8381 16715 8415
rect 16957 8391 16991 8425
rect 17049 8381 17083 8415
rect 17325 8381 17359 8415
rect 17785 8381 17819 8415
rect 17877 8381 17911 8415
rect 18153 8381 18187 8415
rect 20177 8381 20211 8415
rect 20361 8381 20395 8415
rect 20453 8381 20487 8415
rect 20545 8381 20579 8415
rect 20729 8381 20763 8415
rect 8585 8313 8619 8347
rect 9413 8313 9447 8347
rect 9689 8313 9723 8347
rect 11621 8313 11655 8347
rect 15117 8313 15151 8347
rect 18972 8313 19006 8347
rect 20269 8313 20303 8347
rect 8861 8245 8895 8279
rect 10793 8245 10827 8279
rect 11897 8245 11931 8279
rect 12449 8245 12483 8279
rect 12725 8245 12759 8279
rect 14933 8245 14967 8279
rect 15209 8245 15243 8279
rect 16037 8245 16071 8279
rect 16313 8245 16347 8279
rect 16589 8245 16623 8279
rect 16865 8245 16899 8279
rect 20821 8245 20855 8279
rect 8677 8041 8711 8075
rect 10517 8041 10551 8075
rect 11161 8041 11195 8075
rect 13645 8041 13679 8075
rect 14105 8041 14139 8075
rect 14381 8041 14415 8075
rect 14657 8041 14691 8075
rect 15853 8041 15887 8075
rect 19717 8041 19751 8075
rect 9382 7973 9416 8007
rect 11069 7973 11103 8007
rect 13829 7973 13863 8007
rect 15209 7973 15243 8007
rect 19901 7973 19935 8007
rect 8769 7905 8803 7939
rect 9045 7905 9079 7939
rect 10609 7905 10643 7939
rect 11529 7905 11563 7939
rect 11805 7905 11839 7939
rect 12265 7905 12299 7939
rect 12357 7905 12391 7939
rect 12541 7905 12575 7939
rect 12809 7905 12843 7939
rect 12901 7895 12935 7929
rect 13369 7905 13403 7939
rect 13461 7905 13495 7939
rect 13645 7905 13679 7939
rect 13921 7905 13955 7939
rect 14197 7905 14231 7939
rect 14473 7905 14507 7939
rect 14749 7905 14783 7939
rect 15025 7905 15059 7939
rect 15301 7905 15335 7939
rect 15577 7905 15611 7939
rect 15669 7905 15703 7939
rect 15853 7905 15887 7939
rect 16313 7905 16347 7939
rect 16589 7905 16623 7939
rect 16865 7905 16899 7939
rect 17132 7905 17166 7939
rect 18337 7905 18371 7939
rect 18604 7905 18638 7939
rect 20361 7905 20395 7939
rect 9137 7837 9171 7871
rect 12173 7837 12207 7871
rect 20453 7837 20487 7871
rect 13001 7769 13035 7803
rect 14933 7769 14967 7803
rect 16221 7769 16255 7803
rect 8953 7701 8987 7735
rect 10701 7701 10735 7735
rect 11621 7701 11655 7735
rect 11897 7701 11931 7735
rect 12449 7701 12483 7735
rect 12725 7701 12759 7735
rect 13277 7701 13311 7735
rect 15485 7701 15519 7735
rect 16681 7701 16715 7735
rect 18245 7701 18279 7735
rect 19993 7701 20027 7735
rect 9965 7497 9999 7531
rect 13277 7497 13311 7531
rect 18337 7497 18371 7531
rect 19625 7497 19659 7531
rect 19901 7429 19935 7463
rect 13553 7361 13587 7395
rect 15393 7361 15427 7395
rect 9597 7293 9631 7327
rect 9873 7293 9907 7327
rect 10057 7293 10091 7327
rect 10241 7293 10275 7327
rect 10333 7293 10367 7327
rect 10425 7293 10459 7327
rect 10885 7293 10919 7327
rect 10977 7293 11011 7327
rect 13185 7293 13219 7327
rect 15117 7293 15151 7327
rect 17417 7293 17451 7327
rect 17693 7293 17727 7327
rect 17969 7293 18003 7327
rect 18061 7293 18095 7327
rect 18245 7293 18279 7327
rect 18797 7293 18831 7327
rect 19257 7293 19291 7327
rect 19533 7293 19567 7327
rect 19809 7293 19843 7327
rect 9689 7225 9723 7259
rect 11244 7225 11278 7259
rect 12541 7225 12575 7259
rect 13820 7225 13854 7259
rect 15660 7225 15694 7259
rect 16957 7225 16991 7259
rect 17785 7225 17819 7259
rect 19349 7225 19383 7259
rect 10517 7157 10551 7191
rect 10793 7157 10827 7191
rect 12357 7157 12391 7191
rect 12633 7157 12667 7191
rect 14933 7157 14967 7191
rect 15209 7157 15243 7191
rect 16773 7157 16807 7191
rect 17049 7157 17083 7191
rect 17509 7157 17543 7191
rect 18889 7157 18923 7191
rect 13369 6953 13403 6987
rect 13645 6953 13679 6987
rect 13921 6953 13955 6987
rect 14473 6953 14507 6987
rect 15853 6953 15887 6987
rect 16221 6953 16255 6987
rect 17969 6953 18003 6987
rect 14749 6885 14783 6919
rect 10057 6817 10091 6851
rect 10149 6817 10183 6851
rect 10325 6817 10359 6851
rect 10609 6817 10643 6851
rect 10977 6817 11011 6851
rect 11437 6817 11471 6851
rect 11529 6817 11563 6851
rect 11805 6817 11839 6851
rect 12081 6817 12115 6851
rect 12449 6815 12483 6849
rect 12725 6817 12759 6851
rect 13001 6817 13035 6851
rect 13277 6817 13311 6851
rect 13737 6817 13771 6851
rect 14013 6817 14047 6851
rect 14105 6817 14139 6851
rect 15117 6817 15151 6851
rect 15209 6817 15243 6851
rect 15485 6817 15519 6851
rect 15945 6817 15979 6851
rect 16129 6817 16163 6851
rect 16497 6817 16531 6851
rect 16589 6817 16623 6851
rect 16773 6817 16807 6851
rect 17049 6817 17083 6851
rect 17233 6817 17267 6851
rect 17325 6817 17359 6851
rect 17417 6817 17451 6851
rect 17601 6817 17635 6851
rect 18061 6817 18095 6851
rect 18153 6807 18187 6841
rect 18245 6817 18279 6851
rect 18613 6817 18647 6851
rect 11621 6749 11655 6783
rect 11897 6749 11931 6783
rect 12541 6749 12575 6783
rect 11345 6681 11379 6715
rect 12173 6681 12207 6715
rect 15577 6681 15611 6715
rect 18521 6681 18555 6715
rect 10425 6613 10459 6647
rect 10701 6613 10735 6647
rect 11069 6613 11103 6647
rect 12817 6613 12851 6647
rect 13093 6613 13127 6647
rect 14197 6613 14231 6647
rect 16865 6613 16899 6647
rect 17141 6613 17175 6647
rect 17693 6613 17727 6647
rect 10977 6409 11011 6443
rect 11529 6409 11563 6443
rect 11805 6409 11839 6443
rect 13185 6409 13219 6443
rect 13921 6409 13955 6443
rect 14565 6409 14599 6443
rect 16129 6409 16163 6443
rect 13645 6341 13679 6375
rect 11253 6273 11287 6307
rect 10885 6205 10919 6239
rect 11069 6205 11103 6239
rect 11161 6205 11195 6239
rect 11621 6205 11655 6239
rect 11897 6205 11931 6239
rect 11989 6205 12023 6239
rect 12265 6205 12299 6239
rect 12541 6205 12575 6239
rect 12817 6205 12851 6239
rect 13277 6205 13311 6239
rect 13553 6205 13587 6239
rect 14013 6205 14047 6239
rect 14105 6205 14139 6239
rect 14657 6205 14691 6239
rect 14841 6205 14875 6239
rect 15117 6205 15151 6239
rect 15301 6205 15335 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 16037 6205 16071 6239
rect 12081 6069 12115 6103
rect 12357 6069 12391 6103
rect 12633 6069 12667 6103
rect 12909 6069 12943 6103
rect 14197 6069 14231 6103
rect 14933 6069 14967 6103
rect 15117 6069 15151 6103
rect 12265 5865 12299 5899
rect 12725 5865 12759 5899
rect 13921 5865 13955 5899
rect 11345 5797 11379 5831
rect 11253 5729 11287 5763
rect 12357 5729 12391 5763
rect 12633 5729 12667 5763
rect 12909 5729 12943 5763
rect 13093 5729 13127 5763
rect 14013 5729 14047 5763
rect 13001 5661 13035 5695
<< metal1 >>
rect 552 19066 31531 19088
rect 552 19014 8102 19066
rect 8154 19014 8166 19066
rect 8218 19014 8230 19066
rect 8282 19014 8294 19066
rect 8346 19014 8358 19066
rect 8410 19014 15807 19066
rect 15859 19014 15871 19066
rect 15923 19014 15935 19066
rect 15987 19014 15999 19066
rect 16051 19014 16063 19066
rect 16115 19014 23512 19066
rect 23564 19014 23576 19066
rect 23628 19014 23640 19066
rect 23692 19014 23704 19066
rect 23756 19014 23768 19066
rect 23820 19014 31217 19066
rect 31269 19014 31281 19066
rect 31333 19014 31345 19066
rect 31397 19014 31409 19066
rect 31461 19014 31473 19066
rect 31525 19014 31531 19066
rect 552 18992 31531 19014
rect 13538 18912 13544 18964
rect 13596 18912 13602 18964
rect 13556 18816 13584 18912
rect 13817 18819 13875 18825
rect 13817 18816 13829 18819
rect 13556 18788 13829 18816
rect 13817 18785 13829 18788
rect 13863 18785 13875 18819
rect 13817 18779 13875 18785
rect 13630 18572 13636 18624
rect 13688 18572 13694 18624
rect 552 18522 31372 18544
rect 552 18470 4250 18522
rect 4302 18470 4314 18522
rect 4366 18470 4378 18522
rect 4430 18470 4442 18522
rect 4494 18470 4506 18522
rect 4558 18470 11955 18522
rect 12007 18470 12019 18522
rect 12071 18470 12083 18522
rect 12135 18470 12147 18522
rect 12199 18470 12211 18522
rect 12263 18470 19660 18522
rect 19712 18470 19724 18522
rect 19776 18470 19788 18522
rect 19840 18470 19852 18522
rect 19904 18470 19916 18522
rect 19968 18470 27365 18522
rect 27417 18470 27429 18522
rect 27481 18470 27493 18522
rect 27545 18470 27557 18522
rect 27609 18470 27621 18522
rect 27673 18470 31372 18522
rect 552 18448 31372 18470
rect 552 17978 31531 18000
rect 552 17926 8102 17978
rect 8154 17926 8166 17978
rect 8218 17926 8230 17978
rect 8282 17926 8294 17978
rect 8346 17926 8358 17978
rect 8410 17926 15807 17978
rect 15859 17926 15871 17978
rect 15923 17926 15935 17978
rect 15987 17926 15999 17978
rect 16051 17926 16063 17978
rect 16115 17926 23512 17978
rect 23564 17926 23576 17978
rect 23628 17926 23640 17978
rect 23692 17926 23704 17978
rect 23756 17926 23768 17978
rect 23820 17926 31217 17978
rect 31269 17926 31281 17978
rect 31333 17926 31345 17978
rect 31397 17926 31409 17978
rect 31461 17926 31473 17978
rect 31525 17926 31531 17978
rect 552 17904 31531 17926
rect 552 17434 31372 17456
rect 552 17382 4250 17434
rect 4302 17382 4314 17434
rect 4366 17382 4378 17434
rect 4430 17382 4442 17434
rect 4494 17382 4506 17434
rect 4558 17382 11955 17434
rect 12007 17382 12019 17434
rect 12071 17382 12083 17434
rect 12135 17382 12147 17434
rect 12199 17382 12211 17434
rect 12263 17382 19660 17434
rect 19712 17382 19724 17434
rect 19776 17382 19788 17434
rect 19840 17382 19852 17434
rect 19904 17382 19916 17434
rect 19968 17382 27365 17434
rect 27417 17382 27429 17434
rect 27481 17382 27493 17434
rect 27545 17382 27557 17434
rect 27609 17382 27621 17434
rect 27673 17382 31372 17434
rect 552 17360 31372 17382
rect 552 16890 31531 16912
rect 552 16838 8102 16890
rect 8154 16838 8166 16890
rect 8218 16838 8230 16890
rect 8282 16838 8294 16890
rect 8346 16838 8358 16890
rect 8410 16838 15807 16890
rect 15859 16838 15871 16890
rect 15923 16838 15935 16890
rect 15987 16838 15999 16890
rect 16051 16838 16063 16890
rect 16115 16838 23512 16890
rect 23564 16838 23576 16890
rect 23628 16838 23640 16890
rect 23692 16838 23704 16890
rect 23756 16838 23768 16890
rect 23820 16838 31217 16890
rect 31269 16838 31281 16890
rect 31333 16838 31345 16890
rect 31397 16838 31409 16890
rect 31461 16838 31473 16890
rect 31525 16838 31531 16890
rect 552 16816 31531 16838
rect 552 16346 31372 16368
rect 552 16294 4250 16346
rect 4302 16294 4314 16346
rect 4366 16294 4378 16346
rect 4430 16294 4442 16346
rect 4494 16294 4506 16346
rect 4558 16294 11955 16346
rect 12007 16294 12019 16346
rect 12071 16294 12083 16346
rect 12135 16294 12147 16346
rect 12199 16294 12211 16346
rect 12263 16294 19660 16346
rect 19712 16294 19724 16346
rect 19776 16294 19788 16346
rect 19840 16294 19852 16346
rect 19904 16294 19916 16346
rect 19968 16294 27365 16346
rect 27417 16294 27429 16346
rect 27481 16294 27493 16346
rect 27545 16294 27557 16346
rect 27609 16294 27621 16346
rect 27673 16294 31372 16346
rect 552 16272 31372 16294
rect 552 15802 31531 15824
rect 552 15750 8102 15802
rect 8154 15750 8166 15802
rect 8218 15750 8230 15802
rect 8282 15750 8294 15802
rect 8346 15750 8358 15802
rect 8410 15750 15807 15802
rect 15859 15750 15871 15802
rect 15923 15750 15935 15802
rect 15987 15750 15999 15802
rect 16051 15750 16063 15802
rect 16115 15750 23512 15802
rect 23564 15750 23576 15802
rect 23628 15750 23640 15802
rect 23692 15750 23704 15802
rect 23756 15750 23768 15802
rect 23820 15750 31217 15802
rect 31269 15750 31281 15802
rect 31333 15750 31345 15802
rect 31397 15750 31409 15802
rect 31461 15750 31473 15802
rect 31525 15750 31531 15802
rect 552 15728 31531 15750
rect 552 15258 31372 15280
rect 552 15206 4250 15258
rect 4302 15206 4314 15258
rect 4366 15206 4378 15258
rect 4430 15206 4442 15258
rect 4494 15206 4506 15258
rect 4558 15206 11955 15258
rect 12007 15206 12019 15258
rect 12071 15206 12083 15258
rect 12135 15206 12147 15258
rect 12199 15206 12211 15258
rect 12263 15206 19660 15258
rect 19712 15206 19724 15258
rect 19776 15206 19788 15258
rect 19840 15206 19852 15258
rect 19904 15206 19916 15258
rect 19968 15206 27365 15258
rect 27417 15206 27429 15258
rect 27481 15206 27493 15258
rect 27545 15206 27557 15258
rect 27609 15206 27621 15258
rect 27673 15206 31372 15258
rect 552 15184 31372 15206
rect 552 14714 31531 14736
rect 552 14662 8102 14714
rect 8154 14662 8166 14714
rect 8218 14662 8230 14714
rect 8282 14662 8294 14714
rect 8346 14662 8358 14714
rect 8410 14662 15807 14714
rect 15859 14662 15871 14714
rect 15923 14662 15935 14714
rect 15987 14662 15999 14714
rect 16051 14662 16063 14714
rect 16115 14662 23512 14714
rect 23564 14662 23576 14714
rect 23628 14662 23640 14714
rect 23692 14662 23704 14714
rect 23756 14662 23768 14714
rect 23820 14662 31217 14714
rect 31269 14662 31281 14714
rect 31333 14662 31345 14714
rect 31397 14662 31409 14714
rect 31461 14662 31473 14714
rect 31525 14662 31531 14714
rect 552 14640 31531 14662
rect 552 14170 31372 14192
rect 552 14118 4250 14170
rect 4302 14118 4314 14170
rect 4366 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 11955 14170
rect 12007 14118 12019 14170
rect 12071 14118 12083 14170
rect 12135 14118 12147 14170
rect 12199 14118 12211 14170
rect 12263 14118 19660 14170
rect 19712 14118 19724 14170
rect 19776 14118 19788 14170
rect 19840 14118 19852 14170
rect 19904 14118 19916 14170
rect 19968 14118 27365 14170
rect 27417 14118 27429 14170
rect 27481 14118 27493 14170
rect 27545 14118 27557 14170
rect 27609 14118 27621 14170
rect 27673 14118 31372 14170
rect 552 14096 31372 14118
rect 552 13626 31531 13648
rect 552 13574 8102 13626
rect 8154 13574 8166 13626
rect 8218 13574 8230 13626
rect 8282 13574 8294 13626
rect 8346 13574 8358 13626
rect 8410 13574 15807 13626
rect 15859 13574 15871 13626
rect 15923 13574 15935 13626
rect 15987 13574 15999 13626
rect 16051 13574 16063 13626
rect 16115 13574 23512 13626
rect 23564 13574 23576 13626
rect 23628 13574 23640 13626
rect 23692 13574 23704 13626
rect 23756 13574 23768 13626
rect 23820 13574 31217 13626
rect 31269 13574 31281 13626
rect 31333 13574 31345 13626
rect 31397 13574 31409 13626
rect 31461 13574 31473 13626
rect 31525 13574 31531 13626
rect 552 13552 31531 13574
rect 552 13082 31372 13104
rect 552 13030 4250 13082
rect 4302 13030 4314 13082
rect 4366 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 11955 13082
rect 12007 13030 12019 13082
rect 12071 13030 12083 13082
rect 12135 13030 12147 13082
rect 12199 13030 12211 13082
rect 12263 13030 19660 13082
rect 19712 13030 19724 13082
rect 19776 13030 19788 13082
rect 19840 13030 19852 13082
rect 19904 13030 19916 13082
rect 19968 13030 27365 13082
rect 27417 13030 27429 13082
rect 27481 13030 27493 13082
rect 27545 13030 27557 13082
rect 27609 13030 27621 13082
rect 27673 13030 31372 13082
rect 552 13008 31372 13030
rect 552 12538 31531 12560
rect 552 12486 8102 12538
rect 8154 12486 8166 12538
rect 8218 12486 8230 12538
rect 8282 12486 8294 12538
rect 8346 12486 8358 12538
rect 8410 12486 15807 12538
rect 15859 12486 15871 12538
rect 15923 12486 15935 12538
rect 15987 12486 15999 12538
rect 16051 12486 16063 12538
rect 16115 12486 23512 12538
rect 23564 12486 23576 12538
rect 23628 12486 23640 12538
rect 23692 12486 23704 12538
rect 23756 12486 23768 12538
rect 23820 12486 31217 12538
rect 31269 12486 31281 12538
rect 31333 12486 31345 12538
rect 31397 12486 31409 12538
rect 31461 12486 31473 12538
rect 31525 12486 31531 12538
rect 552 12464 31531 12486
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 12250 12424 12256 12436
rect 11664 12396 12256 12424
rect 11664 12384 11670 12396
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 16485 12427 16543 12433
rect 12406 12396 13676 12424
rect 12406 12356 12434 12396
rect 11992 12328 12434 12356
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11992 12297 12020 12328
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 11756 12260 11989 12288
rect 11756 12248 11762 12260
rect 11977 12257 11989 12260
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12136 12288 12194 12289
rect 12136 12283 12296 12288
rect 12136 12249 12148 12283
rect 12182 12260 12296 12283
rect 12182 12252 12204 12260
rect 12182 12249 12194 12252
rect 12136 12243 12194 12249
rect 12268 12220 12296 12260
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 13648 12297 13676 12396
rect 16485 12393 16497 12427
rect 16531 12393 16543 12427
rect 16485 12387 16543 12393
rect 16500 12356 16528 12387
rect 16822 12359 16880 12365
rect 16822 12356 16834 12359
rect 14108 12328 16436 12356
rect 16500 12328 16834 12356
rect 14108 12300 14136 12328
rect 13122 12291 13180 12297
rect 13122 12288 13134 12291
rect 12676 12260 13134 12288
rect 12676 12248 12682 12260
rect 13122 12257 13134 12260
rect 13168 12257 13180 12291
rect 13122 12251 13180 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13817 12291 13875 12297
rect 13817 12288 13829 12291
rect 13679 12260 13829 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13817 12257 13829 12260
rect 13863 12288 13875 12291
rect 13863 12260 14044 12288
rect 13863 12257 13875 12260
rect 13817 12251 13875 12257
rect 13035 12223 13093 12229
rect 13035 12220 13047 12223
rect 12268 12192 13047 12220
rect 13035 12189 13047 12192
rect 13081 12189 13093 12223
rect 13035 12183 13093 12189
rect 10962 12112 10968 12164
rect 11020 12152 11026 12164
rect 12437 12155 12495 12161
rect 12437 12152 12449 12155
rect 11020 12124 12449 12152
rect 11020 12112 11026 12124
rect 12437 12121 12449 12124
rect 12483 12121 12495 12155
rect 12437 12115 12495 12121
rect 14016 12096 14044 12260
rect 14090 12248 14096 12300
rect 14148 12248 14154 12300
rect 14360 12291 14418 12297
rect 14360 12257 14372 12291
rect 14406 12288 14418 12291
rect 14642 12288 14648 12300
rect 14406 12260 14648 12288
rect 14406 12257 14418 12260
rect 14360 12251 14418 12257
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 16298 12248 16304 12300
rect 16356 12248 16362 12300
rect 16408 12288 16436 12328
rect 16822 12325 16834 12328
rect 16868 12325 16880 12359
rect 16822 12319 16880 12325
rect 19426 12316 19432 12368
rect 19484 12316 19490 12368
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16408 12260 16589 12288
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12288 19855 12291
rect 20070 12288 20076 12300
rect 19843 12260 20076 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 11885 12087 11943 12093
rect 11885 12084 11897 12087
rect 11848 12056 11897 12084
rect 11848 12044 11854 12056
rect 11885 12053 11897 12056
rect 11931 12053 11943 12087
rect 11885 12047 11943 12053
rect 12207 12087 12265 12093
rect 12207 12053 12219 12087
rect 12253 12084 12265 12087
rect 12342 12084 12348 12096
rect 12253 12056 12348 12084
rect 12253 12053 12265 12056
rect 12207 12047 12265 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 13538 12044 13544 12096
rect 13596 12044 13602 12096
rect 13906 12044 13912 12096
rect 13964 12044 13970 12096
rect 13998 12044 14004 12096
rect 14056 12044 14062 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 15436 12056 15485 12084
rect 15436 12044 15442 12056
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 15473 12047 15531 12053
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 18782 12084 18788 12096
rect 18003 12056 18788 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 18782 12044 18788 12056
rect 18840 12044 18846 12096
rect 552 11994 31372 12016
rect 552 11942 4250 11994
rect 4302 11942 4314 11994
rect 4366 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 11955 11994
rect 12007 11942 12019 11994
rect 12071 11942 12083 11994
rect 12135 11942 12147 11994
rect 12199 11942 12211 11994
rect 12263 11942 19660 11994
rect 19712 11942 19724 11994
rect 19776 11942 19788 11994
rect 19840 11942 19852 11994
rect 19904 11942 19916 11994
rect 19968 11942 27365 11994
rect 27417 11942 27429 11994
rect 27481 11942 27493 11994
rect 27545 11942 27557 11994
rect 27609 11942 27621 11994
rect 27673 11942 31372 11994
rect 552 11920 31372 11942
rect 13906 11840 13912 11892
rect 13964 11840 13970 11892
rect 14642 11840 14648 11892
rect 14700 11840 14706 11892
rect 16298 11840 16304 11892
rect 16356 11840 16362 11892
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 16991 11852 17325 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 17313 11849 17325 11852
rect 17359 11849 17371 11883
rect 17313 11843 17371 11849
rect 20070 11840 20076 11892
rect 20128 11840 20134 11892
rect 13924 11812 13952 11840
rect 14093 11815 14151 11821
rect 14093 11812 14105 11815
rect 13924 11784 14105 11812
rect 14093 11781 14105 11784
rect 14139 11781 14151 11815
rect 14093 11775 14151 11781
rect 15010 11772 15016 11824
rect 15068 11812 15074 11824
rect 15197 11815 15255 11821
rect 15197 11812 15209 11815
rect 15068 11784 15209 11812
rect 15068 11772 15074 11784
rect 15197 11781 15209 11784
rect 15243 11781 15255 11815
rect 16316 11812 16344 11840
rect 17129 11815 17187 11821
rect 17129 11812 17141 11815
rect 16316 11784 17141 11812
rect 15197 11775 15255 11781
rect 17129 11781 17141 11784
rect 17175 11781 17187 11815
rect 17129 11775 17187 11781
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 14001 11747 14059 11753
rect 8996 11716 11284 11744
rect 8996 11704 9002 11716
rect 10870 11636 10876 11688
rect 10928 11636 10934 11688
rect 11256 11685 11284 11716
rect 14001 11713 14013 11747
rect 14047 11744 14059 11747
rect 14047 11716 14872 11744
rect 14047 11713 14059 11716
rect 14001 11707 14059 11713
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 10980 11608 11008 11639
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 11790 11685 11796 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11480 11648 11529 11676
rect 11480 11636 11486 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11784 11676 11796 11685
rect 11751 11648 11796 11676
rect 11517 11639 11575 11645
rect 11784 11639 11796 11648
rect 11790 11636 11796 11639
rect 11848 11636 11854 11688
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 12989 11679 13047 11685
rect 12989 11676 13001 11679
rect 12216 11648 13001 11676
rect 12216 11636 12222 11648
rect 12989 11645 13001 11648
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 13722 11636 13728 11688
rect 13780 11636 13786 11688
rect 14090 11636 14096 11688
rect 14148 11636 14154 11688
rect 14844 11685 14872 11716
rect 15488 11716 16252 11744
rect 15488 11688 15516 11716
rect 14829 11679 14887 11685
rect 14829 11645 14841 11679
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 15470 11636 15476 11688
rect 15528 11636 15534 11688
rect 16224 11685 16252 11716
rect 16408 11716 18828 11744
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 16298 11676 16304 11688
rect 16255 11648 16304 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 10980 11580 11284 11608
rect 11256 11552 11284 11580
rect 10778 11500 10784 11552
rect 10836 11500 10842 11552
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11146 11540 11152 11552
rect 11103 11512 11152 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11238 11500 11244 11552
rect 11296 11500 11302 11552
rect 11333 11543 11391 11549
rect 11333 11509 11345 11543
rect 11379 11540 11391 11543
rect 11790 11540 11796 11552
rect 11379 11512 11796 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12894 11500 12900 11552
rect 12952 11500 12958 11552
rect 13078 11500 13084 11552
rect 13136 11500 13142 11552
rect 13909 11543 13967 11549
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 14108 11540 14136 11636
rect 14461 11611 14519 11617
rect 14461 11577 14473 11611
rect 14507 11577 14519 11611
rect 14461 11571 14519 11577
rect 13955 11512 14136 11540
rect 14476 11540 14504 11571
rect 15194 11568 15200 11620
rect 15252 11568 15258 11620
rect 16132 11608 16160 11639
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 16408 11685 16436 11716
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 16482 11636 16488 11688
rect 16540 11636 16546 11688
rect 16776 11685 16804 11716
rect 18800 11688 18828 11716
rect 16577 11679 16635 11685
rect 16577 11645 16589 11679
rect 16623 11645 16635 11679
rect 16577 11639 16635 11645
rect 16761 11679 16819 11685
rect 16761 11645 16773 11679
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 16592 11608 16620 11639
rect 16850 11636 16856 11688
rect 16908 11676 16914 11688
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 16908 11648 17601 11676
rect 16908 11636 16914 11648
rect 17589 11645 17601 11648
rect 17635 11645 17647 11679
rect 17589 11639 17647 11645
rect 18414 11636 18420 11688
rect 18472 11676 18478 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18472 11648 18705 11676
rect 18472 11636 18478 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 18949 11679 19007 11685
rect 18949 11676 18961 11679
rect 18840 11648 18961 11676
rect 18840 11636 18846 11648
rect 18949 11645 18961 11648
rect 18995 11645 19007 11679
rect 18949 11639 19007 11645
rect 17281 11611 17339 11617
rect 17281 11608 17293 11611
rect 15396 11580 16620 11608
rect 16684 11580 17293 11608
rect 15396 11552 15424 11580
rect 16224 11552 16252 11580
rect 15378 11540 15384 11552
rect 14476 11512 15384 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 16206 11500 16212 11552
rect 16264 11500 16270 11552
rect 16301 11543 16359 11549
rect 16301 11509 16313 11543
rect 16347 11540 16359 11543
rect 16684 11540 16712 11580
rect 17281 11577 17293 11580
rect 17327 11577 17339 11611
rect 17281 11571 17339 11577
rect 17497 11611 17555 11617
rect 17497 11577 17509 11611
rect 17543 11608 17555 11611
rect 17681 11611 17739 11617
rect 17681 11608 17693 11611
rect 17543 11580 17693 11608
rect 17543 11577 17555 11580
rect 17497 11571 17555 11577
rect 17681 11577 17693 11580
rect 17727 11577 17739 11611
rect 17681 11571 17739 11577
rect 16347 11512 16712 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 552 11450 31531 11472
rect 552 11398 8102 11450
rect 8154 11398 8166 11450
rect 8218 11398 8230 11450
rect 8282 11398 8294 11450
rect 8346 11398 8358 11450
rect 8410 11398 15807 11450
rect 15859 11398 15871 11450
rect 15923 11398 15935 11450
rect 15987 11398 15999 11450
rect 16051 11398 16063 11450
rect 16115 11398 23512 11450
rect 23564 11398 23576 11450
rect 23628 11398 23640 11450
rect 23692 11398 23704 11450
rect 23756 11398 23768 11450
rect 23820 11398 31217 11450
rect 31269 11398 31281 11450
rect 31333 11398 31345 11450
rect 31397 11398 31409 11450
rect 31461 11398 31473 11450
rect 31525 11398 31531 11450
rect 552 11376 31531 11398
rect 11425 11339 11483 11345
rect 11425 11305 11437 11339
rect 11471 11336 11483 11339
rect 11698 11336 11704 11348
rect 11471 11308 11704 11336
rect 11471 11305 11483 11308
rect 11425 11299 11483 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12158 11296 12164 11348
rect 12216 11296 12222 11348
rect 12342 11296 12348 11348
rect 12400 11296 12406 11348
rect 12894 11296 12900 11348
rect 12952 11296 12958 11348
rect 12986 11296 12992 11348
rect 13044 11296 13050 11348
rect 13538 11336 13544 11348
rect 13372 11308 13544 11336
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 10928 11240 11192 11268
rect 10928 11228 10934 11240
rect 10502 11160 10508 11212
rect 10560 11160 10566 11212
rect 11164 11209 11192 11240
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 10796 11132 10824 11163
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 12360 11209 12388 11296
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 11296 11172 11345 11200
rect 11296 11160 11302 11172
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 12069 11203 12127 11209
rect 12069 11169 12081 11203
rect 12115 11169 12127 11203
rect 12069 11163 12127 11169
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 12084 11132 12112 11163
rect 12526 11160 12532 11212
rect 12584 11209 12590 11212
rect 12912 11209 12940 11296
rect 13372 11277 13400 11308
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 13722 11296 13728 11348
rect 13780 11296 13786 11348
rect 14090 11296 14096 11348
rect 14148 11296 14154 11348
rect 15010 11296 15016 11348
rect 15068 11296 15074 11348
rect 15933 11339 15991 11345
rect 15933 11305 15945 11339
rect 15979 11336 15991 11339
rect 16482 11336 16488 11348
rect 15979 11308 16488 11336
rect 15979 11305 15991 11308
rect 15933 11299 15991 11305
rect 16482 11296 16488 11308
rect 16540 11336 16546 11348
rect 19797 11339 19855 11345
rect 16540 11308 18552 11336
rect 16540 11296 16546 11308
rect 13357 11271 13415 11277
rect 13357 11237 13369 11271
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 13630 11228 13636 11280
rect 13688 11228 13694 11280
rect 14108 11268 14136 11296
rect 14820 11271 14878 11277
rect 14108 11240 14596 11268
rect 12584 11203 12607 11209
rect 12595 11200 12607 11203
rect 12897 11203 12955 11209
rect 12595 11172 12848 11200
rect 12595 11169 12607 11172
rect 12584 11163 12607 11169
rect 12584 11160 12590 11163
rect 12820 11132 12848 11172
rect 12897 11169 12909 11203
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 13648 11200 13676 11228
rect 13587 11172 13676 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 13556 11132 13584 11163
rect 13998 11160 14004 11212
rect 14056 11160 14062 11212
rect 14568 11209 14596 11240
rect 14820 11237 14832 11271
rect 14866 11268 14878 11271
rect 15028 11268 15056 11296
rect 18524 11268 18552 11308
rect 19797 11305 19809 11339
rect 19843 11336 19855 11339
rect 19843 11308 20024 11336
rect 19843 11305 19855 11308
rect 19797 11299 19855 11305
rect 19996 11277 20024 11308
rect 20070 11296 20076 11348
rect 20128 11296 20134 11348
rect 18662 11271 18720 11277
rect 18662 11268 18674 11271
rect 14866 11240 15056 11268
rect 16868 11240 18460 11268
rect 18524 11240 18674 11268
rect 14866 11237 14878 11240
rect 14820 11231 14878 11237
rect 14093 11203 14151 11209
rect 14093 11169 14105 11203
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 10796 11104 12388 11132
rect 12820 11104 13584 11132
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 10413 11067 10471 11073
rect 10413 11064 10425 11067
rect 9364 11036 10425 11064
rect 9364 11024 9370 11036
rect 10413 11033 10425 11036
rect 10459 11033 10471 11067
rect 10413 11027 10471 11033
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 11057 11067 11115 11073
rect 11057 11064 11069 11067
rect 10652 11036 11069 11064
rect 10652 11024 10658 11036
rect 11057 11033 11069 11036
rect 11103 11033 11115 11067
rect 11057 11027 11115 11033
rect 12360 11008 12388 11104
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14108 11132 14136 11163
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 16117 11203 16175 11209
rect 16117 11200 16129 11203
rect 15160 11172 16129 11200
rect 15160 11160 15166 11172
rect 16117 11169 16129 11172
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 16574 11160 16580 11212
rect 16632 11160 16638 11212
rect 16868 11209 16896 11240
rect 18432 11212 18460 11240
rect 18662 11237 18674 11240
rect 18708 11237 18720 11271
rect 18662 11231 18720 11237
rect 19981 11271 20039 11277
rect 19981 11237 19993 11271
rect 20027 11237 20039 11271
rect 19981 11231 20039 11237
rect 16853 11203 16911 11209
rect 16853 11169 16865 11203
rect 16899 11169 16911 11203
rect 17109 11203 17167 11209
rect 17109 11200 17121 11203
rect 16853 11163 16911 11169
rect 16960 11172 17121 11200
rect 13872 11104 14136 11132
rect 13872 11092 13878 11104
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 16758 11132 16764 11144
rect 15620 11104 16764 11132
rect 15620 11092 15626 11104
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16960 11132 16988 11172
rect 17109 11169 17121 11172
rect 17155 11169 17167 11203
rect 17109 11163 17167 11169
rect 18414 11160 18420 11212
rect 18472 11160 18478 11212
rect 16868 11104 16988 11132
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 16485 11067 16543 11073
rect 16485 11064 16497 11067
rect 16356 11036 16497 11064
rect 16356 11024 16362 11036
rect 16485 11033 16497 11036
rect 16531 11033 16543 11067
rect 16868 11064 16896 11104
rect 16485 11027 16543 11033
rect 16592 11036 16896 11064
rect 10686 10956 10692 11008
rect 10744 10956 10750 11008
rect 12342 10956 12348 11008
rect 12400 10956 12406 11008
rect 12713 10999 12771 11005
rect 12713 10965 12725 10999
rect 12759 10996 12771 10999
rect 13078 10996 13084 11008
rect 12759 10968 13084 10996
rect 12759 10965 12771 10968
rect 12713 10959 12771 10965
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 13906 10956 13912 11008
rect 13964 10956 13970 11008
rect 14182 10956 14188 11008
rect 14240 10956 14246 11008
rect 16206 10956 16212 11008
rect 16264 10956 16270 11008
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 16592 10996 16620 11036
rect 16448 10968 16620 10996
rect 18233 10999 18291 11005
rect 16448 10956 16454 10968
rect 18233 10965 18245 10999
rect 18279 10996 18291 10999
rect 18598 10996 18604 11008
rect 18279 10968 18604 10996
rect 18279 10965 18291 10968
rect 18233 10959 18291 10965
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 552 10906 31372 10928
rect 552 10854 4250 10906
rect 4302 10854 4314 10906
rect 4366 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 11955 10906
rect 12007 10854 12019 10906
rect 12071 10854 12083 10906
rect 12135 10854 12147 10906
rect 12199 10854 12211 10906
rect 12263 10854 19660 10906
rect 19712 10854 19724 10906
rect 19776 10854 19788 10906
rect 19840 10854 19852 10906
rect 19904 10854 19916 10906
rect 19968 10854 27365 10906
rect 27417 10854 27429 10906
rect 27481 10854 27493 10906
rect 27545 10854 27557 10906
rect 27609 10854 27621 10906
rect 27673 10854 31372 10906
rect 552 10832 31372 10854
rect 13725 10795 13783 10801
rect 10152 10764 11652 10792
rect 9030 10548 9036 10600
rect 9088 10588 9094 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 9088 10560 9413 10588
rect 9088 10548 9094 10560
rect 9401 10557 9413 10560
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 9950 10588 9956 10600
rect 9907 10560 9956 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 9950 10548 9956 10560
rect 10008 10588 10014 10600
rect 10152 10588 10180 10764
rect 11624 10736 11652 10764
rect 13725 10761 13737 10795
rect 13771 10792 13783 10795
rect 13814 10792 13820 10804
rect 13771 10764 13820 10792
rect 13771 10761 13783 10764
rect 13725 10755 13783 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 13906 10752 13912 10804
rect 13964 10752 13970 10804
rect 14001 10795 14059 10801
rect 14001 10761 14013 10795
rect 14047 10792 14059 10795
rect 14182 10792 14188 10804
rect 14047 10764 14188 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 15194 10752 15200 10804
rect 15252 10792 15258 10804
rect 15381 10795 15439 10801
rect 15381 10792 15393 10795
rect 15252 10764 15393 10792
rect 15252 10752 15258 10764
rect 15381 10761 15393 10764
rect 15427 10761 15439 10795
rect 15381 10755 15439 10761
rect 15470 10752 15476 10804
rect 15528 10752 15534 10804
rect 16206 10752 16212 10804
rect 16264 10752 16270 10804
rect 18874 10752 18880 10804
rect 18932 10752 18938 10804
rect 11606 10684 11612 10736
rect 11664 10684 11670 10736
rect 13924 10724 13952 10752
rect 13372 10696 13952 10724
rect 12434 10656 12440 10668
rect 11440 10628 12440 10656
rect 11440 10600 11468 10628
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 13262 10656 13268 10668
rect 12820 10628 13268 10656
rect 10008 10560 10180 10588
rect 10229 10591 10287 10597
rect 10008 10548 10014 10560
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 11422 10588 11428 10600
rect 10275 10560 11428 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 12820 10597 12848 10628
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 12345 10591 12403 10597
rect 12345 10557 12357 10591
rect 12391 10557 12403 10591
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12345 10551 12403 10557
rect 12452 10560 12817 10588
rect 9769 10523 9827 10529
rect 9769 10489 9781 10523
rect 9815 10520 9827 10523
rect 10474 10523 10532 10529
rect 10474 10520 10486 10523
rect 9815 10492 10486 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 10474 10489 10486 10492
rect 10520 10489 10532 10523
rect 11793 10523 11851 10529
rect 11793 10520 11805 10523
rect 10474 10483 10532 10489
rect 11624 10492 11805 10520
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 9456 10424 9505 10452
rect 9456 10412 9462 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 11330 10452 11336 10464
rect 10091 10424 11336 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 11624 10461 11652 10492
rect 11793 10489 11805 10492
rect 11839 10489 11851 10523
rect 11793 10483 11851 10489
rect 12360 10464 12388 10551
rect 12452 10529 12480 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 12437 10523 12495 10529
rect 12437 10489 12449 10523
rect 12483 10489 12495 10523
rect 12437 10483 12495 10489
rect 12912 10464 12940 10551
rect 13170 10548 13176 10600
rect 13228 10548 13234 10600
rect 13372 10597 13400 10696
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 16224 10724 16252 10752
rect 14148 10696 15516 10724
rect 14148 10684 14154 10696
rect 13722 10616 13728 10668
rect 13780 10656 13786 10668
rect 13780 10628 14504 10656
rect 13780 10616 13786 10628
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 13814 10548 13820 10600
rect 13872 10548 13878 10600
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10557 14427 10591
rect 14476 10588 14504 10628
rect 14752 10597 14780 10696
rect 15488 10668 15516 10696
rect 15764 10696 16252 10724
rect 16960 10696 17356 10724
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 14875 10628 15301 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15378 10616 15384 10668
rect 15436 10616 15442 10668
rect 15470 10616 15476 10668
rect 15528 10616 15534 10668
rect 14578 10591 14636 10597
rect 14578 10588 14590 10591
rect 14476 10560 14590 10588
rect 14369 10551 14427 10557
rect 14578 10557 14590 10560
rect 14624 10557 14636 10591
rect 14578 10551 14636 10557
rect 14737 10591 14795 10597
rect 14737 10557 14749 10591
rect 14783 10557 14795 10591
rect 14737 10551 14795 10557
rect 12989 10523 13047 10529
rect 12989 10489 13001 10523
rect 13035 10520 13047 10523
rect 13924 10520 13952 10551
rect 13035 10492 13952 10520
rect 13035 10489 13047 10492
rect 12989 10483 13047 10489
rect 13998 10480 14004 10532
rect 14056 10520 14062 10532
rect 14384 10520 14412 10551
rect 15102 10548 15108 10600
rect 15160 10548 15166 10600
rect 15396 10588 15424 10616
rect 15764 10597 15792 10696
rect 16758 10656 16764 10668
rect 16224 10628 16764 10656
rect 16224 10597 16252 10628
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 15396 10560 15577 10588
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 15749 10591 15807 10597
rect 15749 10557 15761 10591
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10588 15991 10591
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15979 10560 16129 10588
rect 15979 10557 15991 10560
rect 15933 10551 15991 10557
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16577 10591 16635 10597
rect 16577 10557 16589 10591
rect 16623 10588 16635 10591
rect 16666 10588 16672 10600
rect 16623 10560 16672 10588
rect 16623 10557 16635 10560
rect 16577 10551 16635 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 16960 10597 16988 10696
rect 16853 10591 16911 10597
rect 16853 10557 16865 10591
rect 16899 10588 16911 10591
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16899 10560 16957 10588
rect 16899 10557 16911 10560
rect 16853 10551 16911 10557
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10557 17279 10591
rect 17328 10588 17356 10696
rect 17788 10696 19840 10724
rect 17788 10597 17816 10696
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 17920 10628 19288 10656
rect 17920 10616 17926 10628
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 17328 10560 17509 10588
rect 17221 10551 17279 10557
rect 17497 10557 17509 10560
rect 17543 10557 17555 10591
rect 17497 10551 17555 10557
rect 17773 10591 17831 10597
rect 17773 10557 17785 10591
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 15120 10520 15148 10548
rect 14056 10492 15148 10520
rect 15841 10523 15899 10529
rect 14056 10480 14062 10492
rect 15841 10489 15853 10523
rect 15887 10520 15899 10523
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 15887 10492 16773 10520
rect 15887 10489 15899 10492
rect 15841 10483 15899 10489
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 16761 10483 16819 10489
rect 11609 10455 11667 10461
rect 11609 10421 11621 10455
rect 11655 10421 11667 10455
rect 11609 10415 11667 10421
rect 11882 10412 11888 10464
rect 11940 10412 11946 10464
rect 12342 10412 12348 10464
rect 12400 10412 12406 10464
rect 12710 10412 12716 10464
rect 12768 10412 12774 10464
rect 12894 10412 12900 10464
rect 12952 10412 12958 10464
rect 13262 10412 13268 10464
rect 13320 10412 13326 10464
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 14016 10452 14044 10480
rect 13412 10424 14044 10452
rect 13412 10412 13418 10424
rect 14274 10412 14280 10464
rect 14332 10412 14338 10464
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 14507 10455 14565 10461
rect 14507 10452 14519 10455
rect 14424 10424 14519 10452
rect 14424 10412 14430 10424
rect 14507 10421 14519 10424
rect 14553 10421 14565 10455
rect 14507 10415 14565 10421
rect 16482 10412 16488 10464
rect 16540 10412 16546 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16868 10452 16896 10551
rect 17236 10520 17264 10551
rect 17788 10520 17816 10551
rect 18046 10548 18052 10600
rect 18104 10548 18110 10600
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 17052 10492 17264 10520
rect 17512 10492 17816 10520
rect 17865 10523 17923 10529
rect 17052 10461 17080 10492
rect 17512 10464 17540 10492
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 18230 10520 18236 10532
rect 17911 10492 18236 10520
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 18230 10480 18236 10492
rect 18288 10480 18294 10532
rect 18340 10520 18368 10551
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 19260 10597 19288 10628
rect 19812 10597 19840 10696
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18656 10560 18797 10588
rect 18656 10548 18662 10560
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 18785 10551 18843 10557
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19337 10591 19395 10597
rect 19337 10557 19349 10591
rect 19383 10588 19395 10591
rect 19521 10591 19579 10597
rect 19521 10588 19533 10591
rect 19383 10560 19533 10588
rect 19383 10557 19395 10560
rect 19337 10551 19395 10557
rect 19521 10557 19533 10560
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 20530 10588 20536 10600
rect 19843 10560 20536 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 19058 10520 19064 10532
rect 18340 10492 19064 10520
rect 19058 10480 19064 10492
rect 19116 10480 19122 10532
rect 16632 10424 16896 10452
rect 17037 10455 17095 10461
rect 16632 10412 16638 10424
rect 17037 10421 17049 10455
rect 17083 10421 17095 10455
rect 17037 10415 17095 10421
rect 17310 10412 17316 10464
rect 17368 10412 17374 10464
rect 17494 10412 17500 10464
rect 17552 10412 17558 10464
rect 17586 10412 17592 10464
rect 17644 10412 17650 10464
rect 18138 10412 18144 10464
rect 18196 10412 18202 10464
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 19518 10452 19524 10464
rect 18463 10424 19524 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19610 10412 19616 10464
rect 19668 10412 19674 10464
rect 19889 10455 19947 10461
rect 19889 10421 19901 10455
rect 19935 10452 19947 10455
rect 20162 10452 20168 10464
rect 19935 10424 20168 10452
rect 19935 10421 19947 10424
rect 19889 10415 19947 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 552 10362 31531 10384
rect 552 10310 8102 10362
rect 8154 10310 8166 10362
rect 8218 10310 8230 10362
rect 8282 10310 8294 10362
rect 8346 10310 8358 10362
rect 8410 10310 15807 10362
rect 15859 10310 15871 10362
rect 15923 10310 15935 10362
rect 15987 10310 15999 10362
rect 16051 10310 16063 10362
rect 16115 10310 23512 10362
rect 23564 10310 23576 10362
rect 23628 10310 23640 10362
rect 23692 10310 23704 10362
rect 23756 10310 23768 10362
rect 23820 10310 31217 10362
rect 31269 10310 31281 10362
rect 31333 10310 31345 10362
rect 31397 10310 31409 10362
rect 31461 10310 31473 10362
rect 31525 10310 31531 10362
rect 552 10288 31531 10310
rect 9030 10208 9036 10260
rect 9088 10208 9094 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 9447 10220 10149 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 10502 10208 10508 10260
rect 10560 10208 10566 10260
rect 10594 10208 10600 10260
rect 10652 10208 10658 10260
rect 10686 10208 10692 10260
rect 10744 10208 10750 10260
rect 10962 10248 10968 10260
rect 10796 10220 10968 10248
rect 10410 10180 10416 10192
rect 9232 10152 10416 10180
rect 9232 10121 9260 10152
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 8849 10115 8907 10121
rect 8849 10081 8861 10115
rect 8895 10081 8907 10115
rect 8849 10075 8907 10081
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10081 9459 10115
rect 9401 10075 9459 10081
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8260 9880 8769 9908
rect 8260 9868 8266 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8864 9908 8892 10075
rect 9140 9976 9168 10075
rect 9416 10044 9444 10075
rect 9490 10072 9496 10124
rect 9548 10072 9554 10124
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 10520 10112 10548 10208
rect 10612 10121 10640 10208
rect 10796 10121 10824 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11146 10208 11152 10260
rect 11204 10208 11210 10260
rect 11330 10208 11336 10260
rect 11388 10208 11394 10260
rect 11698 10208 11704 10260
rect 11756 10208 11762 10260
rect 12483 10251 12541 10257
rect 12483 10217 12495 10251
rect 12529 10248 12541 10251
rect 12618 10248 12624 10260
rect 12529 10220 12624 10248
rect 12529 10217 12541 10220
rect 12483 10211 12541 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12710 10208 12716 10260
rect 12768 10208 12774 10260
rect 12986 10208 12992 10260
rect 13044 10208 13050 10260
rect 13078 10208 13084 10260
rect 13136 10208 13142 10260
rect 13170 10208 13176 10260
rect 13228 10208 13234 10260
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 13320 10220 13737 10248
rect 13320 10208 13326 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 13725 10211 13783 10217
rect 13814 10208 13820 10260
rect 13872 10208 13878 10260
rect 14274 10208 14280 10260
rect 14332 10208 14338 10260
rect 15289 10251 15347 10257
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 16574 10248 16580 10260
rect 15335 10220 15516 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 10367 10084 10548 10112
rect 10597 10115 10655 10121
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 10597 10081 10609 10115
rect 10643 10081 10655 10115
rect 10597 10075 10655 10081
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 9858 10044 9864 10056
rect 9416 10016 9864 10044
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10244 10044 10272 10075
rect 10962 10072 10968 10124
rect 11020 10072 11026 10124
rect 11164 10112 11192 10208
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 11164 10084 11253 10112
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 11514 10072 11520 10124
rect 11572 10072 11578 10124
rect 11716 10112 11744 10208
rect 11885 10183 11943 10189
rect 11885 10149 11897 10183
rect 11931 10180 11943 10183
rect 13004 10180 13032 10208
rect 11931 10152 13032 10180
rect 13096 10180 13124 10208
rect 13096 10152 13216 10180
rect 11931 10149 11943 10152
rect 11885 10143 11943 10149
rect 11793 10115 11851 10121
rect 11793 10112 11805 10115
rect 11716 10084 11805 10112
rect 11793 10081 11805 10084
rect 11839 10081 11851 10115
rect 11793 10075 11851 10081
rect 12069 10115 12127 10121
rect 12069 10081 12081 10115
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12412 10115 12470 10121
rect 12412 10081 12424 10115
rect 12458 10112 12470 10115
rect 12526 10112 12532 10124
rect 12458 10084 12532 10112
rect 12458 10081 12470 10084
rect 12412 10075 12470 10081
rect 10686 10044 10692 10056
rect 10244 10016 10692 10044
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 12084 10044 12112 10075
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12851 10084 13001 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13188 10112 13216 10152
rect 13357 10115 13415 10121
rect 13188 10111 13308 10112
rect 13357 10111 13369 10115
rect 13188 10084 13369 10111
rect 13280 10083 13369 10084
rect 13081 10075 13139 10081
rect 13357 10081 13369 10083
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10081 13691 10115
rect 13832 10112 13860 10208
rect 14176 10183 14234 10189
rect 14176 10149 14188 10183
rect 14222 10180 14234 10183
rect 14292 10180 14320 10208
rect 15488 10189 15516 10220
rect 16224 10220 16580 10248
rect 14222 10152 14320 10180
rect 15473 10183 15531 10189
rect 14222 10149 14234 10152
rect 14176 10143 14234 10149
rect 15473 10149 15485 10183
rect 15519 10149 15531 10183
rect 15473 10143 15531 10149
rect 15654 10112 15660 10124
rect 13832 10084 15660 10112
rect 13633 10075 13691 10081
rect 11664 10016 12112 10044
rect 12161 10047 12219 10053
rect 11664 10004 11670 10016
rect 12161 10013 12173 10047
rect 12207 10044 12219 10047
rect 12894 10044 12900 10056
rect 12207 10016 12900 10044
rect 12207 10013 12219 10016
rect 12161 10007 12219 10013
rect 12894 10004 12900 10016
rect 12952 10044 12958 10056
rect 13096 10044 13124 10075
rect 13648 10044 13676 10075
rect 15654 10072 15660 10084
rect 15712 10112 15718 10124
rect 16224 10112 16252 10220
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 19610 10208 19616 10260
rect 19668 10208 19674 10260
rect 19705 10251 19763 10257
rect 19705 10217 19717 10251
rect 19751 10248 19763 10251
rect 19751 10220 19932 10248
rect 19751 10217 19763 10220
rect 19705 10211 19763 10217
rect 18592 10183 18650 10189
rect 16592 10152 18368 10180
rect 15712 10084 16252 10112
rect 15712 10072 15718 10084
rect 16298 10072 16304 10124
rect 16356 10072 16362 10124
rect 16592 10121 16620 10152
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10081 16635 10115
rect 16577 10075 16635 10081
rect 16844 10115 16902 10121
rect 16844 10081 16856 10115
rect 16890 10112 16902 10115
rect 17310 10112 17316 10124
rect 16890 10084 17316 10112
rect 16890 10081 16902 10084
rect 16844 10075 16902 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18340 10121 18368 10152
rect 18592 10149 18604 10183
rect 18638 10180 18650 10183
rect 19628 10180 19656 10208
rect 19904 10189 19932 10220
rect 20162 10208 20168 10260
rect 20220 10208 20226 10260
rect 18638 10152 19656 10180
rect 19889 10183 19947 10189
rect 18638 10149 18650 10152
rect 18592 10143 18650 10149
rect 19889 10149 19901 10183
rect 19935 10149 19947 10183
rect 19889 10143 19947 10149
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 18414 10112 18420 10124
rect 18371 10084 18420 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 12952 10016 13676 10044
rect 13909 10047 13967 10053
rect 12952 10004 12958 10016
rect 13909 10013 13921 10047
rect 13955 10013 13967 10047
rect 13909 10007 13967 10013
rect 9490 9976 9496 9988
rect 9140 9948 9496 9976
rect 9490 9936 9496 9948
rect 9548 9976 9554 9988
rect 10226 9976 10232 9988
rect 9548 9948 10232 9976
rect 9548 9936 9554 9948
rect 10226 9936 10232 9948
rect 10284 9976 10290 9988
rect 10502 9976 10508 9988
rect 10284 9948 10508 9976
rect 10284 9936 10290 9948
rect 10502 9936 10508 9948
rect 10560 9976 10566 9988
rect 10962 9976 10968 9988
rect 10560 9948 10968 9976
rect 10560 9936 10566 9948
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 9674 9908 9680 9920
rect 8864 9880 9680 9908
rect 8757 9871 8815 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9861 9911 9919 9917
rect 9861 9877 9873 9911
rect 9907 9908 9919 9911
rect 10042 9908 10048 9920
rect 9907 9880 10048 9908
rect 9907 9877 9919 9880
rect 9861 9871 9919 9877
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 10594 9908 10600 9920
rect 10459 9880 10600 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 11057 9911 11115 9917
rect 11057 9877 11069 9911
rect 11103 9908 11115 9911
rect 11422 9908 11428 9920
rect 11103 9880 11428 9908
rect 11103 9877 11115 9880
rect 11057 9871 11115 9877
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11606 9868 11612 9920
rect 11664 9868 11670 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13538 9908 13544 9920
rect 12492 9880 13544 9908
rect 12492 9868 12498 9880
rect 13538 9868 13544 9880
rect 13596 9908 13602 9920
rect 13924 9908 13952 10007
rect 17862 10004 17868 10056
rect 17920 10044 17926 10056
rect 18248 10044 18276 10075
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 20180 10112 20208 10208
rect 20257 10183 20315 10189
rect 20257 10149 20269 10183
rect 20303 10180 20315 10183
rect 31662 10180 31668 10192
rect 20303 10152 31668 10180
rect 20303 10149 20315 10152
rect 20257 10143 20315 10149
rect 31662 10140 31668 10152
rect 31720 10140 31726 10192
rect 20349 10115 20407 10121
rect 20349 10112 20361 10115
rect 20180 10084 20361 10112
rect 20349 10081 20361 10084
rect 20395 10081 20407 10115
rect 20349 10075 20407 10081
rect 17920 10016 18276 10044
rect 17920 10004 17926 10016
rect 17770 9936 17776 9988
rect 17828 9976 17834 9988
rect 18141 9979 18199 9985
rect 18141 9976 18153 9979
rect 17828 9948 18153 9976
rect 17828 9936 17834 9948
rect 18141 9945 18153 9948
rect 18187 9945 18199 9979
rect 18141 9939 18199 9945
rect 13596 9880 13952 9908
rect 13596 9868 13602 9880
rect 15562 9868 15568 9920
rect 15620 9868 15626 9920
rect 16390 9868 16396 9920
rect 16448 9868 16454 9920
rect 17954 9868 17960 9920
rect 18012 9868 18018 9920
rect 19426 9868 19432 9920
rect 19484 9908 19490 9920
rect 20441 9911 20499 9917
rect 20441 9908 20453 9911
rect 19484 9880 20453 9908
rect 19484 9868 19490 9880
rect 20441 9877 20453 9880
rect 20487 9877 20499 9911
rect 20441 9871 20499 9877
rect 552 9818 31372 9840
rect 552 9766 4250 9818
rect 4302 9766 4314 9818
rect 4366 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 11955 9818
rect 12007 9766 12019 9818
rect 12071 9766 12083 9818
rect 12135 9766 12147 9818
rect 12199 9766 12211 9818
rect 12263 9766 19660 9818
rect 19712 9766 19724 9818
rect 19776 9766 19788 9818
rect 19840 9766 19852 9818
rect 19904 9766 19916 9818
rect 19968 9766 27365 9818
rect 27417 9766 27429 9818
rect 27481 9766 27493 9818
rect 27545 9766 27557 9818
rect 27609 9766 27621 9818
rect 27673 9766 31372 9818
rect 552 9744 31372 9766
rect 9766 9704 9772 9716
rect 9140 9676 9772 9704
rect 8665 9639 8723 9645
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 9140 9636 9168 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 11238 9704 11244 9716
rect 10744 9676 11244 9704
rect 10744 9664 10750 9676
rect 11238 9664 11244 9676
rect 11296 9704 11302 9716
rect 11333 9707 11391 9713
rect 11333 9704 11345 9707
rect 11296 9676 11345 9704
rect 11296 9664 11302 9676
rect 11333 9673 11345 9676
rect 11379 9673 11391 9707
rect 11333 9667 11391 9673
rect 16390 9664 16396 9716
rect 16448 9664 16454 9716
rect 17586 9664 17592 9716
rect 17644 9664 17650 9716
rect 18049 9707 18107 9713
rect 18049 9673 18061 9707
rect 18095 9704 18107 9707
rect 18414 9704 18420 9716
rect 18095 9676 18420 9704
rect 18095 9673 18107 9676
rect 18049 9667 18107 9673
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 19576 9676 20668 9704
rect 19576 9664 19582 9676
rect 8711 9608 9168 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 10134 9596 10140 9648
rect 10192 9636 10198 9648
rect 10873 9639 10931 9645
rect 10873 9636 10885 9639
rect 10192 9608 10885 9636
rect 10192 9596 10198 9608
rect 10873 9605 10885 9608
rect 10919 9605 10931 9639
rect 10873 9599 10931 9605
rect 13909 9639 13967 9645
rect 13909 9605 13921 9639
rect 13955 9636 13967 9639
rect 16574 9636 16580 9648
rect 13955 9608 16580 9636
rect 13955 9605 13967 9608
rect 13909 9599 13967 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 11514 9568 11520 9580
rect 9048 9540 9260 9568
rect 8202 9460 8208 9512
rect 8260 9460 8266 9512
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8812 9472 8861 9500
rect 8812 9460 8818 9472
rect 8849 9469 8861 9472
rect 8895 9500 8907 9503
rect 9048 9500 9076 9540
rect 8895 9472 9076 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 9232 9500 9260 9540
rect 10336 9540 11520 9568
rect 9398 9509 9404 9512
rect 9232 9472 9352 9500
rect 8113 9435 8171 9441
rect 8113 9401 8125 9435
rect 8159 9432 8171 9435
rect 9214 9432 9220 9444
rect 8159 9404 9220 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 9214 9392 9220 9404
rect 9272 9392 9278 9444
rect 9324 9432 9352 9472
rect 9392 9463 9404 9509
rect 9456 9500 9462 9512
rect 10336 9500 10364 9540
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 15286 9568 15292 9580
rect 13556 9540 15292 9568
rect 11330 9500 11336 9512
rect 9456 9472 9492 9500
rect 9646 9472 10364 9500
rect 10428 9472 11336 9500
rect 9398 9460 9404 9463
rect 9456 9460 9462 9472
rect 9646 9432 9674 9472
rect 9324 9404 9674 9432
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 10428 9364 10456 9472
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9500 11483 9503
rect 11606 9500 11612 9512
rect 11471 9472 11612 9500
rect 11471 9469 11483 9472
rect 11425 9463 11483 9469
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 13556 9509 13584 9540
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 17604 9568 17632 9664
rect 18506 9596 18512 9648
rect 18564 9636 18570 9648
rect 18969 9639 19027 9645
rect 18969 9636 18981 9639
rect 18564 9608 18981 9636
rect 18564 9596 18570 9608
rect 18969 9605 18981 9608
rect 19015 9605 19027 9639
rect 18969 9599 19027 9605
rect 19058 9596 19064 9648
rect 19116 9636 19122 9648
rect 19889 9639 19947 9645
rect 19889 9636 19901 9639
rect 19116 9608 19901 9636
rect 19116 9596 19122 9608
rect 19889 9605 19901 9608
rect 19935 9605 19947 9639
rect 19889 9599 19947 9605
rect 16224 9540 17632 9568
rect 13722 9509 13728 9512
rect 13556 9503 13634 9509
rect 13556 9472 13588 9503
rect 13576 9469 13588 9472
rect 13622 9469 13634 9503
rect 13576 9463 13634 9469
rect 13679 9503 13728 9509
rect 13679 9469 13691 9503
rect 13725 9469 13728 9503
rect 13679 9463 13728 9469
rect 13722 9460 13728 9463
rect 13780 9460 13786 9512
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 13998 9500 14004 9512
rect 13863 9472 14004 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9500 14151 9503
rect 14366 9500 14372 9512
rect 14139 9472 14372 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 16224 9509 16252 9540
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 17920 9540 19564 9568
rect 17920 9528 17926 9540
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 16482 9460 16488 9512
rect 16540 9460 16546 9512
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 19536 9509 19564 9540
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 17184 9472 19257 9500
rect 17184 9460 17190 9472
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 19245 9463 19303 9469
rect 19352 9472 19441 9500
rect 10689 9435 10747 9441
rect 10689 9432 10701 9435
rect 10520 9404 10701 9432
rect 10520 9373 10548 9404
rect 10689 9401 10701 9404
rect 10735 9401 10747 9435
rect 10689 9395 10747 9401
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 16577 9435 16635 9441
rect 16577 9432 16589 9435
rect 13320 9404 16589 9432
rect 13320 9392 13326 9404
rect 16577 9401 16589 9404
rect 16623 9401 16635 9435
rect 16577 9395 16635 9401
rect 17954 9392 17960 9444
rect 18012 9432 18018 9444
rect 18785 9435 18843 9441
rect 18785 9432 18797 9435
rect 18012 9404 18797 9432
rect 18012 9392 18018 9404
rect 18785 9401 18797 9404
rect 18831 9401 18843 9435
rect 19352 9432 19380 9472
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19613 9503 19671 9509
rect 19613 9469 19625 9503
rect 19659 9500 19671 9503
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19659 9472 19809 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 20257 9503 20315 9509
rect 20257 9469 20269 9503
rect 20303 9500 20315 9503
rect 20441 9503 20499 9509
rect 20441 9500 20453 9503
rect 20303 9472 20453 9500
rect 20303 9469 20315 9472
rect 20257 9463 20315 9469
rect 20441 9469 20453 9472
rect 20487 9469 20499 9503
rect 20441 9463 20499 9469
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 20640 9509 20668 9676
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 18785 9395 18843 9401
rect 18892 9404 19380 9432
rect 8904 9336 10456 9364
rect 10505 9367 10563 9373
rect 8904 9324 8910 9336
rect 10505 9333 10517 9367
rect 10551 9333 10563 9367
rect 10505 9327 10563 9333
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12434 9364 12440 9376
rect 12023 9336 12440 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 15378 9324 15384 9376
rect 15436 9324 15442 9376
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 17218 9364 17224 9376
rect 16163 9336 17224 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 17218 9324 17224 9336
rect 17276 9364 17282 9376
rect 17494 9364 17500 9376
rect 17276 9336 17500 9364
rect 17276 9324 17282 9336
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 18892 9364 18920 9404
rect 17736 9336 18920 9364
rect 17736 9324 17742 9336
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 19024 9336 19257 9364
rect 19024 9324 19030 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 20165 9367 20223 9373
rect 20165 9333 20177 9367
rect 20211 9364 20223 9367
rect 20717 9367 20775 9373
rect 20717 9364 20729 9367
rect 20211 9336 20729 9364
rect 20211 9333 20223 9336
rect 20165 9327 20223 9333
rect 20717 9333 20729 9336
rect 20763 9333 20775 9367
rect 20717 9327 20775 9333
rect 552 9274 31531 9296
rect 552 9222 8102 9274
rect 8154 9222 8166 9274
rect 8218 9222 8230 9274
rect 8282 9222 8294 9274
rect 8346 9222 8358 9274
rect 8410 9222 15807 9274
rect 15859 9222 15871 9274
rect 15923 9222 15935 9274
rect 15987 9222 15999 9274
rect 16051 9222 16063 9274
rect 16115 9222 23512 9274
rect 23564 9222 23576 9274
rect 23628 9222 23640 9274
rect 23692 9222 23704 9274
rect 23756 9222 23768 9274
rect 23820 9222 31217 9274
rect 31269 9222 31281 9274
rect 31333 9222 31345 9274
rect 31397 9222 31409 9274
rect 31461 9222 31473 9274
rect 31525 9222 31531 9274
rect 552 9200 31531 9222
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 9306 9160 9312 9172
rect 8435 9132 9312 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 10778 9120 10784 9172
rect 10836 9120 10842 9172
rect 10870 9120 10876 9172
rect 10928 9120 10934 9172
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 11882 9160 11888 9172
rect 11572 9132 11888 9160
rect 11572 9120 11578 9132
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 15197 9163 15255 9169
rect 15197 9160 15209 9163
rect 13320 9132 15209 9160
rect 13320 9120 13326 9132
rect 15197 9129 15209 9132
rect 15243 9129 15255 9163
rect 15197 9123 15255 9129
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 15712 9132 15853 9160
rect 15712 9120 15718 9132
rect 15841 9129 15853 9132
rect 15887 9129 15899 9163
rect 15841 9123 15899 9129
rect 16209 9163 16267 9169
rect 16209 9129 16221 9163
rect 16255 9160 16267 9163
rect 16298 9160 16304 9172
rect 16255 9132 16304 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 19613 9163 19671 9169
rect 19613 9129 19625 9163
rect 19659 9160 19671 9163
rect 20073 9163 20131 9169
rect 19659 9132 19840 9160
rect 19659 9129 19671 9132
rect 19613 9123 19671 9129
rect 10796 9092 10824 9120
rect 8404 9064 10824 9092
rect 10888 9092 10916 9120
rect 11977 9095 12035 9101
rect 11977 9092 11989 9095
rect 10888 9064 11989 9092
rect 7837 9027 7895 9033
rect 7837 8993 7849 9027
rect 7883 9024 7895 9027
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 7883 8996 7941 9024
rect 7883 8993 7895 8996
rect 7837 8987 7895 8993
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 7944 8956 7972 8987
rect 8202 8984 8208 9036
rect 8260 8984 8266 9036
rect 8404 9033 8432 9064
rect 11977 9061 11989 9064
rect 12023 9061 12035 9095
rect 11977 9055 12035 9061
rect 13633 9095 13691 9101
rect 13633 9061 13645 9095
rect 13679 9092 13691 9095
rect 15378 9092 15384 9104
rect 13679 9064 15384 9092
rect 13679 9061 13691 9064
rect 13633 9055 13691 9061
rect 15378 9052 15384 9064
rect 15436 9092 15442 9104
rect 16393 9095 16451 9101
rect 16393 9092 16405 9095
rect 15436 9064 16405 9092
rect 15436 9052 15442 9064
rect 16393 9061 16405 9064
rect 16439 9061 16451 9095
rect 16393 9055 16451 9061
rect 18500 9095 18558 9101
rect 18500 9061 18512 9095
rect 18546 9092 18558 9095
rect 19426 9092 19432 9104
rect 18546 9064 19432 9092
rect 18546 9061 18558 9064
rect 18500 9055 18558 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 19812 9101 19840 9132
rect 20073 9129 20085 9163
rect 20119 9160 20131 9163
rect 28258 9160 28264 9172
rect 20119 9132 28264 9160
rect 20119 9129 20131 9132
rect 20073 9123 20131 9129
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 19797 9095 19855 9101
rect 19797 9061 19809 9095
rect 19843 9061 19855 9095
rect 19797 9055 19855 9061
rect 19904 9064 21588 9092
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 8665 9027 8723 9033
rect 8665 8993 8677 9027
rect 8711 9024 8723 9027
rect 8754 9024 8760 9036
rect 8711 8996 8760 9024
rect 8711 8993 8723 8996
rect 8665 8987 8723 8993
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 8846 8984 8852 9036
rect 8904 8984 8910 9036
rect 8938 8984 8944 9036
rect 8996 8984 9002 9036
rect 9033 9027 9091 9033
rect 9033 8993 9045 9027
rect 9079 9024 9091 9027
rect 9122 9024 9128 9036
rect 9079 8996 9128 9024
rect 9079 8993 9091 8996
rect 9033 8987 9091 8993
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 9306 9033 9312 9036
rect 9300 9024 9312 9033
rect 9267 8996 9312 9024
rect 9300 8987 9312 8996
rect 9306 8984 9312 8987
rect 9364 8984 9370 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 10502 9024 10508 9036
rect 9732 8996 10508 9024
rect 9732 8984 9738 8996
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 10686 9024 10692 9036
rect 10643 8996 10692 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10796 8996 11069 9024
rect 8294 8956 8300 8968
rect 7944 8928 8300 8956
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 10796 8956 10824 8996
rect 11057 8993 11069 8996
rect 11103 8993 11115 9027
rect 11057 8987 11115 8993
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11572 8996 11621 9024
rect 11572 8984 11578 8996
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 11756 8996 12434 9024
rect 11756 8984 11762 8996
rect 10428 8928 10824 8956
rect 10428 8897 10456 8928
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8888 7803 8891
rect 10413 8891 10471 8897
rect 7791 8860 9076 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 8754 8820 8760 8832
rect 8619 8792 8760 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9048 8820 9076 8860
rect 10413 8857 10425 8891
rect 10459 8857 10471 8891
rect 10413 8851 10471 8857
rect 10689 8891 10747 8897
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 11238 8888 11244 8900
rect 10735 8860 11244 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 12406 8888 12434 8996
rect 13906 8984 13912 9036
rect 13964 8984 13970 9036
rect 15654 8984 15660 9036
rect 15712 8984 15718 9036
rect 15746 8984 15752 9036
rect 15804 9024 15810 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15804 8996 15945 9024
rect 15804 8984 15810 8996
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 13630 8956 13636 8968
rect 12584 8928 13636 8956
rect 12584 8916 12590 8928
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 15672 8956 15700 8984
rect 16132 8956 16160 8987
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 16908 8996 18245 9024
rect 16908 8984 16914 8996
rect 18233 8993 18245 8996
rect 18279 9024 18291 9027
rect 18322 9024 18328 9036
rect 18279 8996 18328 9024
rect 18279 8993 18291 8996
rect 18233 8987 18291 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 19904 9024 19932 9064
rect 19576 8996 19932 9024
rect 19576 8984 19582 8996
rect 20346 8984 20352 9036
rect 20404 8984 20410 9036
rect 20530 8984 20536 9036
rect 20588 9024 20594 9036
rect 20809 9027 20867 9033
rect 20809 9024 20821 9027
rect 20588 8996 20821 9024
rect 20588 8984 20594 8996
rect 20809 8993 20821 8996
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 21560 9033 21588 9064
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20956 8996 21281 9024
rect 20956 8984 20962 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 21545 9027 21603 9033
rect 21545 8993 21557 9027
rect 21591 8993 21603 9027
rect 21545 8987 21603 8993
rect 15672 8928 16160 8956
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 17862 8956 17868 8968
rect 16632 8928 17868 8956
rect 16632 8916 16638 8928
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 20438 8916 20444 8968
rect 20496 8956 20502 8968
rect 21637 8959 21695 8965
rect 21637 8956 21649 8959
rect 20496 8928 21649 8956
rect 20496 8916 20502 8928
rect 21637 8925 21649 8928
rect 21683 8925 21695 8959
rect 21637 8919 21695 8925
rect 13078 8888 13084 8900
rect 11532 8860 12296 8888
rect 12406 8860 13084 8888
rect 11532 8832 11560 8860
rect 9674 8820 9680 8832
rect 9048 8792 9680 8820
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 11054 8820 11060 8832
rect 9824 8792 11060 8820
rect 9824 8780 9830 8792
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 11514 8780 11520 8832
rect 11572 8780 11578 8832
rect 11698 8780 11704 8832
rect 11756 8780 11762 8832
rect 12268 8820 12296 8860
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13998 8888 14004 8900
rect 13188 8860 14004 8888
rect 12618 8820 12624 8832
rect 12268 8792 12624 8820
rect 12618 8780 12624 8792
rect 12676 8820 12682 8832
rect 13188 8820 13216 8860
rect 13998 8848 14004 8860
rect 14056 8848 14062 8900
rect 20625 8891 20683 8897
rect 20625 8857 20637 8891
rect 20671 8888 20683 8891
rect 28258 8888 28264 8900
rect 20671 8860 28264 8888
rect 20671 8857 20683 8860
rect 20625 8851 20683 8857
rect 28258 8848 28264 8860
rect 28316 8848 28322 8900
rect 12676 8792 13216 8820
rect 12676 8780 12682 8792
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 14642 8820 14648 8832
rect 13320 8792 14648 8820
rect 13320 8780 13326 8792
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 17034 8780 17040 8832
rect 17092 8820 17098 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17092 8792 17693 8820
rect 17092 8780 17098 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 17681 8783 17739 8789
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 19978 8820 19984 8832
rect 18012 8792 19984 8820
rect 18012 8780 18018 8792
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 20901 8823 20959 8829
rect 20901 8820 20913 8823
rect 20588 8792 20913 8820
rect 20588 8780 20594 8792
rect 20901 8789 20913 8792
rect 20947 8789 20959 8823
rect 20901 8783 20959 8789
rect 21358 8780 21364 8832
rect 21416 8780 21422 8832
rect 552 8730 31372 8752
rect 552 8678 4250 8730
rect 4302 8678 4314 8730
rect 4366 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 11955 8730
rect 12007 8678 12019 8730
rect 12071 8678 12083 8730
rect 12135 8678 12147 8730
rect 12199 8678 12211 8730
rect 12263 8678 19660 8730
rect 19712 8678 19724 8730
rect 19776 8678 19788 8730
rect 19840 8678 19852 8730
rect 19904 8678 19916 8730
rect 19968 8678 27365 8730
rect 27417 8678 27429 8730
rect 27481 8678 27493 8730
rect 27545 8678 27557 8730
rect 27609 8678 27621 8730
rect 27673 8678 31372 8730
rect 552 8656 31372 8678
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 9306 8616 9312 8628
rect 8076 8588 9312 8616
rect 8076 8576 8082 8588
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9416 8588 9812 8616
rect 9416 8548 9444 8588
rect 8956 8520 9444 8548
rect 9784 8548 9812 8588
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 9916 8588 10241 8616
rect 9916 8576 9922 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 11146 8616 11152 8628
rect 10551 8588 11152 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8616 11391 8619
rect 11606 8616 11612 8628
rect 11379 8588 11612 8616
rect 11379 8585 11391 8588
rect 11333 8579 11391 8585
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 13814 8616 13820 8628
rect 13136 8588 13820 8616
rect 13136 8576 13142 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 17126 8576 17132 8628
rect 17184 8576 17190 8628
rect 17405 8619 17463 8625
rect 17405 8585 17417 8619
rect 17451 8616 17463 8619
rect 18966 8616 18972 8628
rect 17451 8588 18972 8616
rect 17451 8585 17463 8588
rect 17405 8579 17463 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8616 20131 8619
rect 20346 8616 20352 8628
rect 20119 8588 20352 8616
rect 20119 8585 20131 8588
rect 20073 8579 20131 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 10778 8548 10784 8560
rect 9784 8520 10784 8548
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8846 8480 8852 8492
rect 8159 8452 8852 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8386 8412 8392 8424
rect 8251 8384 8392 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8381 8539 8415
rect 8481 8375 8539 8381
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 8496 8344 8524 8375
rect 8662 8372 8668 8424
rect 8720 8372 8726 8424
rect 8956 8421 8984 8520
rect 10778 8508 10784 8520
rect 10836 8508 10842 8560
rect 11057 8551 11115 8557
rect 11057 8517 11069 8551
rect 11103 8548 11115 8551
rect 11103 8520 11652 8548
rect 11103 8517 11115 8520
rect 11057 8511 11115 8517
rect 11624 8492 11652 8520
rect 11698 8508 11704 8560
rect 11756 8508 11762 8560
rect 12161 8551 12219 8557
rect 12161 8517 12173 8551
rect 12207 8548 12219 8551
rect 12802 8548 12808 8560
rect 12207 8520 12808 8548
rect 12207 8517 12219 8520
rect 12161 8511 12219 8517
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 13262 8508 13268 8560
rect 13320 8508 13326 8560
rect 17678 8508 17684 8560
rect 17736 8508 17742 8560
rect 17957 8551 18015 8557
rect 17957 8517 17969 8551
rect 18003 8548 18015 8551
rect 18046 8548 18052 8560
rect 18003 8520 18052 8548
rect 18003 8517 18015 8520
rect 17957 8511 18015 8517
rect 18046 8508 18052 8520
rect 18104 8508 18110 8560
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 18196 8520 18245 8548
rect 18196 8508 18202 8520
rect 18233 8517 18245 8520
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9398 8480 9404 8492
rect 9171 8452 9404 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 10134 8480 10140 8492
rect 9646 8452 10140 8480
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 9079 8384 9321 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 8076 8316 8524 8344
rect 8076 8304 8082 8316
rect 8570 8304 8576 8356
rect 8628 8304 8634 8356
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8849 8279 8907 8285
rect 8849 8276 8861 8279
rect 8352 8248 8861 8276
rect 8352 8236 8358 8248
rect 8849 8245 8861 8248
rect 8895 8276 8907 8279
rect 9030 8276 9036 8288
rect 8895 8248 9036 8276
rect 8895 8245 8907 8248
rect 8849 8239 8907 8245
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 9324 8276 9352 8375
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9646 8412 9674 8452
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10870 8480 10876 8492
rect 10336 8452 10876 8480
rect 10336 8424 10364 8452
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 11514 8480 11520 8492
rect 11164 8452 11520 8480
rect 9548 8384 9674 8412
rect 9548 8372 9554 8384
rect 9766 8372 9772 8424
rect 9824 8372 9830 8424
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 10226 8412 10232 8424
rect 10091 8384 10232 8412
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10318 8372 10324 8424
rect 10376 8372 10382 8424
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 10502 8412 10508 8424
rect 10459 8384 10508 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 11164 8421 11192 8452
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11606 8440 11612 8492
rect 11664 8440 11670 8492
rect 11716 8480 11744 8508
rect 11716 8452 11836 8480
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10652 8384 10701 8412
rect 10652 8372 10658 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8381 11299 8415
rect 11241 8375 11299 8381
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8412 11759 8415
rect 11808 8412 11836 8452
rect 11747 8384 11836 8412
rect 11900 8452 13492 8480
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 9398 8304 9404 8356
rect 9456 8304 9462 8356
rect 9677 8347 9735 8353
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 10962 8344 10968 8356
rect 9723 8316 10968 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 9766 8276 9772 8288
rect 9324 8248 9772 8276
rect 9766 8236 9772 8248
rect 9824 8236 9830 8288
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 10781 8279 10839 8285
rect 10781 8276 10793 8279
rect 10468 8248 10793 8276
rect 10468 8236 10474 8248
rect 10781 8245 10793 8248
rect 10827 8245 10839 8279
rect 10781 8239 10839 8245
rect 10870 8236 10876 8288
rect 10928 8276 10934 8288
rect 11256 8276 11284 8375
rect 11609 8347 11667 8353
rect 11609 8313 11621 8347
rect 11655 8344 11667 8347
rect 11900 8344 11928 8452
rect 11974 8372 11980 8424
rect 12032 8372 12038 8424
rect 12069 8415 12127 8421
rect 12069 8381 12081 8415
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 11655 8316 11928 8344
rect 11655 8313 11667 8316
rect 11609 8307 11667 8313
rect 12084 8288 12112 8375
rect 12526 8372 12532 8424
rect 12584 8372 12590 8424
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12676 8384 13001 8412
rect 12676 8372 12682 8384
rect 12989 8381 13001 8384
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 13078 8372 13084 8424
rect 13136 8372 13142 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 13280 8384 13369 8412
rect 11790 8276 11796 8288
rect 10928 8248 11796 8276
rect 10928 8236 10934 8248
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 11882 8236 11888 8288
rect 11940 8236 11946 8288
rect 12066 8236 12072 8288
rect 12124 8236 12130 8288
rect 12437 8279 12495 8285
rect 12437 8245 12449 8279
rect 12483 8276 12495 8279
rect 12618 8276 12624 8288
rect 12483 8248 12624 8276
rect 12483 8245 12495 8248
rect 12437 8239 12495 8245
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 12894 8276 12900 8288
rect 12759 8248 12900 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 13280 8276 13308 8384
rect 13357 8381 13369 8384
rect 13403 8381 13415 8415
rect 13464 8412 13492 8452
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 15010 8440 15016 8492
rect 15068 8480 15074 8492
rect 15286 8480 15292 8492
rect 15068 8452 15292 8480
rect 15068 8440 15074 8452
rect 15286 8440 15292 8452
rect 15344 8480 15350 8492
rect 16850 8480 16856 8492
rect 15344 8452 16856 8480
rect 15344 8440 15350 8452
rect 15856 8421 15884 8452
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 18322 8440 18328 8492
rect 18380 8480 18386 8492
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 18380 8452 18705 8480
rect 18380 8440 18386 8452
rect 18693 8449 18705 8452
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 19978 8440 19984 8492
rect 20036 8480 20042 8492
rect 20036 8452 20484 8480
rect 20036 8440 20042 8452
rect 16945 8425 17003 8431
rect 16945 8424 16957 8425
rect 16991 8424 17003 8425
rect 13797 8415 13855 8421
rect 13797 8412 13809 8415
rect 13464 8384 13809 8412
rect 13357 8375 13415 8381
rect 13797 8381 13809 8384
rect 13843 8381 13855 8415
rect 15841 8415 15899 8421
rect 13797 8375 13855 8381
rect 14292 8384 15792 8412
rect 14292 8356 14320 8384
rect 14274 8304 14280 8356
rect 14332 8304 14338 8356
rect 15105 8347 15163 8353
rect 15105 8344 15117 8347
rect 14936 8316 15117 8344
rect 14366 8276 14372 8288
rect 13280 8248 14372 8276
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 14936 8285 14964 8316
rect 15105 8313 15117 8316
rect 15151 8313 15163 8347
rect 15764 8344 15792 8384
rect 15841 8381 15853 8415
rect 15887 8381 15899 8415
rect 15841 8375 15899 8381
rect 16117 8415 16175 8421
rect 16117 8381 16129 8415
rect 16163 8412 16175 8415
rect 16206 8412 16212 8424
rect 16163 8384 16212 8412
rect 16163 8381 16175 8384
rect 16117 8375 16175 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 16393 8415 16451 8421
rect 16393 8381 16405 8415
rect 16439 8412 16451 8415
rect 16574 8412 16580 8424
rect 16439 8384 16580 8412
rect 16439 8381 16451 8384
rect 16393 8375 16451 8381
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 16669 8415 16727 8421
rect 16669 8381 16681 8415
rect 16715 8381 16727 8415
rect 16942 8412 16948 8424
rect 16913 8384 16948 8412
rect 16669 8375 16727 8381
rect 16684 8344 16712 8375
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17037 8415 17095 8421
rect 17037 8381 17049 8415
rect 17083 8412 17095 8415
rect 17313 8415 17371 8421
rect 17083 8384 17163 8412
rect 17083 8381 17095 8384
rect 17037 8375 17095 8381
rect 17135 8356 17163 8384
rect 17313 8381 17325 8415
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 17126 8344 17132 8356
rect 15764 8316 17132 8344
rect 15105 8307 15163 8313
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 17328 8344 17356 8375
rect 17770 8372 17776 8424
rect 17828 8372 17834 8424
rect 17862 8372 17868 8424
rect 17920 8372 17926 8424
rect 18141 8415 18199 8421
rect 18141 8381 18153 8415
rect 18187 8412 18199 8415
rect 18230 8412 18236 8424
rect 18187 8384 18236 8412
rect 18187 8381 18199 8384
rect 18141 8375 18199 8381
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 20456 8421 20484 8452
rect 20165 8415 20223 8421
rect 20165 8412 20177 8415
rect 18800 8384 20177 8412
rect 17276 8316 17356 8344
rect 17276 8304 17282 8316
rect 17402 8304 17408 8356
rect 17460 8344 17466 8356
rect 18800 8344 18828 8384
rect 20165 8381 20177 8384
rect 20211 8381 20223 8415
rect 20165 8375 20223 8381
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8381 20407 8415
rect 20349 8375 20407 8381
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8381 20499 8415
rect 20441 8375 20499 8381
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8412 20591 8415
rect 20717 8415 20775 8421
rect 20717 8412 20729 8415
rect 20579 8384 20729 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20717 8381 20729 8384
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 17460 8316 18828 8344
rect 18960 8347 19018 8353
rect 17460 8304 17466 8316
rect 18960 8313 18972 8347
rect 19006 8344 19018 8347
rect 19426 8344 19432 8356
rect 19006 8316 19432 8344
rect 19006 8313 19018 8316
rect 18960 8307 19018 8313
rect 19426 8304 19432 8316
rect 19484 8304 19490 8356
rect 20254 8304 20260 8356
rect 20312 8304 20318 8356
rect 14921 8279 14979 8285
rect 14921 8245 14933 8279
rect 14967 8245 14979 8279
rect 14921 8239 14979 8245
rect 15194 8236 15200 8288
rect 15252 8236 15258 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 16025 8279 16083 8285
rect 16025 8276 16037 8279
rect 15712 8248 16037 8276
rect 15712 8236 15718 8248
rect 16025 8245 16037 8248
rect 16071 8245 16083 8279
rect 16025 8239 16083 8245
rect 16298 8236 16304 8288
rect 16356 8236 16362 8288
rect 16574 8236 16580 8288
rect 16632 8236 16638 8288
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 16853 8279 16911 8285
rect 16853 8276 16865 8279
rect 16724 8248 16865 8276
rect 16724 8236 16730 8248
rect 16853 8245 16865 8248
rect 16899 8245 16911 8279
rect 16853 8239 16911 8245
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 20364 8276 20392 8375
rect 19392 8248 20392 8276
rect 19392 8236 19398 8248
rect 20806 8236 20812 8288
rect 20864 8236 20870 8288
rect 552 8186 31531 8208
rect 552 8134 8102 8186
rect 8154 8134 8166 8186
rect 8218 8134 8230 8186
rect 8282 8134 8294 8186
rect 8346 8134 8358 8186
rect 8410 8134 15807 8186
rect 15859 8134 15871 8186
rect 15923 8134 15935 8186
rect 15987 8134 15999 8186
rect 16051 8134 16063 8186
rect 16115 8134 23512 8186
rect 23564 8134 23576 8186
rect 23628 8134 23640 8186
rect 23692 8134 23704 8186
rect 23756 8134 23768 8186
rect 23820 8134 31217 8186
rect 31269 8134 31281 8186
rect 31333 8134 31345 8186
rect 31397 8134 31409 8186
rect 31461 8134 31473 8186
rect 31525 8134 31531 8186
rect 552 8112 31531 8134
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 8536 8044 8677 8072
rect 8536 8032 8542 8044
rect 8665 8041 8677 8044
rect 8711 8041 8723 8075
rect 9030 8072 9036 8084
rect 8665 8035 8723 8041
rect 8772 8044 9036 8072
rect 8772 7945 8800 8044
rect 9030 8032 9036 8044
rect 9088 8072 9094 8084
rect 10505 8075 10563 8081
rect 9088 8044 9628 8072
rect 9088 8032 9094 8044
rect 9600 8016 9628 8044
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 10551 8044 11100 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 8846 7964 8852 8016
rect 8904 8004 8910 8016
rect 9370 8007 9428 8013
rect 9370 8004 9382 8007
rect 8904 7976 9382 8004
rect 8904 7964 8910 7976
rect 9370 7973 9382 7976
rect 9416 7973 9428 8007
rect 9370 7967 9428 7973
rect 9582 7964 9588 8016
rect 9640 7964 9646 8016
rect 9766 8004 9772 8016
rect 9692 7976 9772 8004
rect 8757 7939 8815 7945
rect 8757 7905 8769 7939
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 9033 7939 9091 7945
rect 9033 7905 9045 7939
rect 9079 7936 9091 7939
rect 9692 7936 9720 7976
rect 9766 7964 9772 7976
rect 9824 8004 9830 8016
rect 10686 8004 10692 8016
rect 9824 7976 10692 8004
rect 9824 7964 9830 7976
rect 10686 7964 10692 7976
rect 10744 8004 10750 8016
rect 10870 8004 10876 8016
rect 10744 7976 10876 8004
rect 10744 7964 10750 7976
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 11072 8013 11100 8044
rect 11146 8032 11152 8084
rect 11204 8032 11210 8084
rect 11238 8032 11244 8084
rect 11296 8032 11302 8084
rect 11422 8032 11428 8084
rect 11480 8032 11486 8084
rect 11882 8032 11888 8084
rect 11940 8032 11946 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 13446 8072 13452 8084
rect 12124 8044 13452 8072
rect 12124 8032 12130 8044
rect 11057 8007 11115 8013
rect 11057 7973 11069 8007
rect 11103 7973 11115 8007
rect 11057 7967 11115 7973
rect 9079 7908 9720 7936
rect 9079 7905 9091 7908
rect 9033 7899 9091 7905
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10502 7936 10508 7948
rect 10008 7908 10508 7936
rect 10008 7896 10014 7908
rect 10502 7896 10508 7908
rect 10560 7936 10566 7948
rect 10597 7939 10655 7945
rect 10597 7936 10609 7939
rect 10560 7908 10609 7936
rect 10560 7896 10566 7908
rect 10597 7905 10609 7908
rect 10643 7936 10655 7939
rect 10962 7936 10968 7948
rect 10643 7908 10968 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11256 7936 11284 8032
rect 11440 8004 11468 8032
rect 11900 8004 11928 8032
rect 11440 7976 11836 8004
rect 11900 7976 12388 8004
rect 11808 7945 11836 7976
rect 12360 7945 12388 7976
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 11256 7908 11529 7936
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 12253 7939 12311 7945
rect 12253 7905 12265 7939
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7905 12587 7939
rect 12728 7936 12756 8044
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13679 8044 14105 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14366 8032 14372 8084
rect 14424 8032 14430 8084
rect 14642 8032 14648 8084
rect 14700 8032 14706 8084
rect 15562 8072 15568 8084
rect 14752 8044 15568 8072
rect 12894 7964 12900 8016
rect 12952 7964 12958 8016
rect 13372 7976 13584 8004
rect 12797 7939 12855 7945
rect 12797 7936 12809 7939
rect 12728 7908 12809 7936
rect 12529 7899 12587 7905
rect 12797 7905 12809 7908
rect 12843 7905 12855 7939
rect 12912 7935 12940 7964
rect 13372 7945 13400 7976
rect 13357 7939 13415 7945
rect 12797 7899 12855 7905
rect 12889 7929 12947 7935
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 11422 7868 11428 7880
rect 10376 7840 11428 7868
rect 10376 7828 10382 7840
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 12268 7868 12296 7899
rect 12434 7868 12440 7880
rect 12268 7840 12440 7868
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 12544 7868 12572 7899
rect 12889 7895 12901 7929
rect 12935 7895 12947 7929
rect 13357 7905 13369 7939
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 12889 7889 12947 7895
rect 12544 7840 12664 7868
rect 12066 7800 12072 7812
rect 10888 7772 12072 7800
rect 10888 7744 10916 7772
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 12526 7800 12532 7812
rect 12308 7772 12532 7800
rect 12308 7760 12314 7772
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 12636 7800 12664 7840
rect 12989 7803 13047 7809
rect 12989 7800 13001 7803
rect 12636 7772 13001 7800
rect 12989 7769 13001 7772
rect 13035 7769 13047 7803
rect 12989 7763 13047 7769
rect 8941 7735 8999 7741
rect 8941 7701 8953 7735
rect 8987 7732 8999 7735
rect 9766 7732 9772 7744
rect 8987 7704 9772 7732
rect 8987 7701 8999 7704
rect 8941 7695 8999 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10686 7692 10692 7744
rect 10744 7692 10750 7744
rect 10870 7692 10876 7744
rect 10928 7692 10934 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11606 7732 11612 7744
rect 11020 7704 11612 7732
rect 11020 7692 11026 7704
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 11885 7735 11943 7741
rect 11885 7701 11897 7735
rect 11931 7732 11943 7735
rect 12342 7732 12348 7744
rect 11931 7704 12348 7732
rect 11931 7701 11943 7704
rect 11885 7695 11943 7701
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7732 12495 7735
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 12483 7704 12725 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 12713 7695 12771 7701
rect 13262 7692 13268 7744
rect 13320 7692 13326 7744
rect 13464 7732 13492 7899
rect 13556 7800 13584 7976
rect 13814 7964 13820 8016
rect 13872 7964 13878 8016
rect 13998 7964 14004 8016
rect 14056 8004 14062 8016
rect 14056 7976 14504 8004
rect 14056 7964 14062 7976
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 13909 7939 13967 7945
rect 13909 7905 13921 7939
rect 13955 7936 13967 7939
rect 14090 7936 14096 7948
rect 13955 7908 14096 7936
rect 13955 7905 13967 7908
rect 13909 7899 13967 7905
rect 13648 7868 13676 7899
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14182 7896 14188 7948
rect 14240 7896 14246 7948
rect 14366 7896 14372 7948
rect 14424 7936 14430 7948
rect 14476 7945 14504 7976
rect 14752 7945 14780 8044
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 15654 8032 15660 8084
rect 15712 8032 15718 8084
rect 15841 8075 15899 8081
rect 15841 8041 15853 8075
rect 15887 8072 15899 8075
rect 16298 8072 16304 8084
rect 15887 8044 16304 8072
rect 15887 8041 15899 8044
rect 15841 8035 15899 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 16574 8032 16580 8084
rect 16632 8032 16638 8084
rect 17218 8072 17224 8084
rect 16776 8044 17224 8072
rect 15197 8007 15255 8013
rect 15197 8004 15209 8007
rect 15028 7976 15209 8004
rect 15028 7945 15056 7976
rect 15197 7973 15209 7976
rect 15243 7973 15255 8007
rect 15197 7967 15255 7973
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 14424 7908 14473 7936
rect 14424 7896 14430 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7905 14795 7939
rect 14737 7899 14795 7905
rect 15013 7939 15071 7945
rect 15013 7905 15025 7939
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 15102 7896 15108 7948
rect 15160 7936 15166 7948
rect 15672 7945 15700 8032
rect 16592 8004 16620 8032
rect 15856 7976 16620 8004
rect 15856 7945 15884 7976
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 15160 7908 15301 7936
rect 15160 7896 15166 7908
rect 15289 7905 15301 7908
rect 15335 7936 15347 7939
rect 15565 7939 15623 7945
rect 15335 7908 15516 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15488 7880 15516 7908
rect 15565 7905 15577 7939
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 15194 7868 15200 7880
rect 13648 7840 15200 7868
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 15580 7868 15608 7899
rect 16298 7896 16304 7948
rect 16356 7896 16362 7948
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 16776 7936 16804 8044
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 19705 8075 19763 8081
rect 19705 8041 19717 8075
rect 19751 8041 19763 8075
rect 19705 8035 19763 8041
rect 19720 8004 19748 8035
rect 19889 8007 19947 8013
rect 19889 8004 19901 8007
rect 16868 7976 18368 8004
rect 19720 7976 19901 8004
rect 16868 7948 16896 7976
rect 16623 7908 16804 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 16850 7896 16856 7948
rect 16908 7896 16914 7948
rect 18340 7945 18368 7976
rect 19889 7973 19901 7976
rect 19935 7973 19947 8007
rect 19889 7967 19947 7973
rect 17120 7939 17178 7945
rect 17120 7905 17132 7939
rect 17166 7936 17178 7939
rect 18325 7939 18383 7945
rect 17166 7908 18276 7936
rect 17166 7905 17178 7908
rect 17120 7899 17178 7905
rect 16666 7868 16672 7880
rect 15580 7840 16672 7868
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 17954 7828 17960 7880
rect 18012 7828 18018 7880
rect 18248 7868 18276 7908
rect 18325 7905 18337 7939
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 18592 7939 18650 7945
rect 18592 7905 18604 7939
rect 18638 7936 18650 7939
rect 18638 7908 19564 7936
rect 18638 7905 18650 7908
rect 18592 7899 18650 7905
rect 19536 7868 19564 7908
rect 20346 7896 20352 7948
rect 20404 7896 20410 7948
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 18248 7840 18368 7868
rect 19536 7840 20453 7868
rect 13998 7800 14004 7812
rect 13556 7772 14004 7800
rect 13998 7760 14004 7772
rect 14056 7760 14062 7812
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7800 14979 7803
rect 16209 7803 16267 7809
rect 16209 7800 16221 7803
rect 14967 7772 16221 7800
rect 14967 7769 14979 7772
rect 14921 7763 14979 7769
rect 16209 7769 16221 7772
rect 16255 7769 16267 7803
rect 16574 7800 16580 7812
rect 16209 7763 16267 7769
rect 16316 7772 16580 7800
rect 15378 7732 15384 7744
rect 13464 7704 15384 7732
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 15470 7692 15476 7744
rect 15528 7732 15534 7744
rect 16316 7732 16344 7772
rect 16574 7760 16580 7772
rect 16632 7800 16638 7812
rect 16632 7772 16804 7800
rect 16632 7760 16638 7772
rect 15528 7704 16344 7732
rect 15528 7692 15534 7704
rect 16666 7692 16672 7744
rect 16724 7692 16730 7744
rect 16776 7732 16804 7772
rect 17972 7732 18000 7828
rect 16776 7704 18000 7732
rect 18230 7692 18236 7744
rect 18288 7692 18294 7744
rect 18340 7732 18368 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 20806 7800 20812 7812
rect 19260 7772 20812 7800
rect 19260 7732 19288 7772
rect 20806 7760 20812 7772
rect 20864 7760 20870 7812
rect 18340 7704 19288 7732
rect 19978 7692 19984 7744
rect 20036 7692 20042 7744
rect 552 7642 31372 7664
rect 552 7590 4250 7642
rect 4302 7590 4314 7642
rect 4366 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 11955 7642
rect 12007 7590 12019 7642
rect 12071 7590 12083 7642
rect 12135 7590 12147 7642
rect 12199 7590 12211 7642
rect 12263 7590 19660 7642
rect 19712 7590 19724 7642
rect 19776 7590 19788 7642
rect 19840 7590 19852 7642
rect 19904 7590 19916 7642
rect 19968 7590 27365 7642
rect 27417 7590 27429 7642
rect 27481 7590 27493 7642
rect 27545 7590 27557 7642
rect 27609 7590 27621 7642
rect 27673 7590 31372 7642
rect 552 7568 31372 7590
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 11146 7528 11152 7540
rect 9999 7500 11152 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 12710 7528 12716 7540
rect 11296 7500 12716 7528
rect 11296 7488 11302 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 13262 7488 13268 7540
rect 13320 7488 13326 7540
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 15102 7528 15108 7540
rect 14240 7500 15108 7528
rect 14240 7488 14246 7500
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 16666 7488 16672 7540
rect 16724 7488 16730 7540
rect 18230 7488 18236 7540
rect 18288 7488 18294 7540
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 19334 7528 19340 7540
rect 18371 7500 19340 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19426 7488 19432 7540
rect 19484 7488 19490 7540
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7528 19671 7531
rect 20346 7528 20352 7540
rect 19659 7500 20352 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 9122 7420 9128 7472
rect 9180 7460 9186 7472
rect 10962 7460 10968 7472
rect 9180 7432 10968 7460
rect 9180 7420 9186 7432
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 12434 7420 12440 7472
rect 12492 7460 12498 7472
rect 13354 7460 13360 7472
rect 12492 7432 13360 7460
rect 12492 7420 12498 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 9950 7392 9956 7404
rect 9600 7364 9956 7392
rect 9600 7333 9628 7364
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 13538 7392 13544 7404
rect 10060 7364 11100 7392
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9858 7284 9864 7336
rect 9916 7284 9922 7336
rect 10060 7333 10088 7364
rect 11072 7336 11100 7364
rect 12406 7364 13544 7392
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 10226 7284 10232 7336
rect 10284 7284 10290 7336
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 10413 7327 10471 7333
rect 10413 7293 10425 7327
rect 10459 7324 10471 7327
rect 10459 7296 10548 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 9677 7259 9735 7265
rect 9677 7225 9689 7259
rect 9723 7256 9735 7259
rect 9950 7256 9956 7268
rect 9723 7228 9956 7256
rect 9723 7225 9735 7228
rect 9677 7219 9735 7225
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10336 7188 10364 7287
rect 10520 7256 10548 7296
rect 10870 7284 10876 7336
rect 10928 7284 10934 7336
rect 10962 7284 10968 7336
rect 11020 7284 11026 7336
rect 11054 7284 11060 7336
rect 11112 7284 11118 7336
rect 12406 7324 12434 7364
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 15010 7352 15016 7404
rect 15068 7392 15074 7404
rect 15381 7395 15439 7401
rect 15381 7392 15393 7395
rect 15068 7364 15393 7392
rect 15068 7352 15074 7364
rect 15381 7361 15393 7364
rect 15427 7361 15439 7395
rect 16684 7392 16712 7488
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 17000 7432 18000 7460
rect 17000 7420 17006 7432
rect 16684 7364 17724 7392
rect 15381 7355 15439 7361
rect 11164 7296 12434 7324
rect 10594 7256 10600 7268
rect 10520 7228 10600 7256
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 10980 7256 11008 7284
rect 11164 7256 11192 7296
rect 12618 7284 12624 7336
rect 12676 7284 12682 7336
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 12860 7296 13185 7324
rect 12860 7284 12866 7296
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 14090 7284 14096 7336
rect 14148 7324 14154 7336
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14148 7296 15117 7324
rect 14148 7284 14154 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 10980 7228 11192 7256
rect 11232 7259 11290 7265
rect 11232 7225 11244 7259
rect 11278 7256 11290 7259
rect 11330 7256 11336 7268
rect 11278 7228 11336 7256
rect 11278 7225 11290 7228
rect 11232 7219 11290 7225
rect 11330 7216 11336 7228
rect 11388 7216 11394 7268
rect 12529 7259 12587 7265
rect 12529 7256 12541 7259
rect 12360 7228 12541 7256
rect 10284 7160 10364 7188
rect 10284 7148 10290 7160
rect 10502 7148 10508 7200
rect 10560 7148 10566 7200
rect 10778 7148 10784 7200
rect 10836 7148 10842 7200
rect 12360 7197 12388 7228
rect 12529 7225 12541 7228
rect 12575 7225 12587 7259
rect 12636 7256 12664 7284
rect 13814 7265 13820 7268
rect 12636 7228 13768 7256
rect 12529 7219 12587 7225
rect 13740 7200 13768 7228
rect 13808 7219 13820 7265
rect 13814 7216 13820 7219
rect 13872 7216 13878 7268
rect 15120 7256 15148 7287
rect 17126 7284 17132 7336
rect 17184 7324 17190 7336
rect 17310 7324 17316 7336
rect 17184 7296 17316 7324
rect 17184 7284 17190 7296
rect 17310 7284 17316 7296
rect 17368 7324 17374 7336
rect 17696 7333 17724 7364
rect 17972 7333 18000 7432
rect 18248 7392 18276 7488
rect 19058 7420 19064 7472
rect 19116 7420 19122 7472
rect 19444 7460 19472 7488
rect 19889 7463 19947 7469
rect 19889 7460 19901 7463
rect 19444 7432 19901 7460
rect 19889 7429 19901 7432
rect 19935 7429 19947 7463
rect 19889 7423 19947 7429
rect 18248 7364 18828 7392
rect 18800 7333 18828 7364
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 17368 7296 17417 7324
rect 17368 7284 17374 7296
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 17681 7327 17739 7333
rect 17681 7293 17693 7327
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7324 18107 7327
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 18095 7296 18245 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18233 7293 18245 7296
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 18785 7327 18843 7333
rect 18785 7293 18797 7327
rect 18831 7293 18843 7327
rect 18785 7287 18843 7293
rect 19076 7324 19104 7420
rect 20622 7392 20628 7404
rect 19536 7364 20628 7392
rect 19245 7327 19303 7333
rect 19245 7324 19257 7327
rect 19076 7296 19257 7324
rect 15654 7265 15660 7268
rect 15120 7228 15516 7256
rect 12345 7191 12403 7197
rect 12345 7157 12357 7191
rect 12391 7157 12403 7191
rect 12345 7151 12403 7157
rect 12618 7148 12624 7200
rect 12676 7148 12682 7200
rect 13722 7148 13728 7200
rect 13780 7148 13786 7200
rect 14918 7148 14924 7200
rect 14976 7148 14982 7200
rect 15197 7191 15255 7197
rect 15197 7157 15209 7191
rect 15243 7188 15255 7191
rect 15378 7188 15384 7200
rect 15243 7160 15384 7188
rect 15243 7157 15255 7160
rect 15197 7151 15255 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 15488 7188 15516 7228
rect 15648 7219 15660 7265
rect 15654 7216 15660 7219
rect 15712 7216 15718 7268
rect 16666 7216 16672 7268
rect 16724 7216 16730 7268
rect 16945 7259 17003 7265
rect 16945 7225 16957 7259
rect 16991 7225 17003 7259
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 16945 7219 17003 7225
rect 17420 7228 17785 7256
rect 16684 7188 16712 7216
rect 15488 7160 16712 7188
rect 16761 7191 16819 7197
rect 16761 7157 16773 7191
rect 16807 7188 16819 7191
rect 16960 7188 16988 7219
rect 16807 7160 16988 7188
rect 16807 7157 16819 7160
rect 16761 7151 16819 7157
rect 17034 7148 17040 7200
rect 17092 7148 17098 7200
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 17420 7188 17448 7228
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 17972 7256 18000 7287
rect 18138 7256 18144 7268
rect 17972 7228 18144 7256
rect 17773 7219 17831 7225
rect 18138 7216 18144 7228
rect 18196 7256 18202 7268
rect 19076 7256 19104 7296
rect 19245 7293 19257 7296
rect 19291 7293 19303 7327
rect 19245 7287 19303 7293
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 19536 7333 19564 7364
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 19521 7327 19579 7333
rect 19521 7324 19533 7327
rect 19484 7296 19533 7324
rect 19484 7284 19490 7296
rect 19521 7293 19533 7296
rect 19567 7293 19579 7327
rect 19521 7287 19579 7293
rect 19797 7327 19855 7333
rect 19797 7293 19809 7327
rect 19843 7293 19855 7327
rect 19797 7287 19855 7293
rect 18196 7228 19104 7256
rect 19337 7259 19395 7265
rect 18196 7216 18202 7228
rect 19337 7225 19349 7259
rect 19383 7256 19395 7259
rect 19812 7256 19840 7287
rect 19383 7228 19840 7256
rect 19383 7225 19395 7228
rect 19337 7219 19395 7225
rect 17276 7160 17448 7188
rect 17276 7148 17282 7160
rect 17494 7148 17500 7200
rect 17552 7148 17558 7200
rect 18874 7148 18880 7200
rect 18932 7148 18938 7200
rect 552 7098 31531 7120
rect 552 7046 8102 7098
rect 8154 7046 8166 7098
rect 8218 7046 8230 7098
rect 8282 7046 8294 7098
rect 8346 7046 8358 7098
rect 8410 7046 15807 7098
rect 15859 7046 15871 7098
rect 15923 7046 15935 7098
rect 15987 7046 15999 7098
rect 16051 7046 16063 7098
rect 16115 7046 23512 7098
rect 23564 7046 23576 7098
rect 23628 7046 23640 7098
rect 23692 7046 23704 7098
rect 23756 7046 23768 7098
rect 23820 7046 31217 7098
rect 31269 7046 31281 7098
rect 31333 7046 31345 7098
rect 31397 7046 31409 7098
rect 31461 7046 31473 7098
rect 31525 7046 31531 7098
rect 552 7024 31531 7046
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 11238 6984 11244 6996
rect 9916 6956 11244 6984
rect 9916 6944 9922 6956
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 11422 6944 11428 6996
rect 11480 6944 11486 6996
rect 11698 6944 11704 6996
rect 11756 6944 11762 6996
rect 11882 6944 11888 6996
rect 11940 6984 11946 6996
rect 11940 6956 12664 6984
rect 11940 6944 11946 6956
rect 8570 6808 8576 6860
rect 8628 6808 8634 6860
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9732 6820 10057 6848
rect 9732 6808 9738 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10134 6808 10140 6860
rect 10192 6808 10198 6860
rect 10313 6851 10371 6857
rect 10313 6817 10325 6851
rect 10359 6848 10371 6851
rect 10410 6848 10416 6860
rect 10359 6820 10416 6848
rect 10359 6817 10371 6820
rect 10313 6811 10371 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10594 6808 10600 6860
rect 10652 6808 10658 6860
rect 10778 6808 10784 6860
rect 10836 6838 10842 6860
rect 11440 6857 11468 6944
rect 10965 6851 11023 6857
rect 10965 6838 10977 6851
rect 10836 6817 10977 6838
rect 11011 6817 11023 6851
rect 10836 6811 11023 6817
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 11716 6848 11744 6944
rect 11808 6888 12480 6916
rect 11808 6857 11836 6888
rect 11563 6820 11744 6848
rect 11793 6851 11851 6857
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 11793 6817 11805 6851
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 10836 6810 11008 6811
rect 10836 6808 10842 6810
rect 8588 6780 8616 6808
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 8588 6752 11621 6780
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 11808 6780 11836 6811
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12069 6851 12127 6857
rect 12452 6855 12480 6888
rect 12526 6876 12532 6928
rect 12584 6876 12590 6928
rect 12636 6916 12664 6956
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 13357 6987 13415 6993
rect 13357 6984 13369 6987
rect 12952 6956 13369 6984
rect 12952 6944 12958 6956
rect 13357 6953 13369 6956
rect 13403 6953 13415 6987
rect 13357 6947 13415 6953
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13504 6956 13645 6984
rect 13504 6944 13510 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 13909 6987 13967 6993
rect 13909 6953 13921 6987
rect 13955 6984 13967 6987
rect 13998 6984 14004 6996
rect 13955 6956 14004 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14366 6984 14372 6996
rect 14148 6956 14372 6984
rect 14148 6944 14154 6956
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 14458 6944 14464 6996
rect 14516 6944 14522 6996
rect 15102 6944 15108 6996
rect 15160 6944 15166 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15841 6987 15899 6993
rect 15841 6984 15853 6987
rect 15252 6956 15853 6984
rect 15252 6944 15258 6956
rect 15841 6953 15853 6956
rect 15887 6953 15899 6987
rect 15841 6947 15899 6953
rect 16209 6987 16267 6993
rect 16209 6953 16221 6987
rect 16255 6984 16267 6987
rect 16298 6984 16304 6996
rect 16255 6956 16304 6984
rect 16255 6953 16267 6956
rect 16209 6947 16267 6953
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 16574 6944 16580 6996
rect 16632 6944 16638 6996
rect 16666 6944 16672 6996
rect 16724 6984 16730 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 16724 6956 17969 6984
rect 16724 6944 16730 6956
rect 13538 6916 13544 6928
rect 12636 6888 13544 6916
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 14737 6919 14795 6925
rect 13648 6888 14228 6916
rect 12069 6848 12081 6851
rect 12032 6820 12081 6848
rect 12032 6808 12038 6820
rect 12069 6817 12081 6820
rect 12115 6817 12127 6851
rect 12069 6811 12127 6817
rect 12437 6849 12495 6855
rect 12437 6815 12449 6849
rect 12483 6815 12495 6849
rect 12544 6848 12572 6876
rect 13648 6860 13676 6888
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12544 6820 12725 6848
rect 12437 6809 12495 6815
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 11609 6743 11667 6749
rect 11716 6752 11836 6780
rect 11885 6783 11943 6789
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 9858 6712 9864 6724
rect 8720 6684 9864 6712
rect 8720 6672 8726 6684
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 11333 6715 11391 6721
rect 11333 6712 11345 6715
rect 10928 6684 11345 6712
rect 10928 6672 10934 6684
rect 11333 6681 11345 6684
rect 11379 6681 11391 6715
rect 11333 6675 11391 6681
rect 11514 6672 11520 6724
rect 11572 6672 11578 6724
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 10689 6647 10747 6653
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 10962 6644 10968 6656
rect 10735 6616 10968 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11057 6647 11115 6653
rect 11057 6613 11069 6647
rect 11103 6644 11115 6647
rect 11532 6644 11560 6672
rect 11716 6656 11744 6752
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12529 6783 12587 6789
rect 11931 6752 12434 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 11103 6616 11560 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11698 6604 11704 6656
rect 11756 6604 11762 6656
rect 12406 6644 12434 6752
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 13004 6780 13032 6811
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 13228 6820 13277 6848
rect 13228 6808 13234 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13630 6808 13636 6860
rect 13688 6808 13694 6860
rect 13725 6851 13783 6857
rect 13725 6817 13737 6851
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 12575 6752 13032 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 13740 6712 13768 6811
rect 13998 6808 14004 6860
rect 14056 6808 14062 6860
rect 14093 6851 14151 6857
rect 14093 6817 14105 6851
rect 14139 6817 14151 6851
rect 14200 6848 14228 6888
rect 14737 6885 14749 6919
rect 14783 6916 14795 6919
rect 14918 6916 14924 6928
rect 14783 6888 14924 6916
rect 14783 6885 14795 6888
rect 14737 6879 14795 6885
rect 14918 6876 14924 6888
rect 14976 6876 14982 6928
rect 15120 6916 15148 6944
rect 15120 6888 15240 6916
rect 15212 6857 15240 6888
rect 15378 6876 15384 6928
rect 15436 6876 15442 6928
rect 15562 6876 15568 6928
rect 15620 6916 15626 6928
rect 15620 6888 16528 6916
rect 15620 6876 15626 6888
rect 15105 6851 15163 6857
rect 15105 6848 15117 6851
rect 14200 6820 15117 6848
rect 14093 6811 14151 6817
rect 15105 6817 15117 6820
rect 15151 6817 15163 6851
rect 15105 6811 15163 6817
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6817 15255 6851
rect 15396 6848 15424 6876
rect 16500 6857 16528 6888
rect 16592 6857 16620 6944
rect 15473 6851 15531 6857
rect 15473 6848 15485 6851
rect 15396 6820 15485 6848
rect 15197 6811 15255 6817
rect 15473 6817 15485 6820
rect 15519 6817 15531 6851
rect 15473 6811 15531 6817
rect 15933 6851 15991 6857
rect 15933 6817 15945 6851
rect 15979 6817 15991 6851
rect 15933 6811 15991 6817
rect 16117 6851 16175 6857
rect 16117 6817 16129 6851
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6817 16635 6851
rect 16577 6811 16635 6817
rect 14108 6780 14136 6811
rect 14274 6780 14280 6792
rect 14108 6752 14280 6780
rect 14274 6740 14280 6752
rect 14332 6780 14338 6792
rect 15948 6780 15976 6811
rect 14332 6752 15976 6780
rect 16132 6780 16160 6811
rect 16684 6780 16712 6944
rect 16942 6876 16948 6928
rect 17000 6876 17006 6928
rect 17494 6916 17500 6928
rect 17052 6888 17500 6916
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 16960 6848 16988 6876
rect 17052 6857 17080 6888
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 16807 6820 16988 6848
rect 17037 6851 17095 6857
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 17037 6817 17049 6851
rect 17083 6817 17095 6851
rect 17037 6811 17095 6817
rect 17218 6808 17224 6860
rect 17276 6808 17282 6860
rect 17310 6808 17316 6860
rect 17368 6808 17374 6860
rect 17402 6808 17408 6860
rect 17460 6808 17466 6860
rect 17604 6857 17632 6956
rect 17957 6953 17969 6956
rect 18003 6984 18015 6987
rect 19426 6984 19432 6996
rect 18003 6956 19432 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 19518 6944 19524 6996
rect 19576 6944 19582 6996
rect 18138 6876 18144 6928
rect 18196 6876 18202 6928
rect 19536 6916 19564 6944
rect 18524 6888 19564 6916
rect 20180 6888 20392 6916
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6817 17647 6851
rect 17589 6811 17647 6817
rect 18046 6808 18052 6860
rect 18104 6808 18110 6860
rect 18156 6847 18184 6876
rect 18233 6851 18291 6857
rect 18141 6841 18199 6847
rect 18141 6807 18153 6841
rect 18187 6807 18199 6841
rect 18233 6817 18245 6851
rect 18279 6848 18291 6851
rect 18524 6848 18552 6888
rect 18279 6820 18552 6848
rect 18601 6851 18659 6857
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 18601 6817 18613 6851
rect 18647 6848 18659 6851
rect 20180 6848 20208 6888
rect 18647 6820 20208 6848
rect 18647 6817 18659 6820
rect 18601 6811 18659 6817
rect 20254 6808 20260 6860
rect 20312 6808 20318 6860
rect 20364 6848 20392 6888
rect 21358 6848 21364 6860
rect 20364 6820 21364 6848
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 18141 6801 18199 6807
rect 20272 6780 20300 6808
rect 16132 6752 16712 6780
rect 18248 6752 20300 6780
rect 14332 6740 14338 6752
rect 14550 6712 14556 6724
rect 13740 6684 14556 6712
rect 14550 6672 14556 6684
rect 14608 6672 14614 6724
rect 15470 6672 15476 6724
rect 15528 6712 15534 6724
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 15528 6684 15577 6712
rect 15528 6672 15534 6684
rect 15565 6681 15577 6684
rect 15611 6681 15623 6715
rect 15565 6675 15623 6681
rect 12526 6644 12532 6656
rect 12406 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12805 6647 12863 6653
rect 12805 6613 12817 6647
rect 12851 6644 12863 6647
rect 13081 6647 13139 6653
rect 13081 6644 13093 6647
rect 12851 6616 13093 6644
rect 12851 6613 12863 6616
rect 12805 6607 12863 6613
rect 13081 6613 13093 6616
rect 13127 6613 13139 6647
rect 13081 6607 13139 6613
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 15102 6644 15108 6656
rect 14231 6616 15108 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 17129 6647 17187 6653
rect 17129 6644 17141 6647
rect 16899 6616 17141 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 17129 6613 17141 6616
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 17681 6647 17739 6653
rect 17681 6613 17693 6647
rect 17727 6644 17739 6647
rect 18248 6644 18276 6752
rect 20438 6740 20444 6792
rect 20496 6740 20502 6792
rect 20530 6740 20536 6792
rect 20588 6740 20594 6792
rect 18509 6715 18567 6721
rect 18509 6681 18521 6715
rect 18555 6712 18567 6715
rect 20456 6712 20484 6740
rect 18555 6684 20484 6712
rect 18555 6681 18567 6684
rect 18509 6675 18567 6681
rect 17727 6616 18276 6644
rect 17727 6613 17739 6616
rect 17681 6607 17739 6613
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 20548 6644 20576 6740
rect 18380 6616 20576 6644
rect 18380 6604 18386 6616
rect 552 6554 31372 6576
rect 552 6502 4250 6554
rect 4302 6502 4314 6554
rect 4366 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 11955 6554
rect 12007 6502 12019 6554
rect 12071 6502 12083 6554
rect 12135 6502 12147 6554
rect 12199 6502 12211 6554
rect 12263 6502 19660 6554
rect 19712 6502 19724 6554
rect 19776 6502 19788 6554
rect 19840 6502 19852 6554
rect 19904 6502 19916 6554
rect 19968 6502 27365 6554
rect 27417 6502 27429 6554
rect 27481 6502 27493 6554
rect 27545 6502 27557 6554
rect 27609 6502 27621 6554
rect 27673 6502 31372 6554
rect 552 6480 31372 6502
rect 10134 6400 10140 6452
rect 10192 6400 10198 6452
rect 10410 6400 10416 6452
rect 10468 6400 10474 6452
rect 10502 6400 10508 6452
rect 10560 6400 10566 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10612 6412 10977 6440
rect 10152 6168 10180 6400
rect 10428 6236 10456 6400
rect 10520 6304 10548 6400
rect 10612 6384 10640 6412
rect 10965 6409 10977 6412
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11204 6412 11529 6440
rect 11204 6400 11210 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11756 6412 11805 6440
rect 11756 6400 11762 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 12768 6412 13185 6440
rect 12768 6400 12774 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13909 6443 13967 6449
rect 13909 6440 13921 6443
rect 13412 6412 13921 6440
rect 13412 6400 13418 6412
rect 13909 6409 13921 6412
rect 13955 6409 13967 6443
rect 13909 6403 13967 6409
rect 14366 6400 14372 6452
rect 14424 6400 14430 6452
rect 14550 6400 14556 6452
rect 14608 6400 14614 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 16117 6443 16175 6449
rect 16117 6440 16129 6443
rect 15712 6412 16129 6440
rect 15712 6400 15718 6412
rect 16117 6409 16129 6412
rect 16163 6409 16175 6443
rect 16117 6403 16175 6409
rect 10594 6332 10600 6384
rect 10652 6332 10658 6384
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 12342 6372 12348 6384
rect 11480 6344 12348 6372
rect 11480 6332 11486 6344
rect 12342 6332 12348 6344
rect 12400 6372 12406 6384
rect 12400 6344 12572 6372
rect 12400 6332 12406 6344
rect 10520 6276 11192 6304
rect 11164 6245 11192 6276
rect 11238 6264 11244 6316
rect 11296 6264 11302 6316
rect 11514 6264 11520 6316
rect 11572 6304 11578 6316
rect 11572 6276 11652 6304
rect 11572 6264 11578 6276
rect 11624 6245 11652 6276
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 11756 6276 11928 6304
rect 11756 6264 11762 6276
rect 11900 6245 11928 6276
rect 12544 6245 12572 6344
rect 13446 6332 13452 6384
rect 13504 6332 13510 6384
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 13633 6375 13691 6381
rect 13633 6372 13645 6375
rect 13596 6344 13645 6372
rect 13596 6332 13602 6344
rect 13633 6341 13645 6344
rect 13679 6341 13691 6375
rect 13633 6335 13691 6341
rect 13464 6304 13492 6332
rect 14384 6304 14412 6400
rect 13464 6276 14044 6304
rect 14384 6276 15792 6304
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10428 6208 10885 6236
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 11149 6239 11207 6245
rect 11149 6205 11161 6239
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 11609 6239 11667 6245
rect 11609 6205 11621 6239
rect 11655 6205 11667 6239
rect 11609 6199 11667 6205
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 11977 6239 12035 6245
rect 11977 6236 11989 6239
rect 11931 6208 11989 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 11977 6205 11989 6208
rect 12023 6205 12035 6239
rect 11977 6199 12035 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 12529 6199 12587 6205
rect 11072 6168 11100 6199
rect 12268 6168 12296 6199
rect 12802 6196 12808 6248
rect 12860 6196 12866 6248
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6236 13323 6239
rect 13464 6236 13492 6276
rect 13311 6208 13492 6236
rect 13541 6239 13599 6245
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 13541 6205 13553 6239
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 10152 6140 11100 6168
rect 11992 6140 12296 6168
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 11992 6100 12020 6140
rect 12986 6128 12992 6180
rect 13044 6168 13050 6180
rect 13556 6168 13584 6199
rect 13722 6196 13728 6248
rect 13780 6196 13786 6248
rect 14016 6245 14044 6276
rect 14001 6239 14059 6245
rect 14001 6205 14013 6239
rect 14047 6236 14059 6239
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 14047 6208 14105 6236
rect 14047 6205 14059 6208
rect 14001 6199 14059 6205
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 14844 6245 14872 6276
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14240 6208 14657 6236
rect 14240 6196 14246 6208
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 15102 6196 15108 6248
rect 15160 6196 15166 6248
rect 15764 6245 15792 6276
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15887 6208 16037 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 13044 6140 13584 6168
rect 13740 6168 13768 6196
rect 15304 6168 15332 6199
rect 13740 6140 15332 6168
rect 13044 6128 13050 6140
rect 10744 6072 12020 6100
rect 10744 6060 10750 6072
rect 12066 6060 12072 6112
rect 12124 6060 12130 6112
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 12345 6103 12403 6109
rect 12345 6100 12357 6103
rect 12216 6072 12357 6100
rect 12216 6060 12222 6072
rect 12345 6069 12357 6072
rect 12391 6069 12403 6103
rect 12345 6063 12403 6069
rect 12618 6060 12624 6112
rect 12676 6060 12682 6112
rect 12894 6060 12900 6112
rect 12952 6060 12958 6112
rect 14182 6060 14188 6112
rect 14240 6060 14246 6112
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 14967 6072 15117 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 552 6010 31531 6032
rect 552 5958 8102 6010
rect 8154 5958 8166 6010
rect 8218 5958 8230 6010
rect 8282 5958 8294 6010
rect 8346 5958 8358 6010
rect 8410 5958 15807 6010
rect 15859 5958 15871 6010
rect 15923 5958 15935 6010
rect 15987 5958 15999 6010
rect 16051 5958 16063 6010
rect 16115 5958 23512 6010
rect 23564 5958 23576 6010
rect 23628 5958 23640 6010
rect 23692 5958 23704 6010
rect 23756 5958 23768 6010
rect 23820 5958 31217 6010
rect 31269 5958 31281 6010
rect 31333 5958 31345 6010
rect 31397 5958 31409 6010
rect 31461 5958 31473 6010
rect 31525 5958 31531 6010
rect 552 5936 31531 5958
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 10778 5896 10784 5908
rect 8812 5868 10784 5896
rect 8812 5856 8818 5868
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 11112 5868 12265 5896
rect 11112 5856 11118 5868
rect 12253 5865 12265 5868
rect 12299 5865 12311 5899
rect 12253 5859 12311 5865
rect 12342 5856 12348 5908
rect 12400 5856 12406 5908
rect 12618 5856 12624 5908
rect 12676 5856 12682 5908
rect 12713 5899 12771 5905
rect 12713 5865 12725 5899
rect 12759 5896 12771 5899
rect 12894 5896 12900 5908
rect 12759 5868 12900 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 13909 5899 13967 5905
rect 13909 5896 13921 5899
rect 13872 5868 13921 5896
rect 13872 5856 13878 5868
rect 13909 5865 13921 5868
rect 13955 5865 13967 5899
rect 13909 5859 13967 5865
rect 14182 5856 14188 5908
rect 14240 5856 14246 5908
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 9824 5800 11284 5828
rect 9824 5788 9830 5800
rect 11256 5769 11284 5800
rect 11330 5788 11336 5840
rect 11388 5788 11394 5840
rect 12360 5769 12388 5856
rect 12636 5828 12664 5856
rect 12636 5800 12940 5828
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 12345 5763 12403 5769
rect 11241 5723 11299 5729
rect 11440 5732 12296 5760
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 11440 5692 11468 5732
rect 9456 5664 11468 5692
rect 12268 5692 12296 5732
rect 12345 5729 12357 5763
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 12912 5769 12940 5800
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12584 5732 12633 5760
rect 12584 5720 12590 5732
rect 12621 5729 12633 5732
rect 12667 5729 12679 5763
rect 12621 5723 12679 5729
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 13078 5720 13084 5772
rect 13136 5720 13142 5772
rect 14001 5763 14059 5769
rect 14001 5729 14013 5763
rect 14047 5760 14059 5763
rect 14200 5760 14228 5856
rect 14047 5732 14228 5760
rect 14047 5729 14059 5732
rect 14001 5723 14059 5729
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12268 5664 13001 5692
rect 9456 5652 9462 5664
rect 12989 5661 13001 5664
rect 13035 5661 13047 5695
rect 12989 5655 13047 5661
rect 8938 5584 8944 5636
rect 8996 5624 9002 5636
rect 12066 5624 12072 5636
rect 8996 5596 12072 5624
rect 8996 5584 9002 5596
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 12158 5556 12164 5568
rect 8076 5528 12164 5556
rect 8076 5516 8082 5528
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 552 5466 31372 5488
rect 552 5414 4250 5466
rect 4302 5414 4314 5466
rect 4366 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 11955 5466
rect 12007 5414 12019 5466
rect 12071 5414 12083 5466
rect 12135 5414 12147 5466
rect 12199 5414 12211 5466
rect 12263 5414 19660 5466
rect 19712 5414 19724 5466
rect 19776 5414 19788 5466
rect 19840 5414 19852 5466
rect 19904 5414 19916 5466
rect 19968 5414 27365 5466
rect 27417 5414 27429 5466
rect 27481 5414 27493 5466
rect 27545 5414 27557 5466
rect 27609 5414 27621 5466
rect 27673 5414 31372 5466
rect 552 5392 31372 5414
rect 552 4922 31531 4944
rect 552 4870 8102 4922
rect 8154 4870 8166 4922
rect 8218 4870 8230 4922
rect 8282 4870 8294 4922
rect 8346 4870 8358 4922
rect 8410 4870 15807 4922
rect 15859 4870 15871 4922
rect 15923 4870 15935 4922
rect 15987 4870 15999 4922
rect 16051 4870 16063 4922
rect 16115 4870 23512 4922
rect 23564 4870 23576 4922
rect 23628 4870 23640 4922
rect 23692 4870 23704 4922
rect 23756 4870 23768 4922
rect 23820 4870 31217 4922
rect 31269 4870 31281 4922
rect 31333 4870 31345 4922
rect 31397 4870 31409 4922
rect 31461 4870 31473 4922
rect 31525 4870 31531 4922
rect 552 4848 31531 4870
rect 552 4378 31372 4400
rect 552 4326 4250 4378
rect 4302 4326 4314 4378
rect 4366 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 11955 4378
rect 12007 4326 12019 4378
rect 12071 4326 12083 4378
rect 12135 4326 12147 4378
rect 12199 4326 12211 4378
rect 12263 4326 19660 4378
rect 19712 4326 19724 4378
rect 19776 4326 19788 4378
rect 19840 4326 19852 4378
rect 19904 4326 19916 4378
rect 19968 4326 27365 4378
rect 27417 4326 27429 4378
rect 27481 4326 27493 4378
rect 27545 4326 27557 4378
rect 27609 4326 27621 4378
rect 27673 4326 31372 4378
rect 552 4304 31372 4326
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 15286 4128 15292 4140
rect 14240 4100 15292 4128
rect 14240 4088 14246 4100
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 552 3834 31531 3856
rect 552 3782 8102 3834
rect 8154 3782 8166 3834
rect 8218 3782 8230 3834
rect 8282 3782 8294 3834
rect 8346 3782 8358 3834
rect 8410 3782 15807 3834
rect 15859 3782 15871 3834
rect 15923 3782 15935 3834
rect 15987 3782 15999 3834
rect 16051 3782 16063 3834
rect 16115 3782 23512 3834
rect 23564 3782 23576 3834
rect 23628 3782 23640 3834
rect 23692 3782 23704 3834
rect 23756 3782 23768 3834
rect 23820 3782 31217 3834
rect 31269 3782 31281 3834
rect 31333 3782 31345 3834
rect 31397 3782 31409 3834
rect 31461 3782 31473 3834
rect 31525 3782 31531 3834
rect 552 3760 31531 3782
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 13906 3516 13912 3528
rect 9732 3488 13912 3516
rect 9732 3476 9738 3488
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 552 3290 31372 3312
rect 552 3238 4250 3290
rect 4302 3238 4314 3290
rect 4366 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 11955 3290
rect 12007 3238 12019 3290
rect 12071 3238 12083 3290
rect 12135 3238 12147 3290
rect 12199 3238 12211 3290
rect 12263 3238 19660 3290
rect 19712 3238 19724 3290
rect 19776 3238 19788 3290
rect 19840 3238 19852 3290
rect 19904 3238 19916 3290
rect 19968 3238 27365 3290
rect 27417 3238 27429 3290
rect 27481 3238 27493 3290
rect 27545 3238 27557 3290
rect 27609 3238 27621 3290
rect 27673 3238 31372 3290
rect 552 3216 31372 3238
rect 552 2746 31531 2768
rect 552 2694 8102 2746
rect 8154 2694 8166 2746
rect 8218 2694 8230 2746
rect 8282 2694 8294 2746
rect 8346 2694 8358 2746
rect 8410 2694 15807 2746
rect 15859 2694 15871 2746
rect 15923 2694 15935 2746
rect 15987 2694 15999 2746
rect 16051 2694 16063 2746
rect 16115 2694 23512 2746
rect 23564 2694 23576 2746
rect 23628 2694 23640 2746
rect 23692 2694 23704 2746
rect 23756 2694 23768 2746
rect 23820 2694 31217 2746
rect 31269 2694 31281 2746
rect 31333 2694 31345 2746
rect 31397 2694 31409 2746
rect 31461 2694 31473 2746
rect 31525 2694 31531 2746
rect 552 2672 31531 2694
rect 552 2202 31372 2224
rect 552 2150 4250 2202
rect 4302 2150 4314 2202
rect 4366 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 11955 2202
rect 12007 2150 12019 2202
rect 12071 2150 12083 2202
rect 12135 2150 12147 2202
rect 12199 2150 12211 2202
rect 12263 2150 19660 2202
rect 19712 2150 19724 2202
rect 19776 2150 19788 2202
rect 19840 2150 19852 2202
rect 19904 2150 19916 2202
rect 19968 2150 27365 2202
rect 27417 2150 27429 2202
rect 27481 2150 27493 2202
rect 27545 2150 27557 2202
rect 27609 2150 27621 2202
rect 27673 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31531 1680
rect 552 1606 8102 1658
rect 8154 1606 8166 1658
rect 8218 1606 8230 1658
rect 8282 1606 8294 1658
rect 8346 1606 8358 1658
rect 8410 1606 15807 1658
rect 15859 1606 15871 1658
rect 15923 1606 15935 1658
rect 15987 1606 15999 1658
rect 16051 1606 16063 1658
rect 16115 1606 23512 1658
rect 23564 1606 23576 1658
rect 23628 1606 23640 1658
rect 23692 1606 23704 1658
rect 23756 1606 23768 1658
rect 23820 1606 31217 1658
rect 31269 1606 31281 1658
rect 31333 1606 31345 1658
rect 31397 1606 31409 1658
rect 31461 1606 31473 1658
rect 31525 1606 31531 1658
rect 552 1584 31531 1606
rect 552 1114 31372 1136
rect 552 1062 4250 1114
rect 4302 1062 4314 1114
rect 4366 1062 4378 1114
rect 4430 1062 4442 1114
rect 4494 1062 4506 1114
rect 4558 1062 11955 1114
rect 12007 1062 12019 1114
rect 12071 1062 12083 1114
rect 12135 1062 12147 1114
rect 12199 1062 12211 1114
rect 12263 1062 19660 1114
rect 19712 1062 19724 1114
rect 19776 1062 19788 1114
rect 19840 1062 19852 1114
rect 19904 1062 19916 1114
rect 19968 1062 27365 1114
rect 27417 1062 27429 1114
rect 27481 1062 27493 1114
rect 27545 1062 27557 1114
rect 27609 1062 27621 1114
rect 27673 1062 31372 1114
rect 552 1040 31372 1062
rect 552 570 31531 592
rect 552 518 8102 570
rect 8154 518 8166 570
rect 8218 518 8230 570
rect 8282 518 8294 570
rect 8346 518 8358 570
rect 8410 518 15807 570
rect 15859 518 15871 570
rect 15923 518 15935 570
rect 15987 518 15999 570
rect 16051 518 16063 570
rect 16115 518 23512 570
rect 23564 518 23576 570
rect 23628 518 23640 570
rect 23692 518 23704 570
rect 23756 518 23768 570
rect 23820 518 31217 570
rect 31269 518 31281 570
rect 31333 518 31345 570
rect 31397 518 31409 570
rect 31461 518 31473 570
rect 31525 518 31531 570
rect 552 496 31531 518
<< via1 >>
rect 8102 19014 8154 19066
rect 8166 19014 8218 19066
rect 8230 19014 8282 19066
rect 8294 19014 8346 19066
rect 8358 19014 8410 19066
rect 15807 19014 15859 19066
rect 15871 19014 15923 19066
rect 15935 19014 15987 19066
rect 15999 19014 16051 19066
rect 16063 19014 16115 19066
rect 23512 19014 23564 19066
rect 23576 19014 23628 19066
rect 23640 19014 23692 19066
rect 23704 19014 23756 19066
rect 23768 19014 23820 19066
rect 31217 19014 31269 19066
rect 31281 19014 31333 19066
rect 31345 19014 31397 19066
rect 31409 19014 31461 19066
rect 31473 19014 31525 19066
rect 13544 18912 13596 18964
rect 13636 18615 13688 18624
rect 13636 18581 13645 18615
rect 13645 18581 13679 18615
rect 13679 18581 13688 18615
rect 13636 18572 13688 18581
rect 4250 18470 4302 18522
rect 4314 18470 4366 18522
rect 4378 18470 4430 18522
rect 4442 18470 4494 18522
rect 4506 18470 4558 18522
rect 11955 18470 12007 18522
rect 12019 18470 12071 18522
rect 12083 18470 12135 18522
rect 12147 18470 12199 18522
rect 12211 18470 12263 18522
rect 19660 18470 19712 18522
rect 19724 18470 19776 18522
rect 19788 18470 19840 18522
rect 19852 18470 19904 18522
rect 19916 18470 19968 18522
rect 27365 18470 27417 18522
rect 27429 18470 27481 18522
rect 27493 18470 27545 18522
rect 27557 18470 27609 18522
rect 27621 18470 27673 18522
rect 8102 17926 8154 17978
rect 8166 17926 8218 17978
rect 8230 17926 8282 17978
rect 8294 17926 8346 17978
rect 8358 17926 8410 17978
rect 15807 17926 15859 17978
rect 15871 17926 15923 17978
rect 15935 17926 15987 17978
rect 15999 17926 16051 17978
rect 16063 17926 16115 17978
rect 23512 17926 23564 17978
rect 23576 17926 23628 17978
rect 23640 17926 23692 17978
rect 23704 17926 23756 17978
rect 23768 17926 23820 17978
rect 31217 17926 31269 17978
rect 31281 17926 31333 17978
rect 31345 17926 31397 17978
rect 31409 17926 31461 17978
rect 31473 17926 31525 17978
rect 4250 17382 4302 17434
rect 4314 17382 4366 17434
rect 4378 17382 4430 17434
rect 4442 17382 4494 17434
rect 4506 17382 4558 17434
rect 11955 17382 12007 17434
rect 12019 17382 12071 17434
rect 12083 17382 12135 17434
rect 12147 17382 12199 17434
rect 12211 17382 12263 17434
rect 19660 17382 19712 17434
rect 19724 17382 19776 17434
rect 19788 17382 19840 17434
rect 19852 17382 19904 17434
rect 19916 17382 19968 17434
rect 27365 17382 27417 17434
rect 27429 17382 27481 17434
rect 27493 17382 27545 17434
rect 27557 17382 27609 17434
rect 27621 17382 27673 17434
rect 8102 16838 8154 16890
rect 8166 16838 8218 16890
rect 8230 16838 8282 16890
rect 8294 16838 8346 16890
rect 8358 16838 8410 16890
rect 15807 16838 15859 16890
rect 15871 16838 15923 16890
rect 15935 16838 15987 16890
rect 15999 16838 16051 16890
rect 16063 16838 16115 16890
rect 23512 16838 23564 16890
rect 23576 16838 23628 16890
rect 23640 16838 23692 16890
rect 23704 16838 23756 16890
rect 23768 16838 23820 16890
rect 31217 16838 31269 16890
rect 31281 16838 31333 16890
rect 31345 16838 31397 16890
rect 31409 16838 31461 16890
rect 31473 16838 31525 16890
rect 4250 16294 4302 16346
rect 4314 16294 4366 16346
rect 4378 16294 4430 16346
rect 4442 16294 4494 16346
rect 4506 16294 4558 16346
rect 11955 16294 12007 16346
rect 12019 16294 12071 16346
rect 12083 16294 12135 16346
rect 12147 16294 12199 16346
rect 12211 16294 12263 16346
rect 19660 16294 19712 16346
rect 19724 16294 19776 16346
rect 19788 16294 19840 16346
rect 19852 16294 19904 16346
rect 19916 16294 19968 16346
rect 27365 16294 27417 16346
rect 27429 16294 27481 16346
rect 27493 16294 27545 16346
rect 27557 16294 27609 16346
rect 27621 16294 27673 16346
rect 8102 15750 8154 15802
rect 8166 15750 8218 15802
rect 8230 15750 8282 15802
rect 8294 15750 8346 15802
rect 8358 15750 8410 15802
rect 15807 15750 15859 15802
rect 15871 15750 15923 15802
rect 15935 15750 15987 15802
rect 15999 15750 16051 15802
rect 16063 15750 16115 15802
rect 23512 15750 23564 15802
rect 23576 15750 23628 15802
rect 23640 15750 23692 15802
rect 23704 15750 23756 15802
rect 23768 15750 23820 15802
rect 31217 15750 31269 15802
rect 31281 15750 31333 15802
rect 31345 15750 31397 15802
rect 31409 15750 31461 15802
rect 31473 15750 31525 15802
rect 4250 15206 4302 15258
rect 4314 15206 4366 15258
rect 4378 15206 4430 15258
rect 4442 15206 4494 15258
rect 4506 15206 4558 15258
rect 11955 15206 12007 15258
rect 12019 15206 12071 15258
rect 12083 15206 12135 15258
rect 12147 15206 12199 15258
rect 12211 15206 12263 15258
rect 19660 15206 19712 15258
rect 19724 15206 19776 15258
rect 19788 15206 19840 15258
rect 19852 15206 19904 15258
rect 19916 15206 19968 15258
rect 27365 15206 27417 15258
rect 27429 15206 27481 15258
rect 27493 15206 27545 15258
rect 27557 15206 27609 15258
rect 27621 15206 27673 15258
rect 8102 14662 8154 14714
rect 8166 14662 8218 14714
rect 8230 14662 8282 14714
rect 8294 14662 8346 14714
rect 8358 14662 8410 14714
rect 15807 14662 15859 14714
rect 15871 14662 15923 14714
rect 15935 14662 15987 14714
rect 15999 14662 16051 14714
rect 16063 14662 16115 14714
rect 23512 14662 23564 14714
rect 23576 14662 23628 14714
rect 23640 14662 23692 14714
rect 23704 14662 23756 14714
rect 23768 14662 23820 14714
rect 31217 14662 31269 14714
rect 31281 14662 31333 14714
rect 31345 14662 31397 14714
rect 31409 14662 31461 14714
rect 31473 14662 31525 14714
rect 4250 14118 4302 14170
rect 4314 14118 4366 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 11955 14118 12007 14170
rect 12019 14118 12071 14170
rect 12083 14118 12135 14170
rect 12147 14118 12199 14170
rect 12211 14118 12263 14170
rect 19660 14118 19712 14170
rect 19724 14118 19776 14170
rect 19788 14118 19840 14170
rect 19852 14118 19904 14170
rect 19916 14118 19968 14170
rect 27365 14118 27417 14170
rect 27429 14118 27481 14170
rect 27493 14118 27545 14170
rect 27557 14118 27609 14170
rect 27621 14118 27673 14170
rect 8102 13574 8154 13626
rect 8166 13574 8218 13626
rect 8230 13574 8282 13626
rect 8294 13574 8346 13626
rect 8358 13574 8410 13626
rect 15807 13574 15859 13626
rect 15871 13574 15923 13626
rect 15935 13574 15987 13626
rect 15999 13574 16051 13626
rect 16063 13574 16115 13626
rect 23512 13574 23564 13626
rect 23576 13574 23628 13626
rect 23640 13574 23692 13626
rect 23704 13574 23756 13626
rect 23768 13574 23820 13626
rect 31217 13574 31269 13626
rect 31281 13574 31333 13626
rect 31345 13574 31397 13626
rect 31409 13574 31461 13626
rect 31473 13574 31525 13626
rect 4250 13030 4302 13082
rect 4314 13030 4366 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 11955 13030 12007 13082
rect 12019 13030 12071 13082
rect 12083 13030 12135 13082
rect 12147 13030 12199 13082
rect 12211 13030 12263 13082
rect 19660 13030 19712 13082
rect 19724 13030 19776 13082
rect 19788 13030 19840 13082
rect 19852 13030 19904 13082
rect 19916 13030 19968 13082
rect 27365 13030 27417 13082
rect 27429 13030 27481 13082
rect 27493 13030 27545 13082
rect 27557 13030 27609 13082
rect 27621 13030 27673 13082
rect 8102 12486 8154 12538
rect 8166 12486 8218 12538
rect 8230 12486 8282 12538
rect 8294 12486 8346 12538
rect 8358 12486 8410 12538
rect 15807 12486 15859 12538
rect 15871 12486 15923 12538
rect 15935 12486 15987 12538
rect 15999 12486 16051 12538
rect 16063 12486 16115 12538
rect 23512 12486 23564 12538
rect 23576 12486 23628 12538
rect 23640 12486 23692 12538
rect 23704 12486 23756 12538
rect 23768 12486 23820 12538
rect 31217 12486 31269 12538
rect 31281 12486 31333 12538
rect 31345 12486 31397 12538
rect 31409 12486 31461 12538
rect 31473 12486 31525 12538
rect 11612 12384 11664 12436
rect 12256 12384 12308 12436
rect 11704 12248 11756 12300
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 12624 12248 12676 12300
rect 10968 12112 11020 12164
rect 14096 12291 14148 12300
rect 14096 12257 14105 12291
rect 14105 12257 14139 12291
rect 14139 12257 14148 12291
rect 14096 12248 14148 12257
rect 14648 12248 14700 12300
rect 16304 12291 16356 12300
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 19432 12359 19484 12368
rect 19432 12325 19441 12359
rect 19441 12325 19475 12359
rect 19475 12325 19484 12359
rect 19432 12316 19484 12325
rect 20076 12248 20128 12300
rect 11796 12044 11848 12096
rect 12348 12044 12400 12096
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 14004 12044 14056 12096
rect 15384 12044 15436 12096
rect 18788 12044 18840 12096
rect 4250 11942 4302 11994
rect 4314 11942 4366 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 11955 11942 12007 11994
rect 12019 11942 12071 11994
rect 12083 11942 12135 11994
rect 12147 11942 12199 11994
rect 12211 11942 12263 11994
rect 19660 11942 19712 11994
rect 19724 11942 19776 11994
rect 19788 11942 19840 11994
rect 19852 11942 19904 11994
rect 19916 11942 19968 11994
rect 27365 11942 27417 11994
rect 27429 11942 27481 11994
rect 27493 11942 27545 11994
rect 27557 11942 27609 11994
rect 27621 11942 27673 11994
rect 13912 11840 13964 11892
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 16304 11840 16356 11892
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 15016 11772 15068 11824
rect 8944 11704 8996 11756
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 11428 11636 11480 11688
rect 11796 11679 11848 11688
rect 11796 11645 11830 11679
rect 11830 11645 11848 11679
rect 11796 11636 11848 11645
rect 12164 11636 12216 11688
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 14096 11636 14148 11688
rect 15476 11679 15528 11688
rect 15476 11645 15485 11679
rect 15485 11645 15519 11679
rect 15519 11645 15528 11679
rect 15476 11636 15528 11645
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11152 11500 11204 11552
rect 11244 11500 11296 11552
rect 11796 11500 11848 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 15200 11611 15252 11620
rect 15200 11577 15209 11611
rect 15209 11577 15243 11611
rect 15243 11577 15252 11611
rect 15200 11568 15252 11577
rect 16304 11636 16356 11688
rect 16488 11679 16540 11688
rect 16488 11645 16497 11679
rect 16497 11645 16531 11679
rect 16531 11645 16540 11679
rect 16488 11636 16540 11645
rect 16856 11636 16908 11688
rect 18420 11636 18472 11688
rect 18788 11636 18840 11688
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 16212 11500 16264 11552
rect 8102 11398 8154 11450
rect 8166 11398 8218 11450
rect 8230 11398 8282 11450
rect 8294 11398 8346 11450
rect 8358 11398 8410 11450
rect 15807 11398 15859 11450
rect 15871 11398 15923 11450
rect 15935 11398 15987 11450
rect 15999 11398 16051 11450
rect 16063 11398 16115 11450
rect 23512 11398 23564 11450
rect 23576 11398 23628 11450
rect 23640 11398 23692 11450
rect 23704 11398 23756 11450
rect 23768 11398 23820 11450
rect 31217 11398 31269 11450
rect 31281 11398 31333 11450
rect 31345 11398 31397 11450
rect 31409 11398 31461 11450
rect 31473 11398 31525 11450
rect 11704 11296 11756 11348
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 12348 11296 12400 11348
rect 12900 11296 12952 11348
rect 12992 11339 13044 11348
rect 12992 11305 13001 11339
rect 13001 11305 13035 11339
rect 13035 11305 13044 11339
rect 12992 11296 13044 11305
rect 10876 11228 10928 11280
rect 10508 11203 10560 11212
rect 10508 11169 10517 11203
rect 10517 11169 10551 11203
rect 10551 11169 10560 11203
rect 10508 11160 10560 11169
rect 11244 11160 11296 11212
rect 12532 11203 12584 11212
rect 13544 11296 13596 11348
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 14096 11296 14148 11348
rect 15016 11296 15068 11348
rect 16488 11296 16540 11348
rect 13636 11228 13688 11280
rect 12532 11169 12561 11203
rect 12561 11169 12584 11203
rect 12532 11160 12584 11169
rect 14004 11203 14056 11212
rect 14004 11169 14013 11203
rect 14013 11169 14047 11203
rect 14047 11169 14056 11203
rect 14004 11160 14056 11169
rect 20076 11339 20128 11348
rect 20076 11305 20085 11339
rect 20085 11305 20119 11339
rect 20119 11305 20128 11339
rect 20076 11296 20128 11305
rect 9312 11024 9364 11076
rect 10600 11024 10652 11076
rect 13820 11092 13872 11144
rect 15108 11160 15160 11212
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 15568 11092 15620 11144
rect 16764 11092 16816 11144
rect 18420 11203 18472 11212
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 16304 11024 16356 11076
rect 10692 10999 10744 11008
rect 10692 10965 10701 10999
rect 10701 10965 10735 10999
rect 10735 10965 10744 10999
rect 10692 10956 10744 10965
rect 12348 10956 12400 11008
rect 13084 10956 13136 11008
rect 13912 10999 13964 11008
rect 13912 10965 13921 10999
rect 13921 10965 13955 10999
rect 13955 10965 13964 10999
rect 13912 10956 13964 10965
rect 14188 10999 14240 11008
rect 14188 10965 14197 10999
rect 14197 10965 14231 10999
rect 14231 10965 14240 10999
rect 14188 10956 14240 10965
rect 16212 10999 16264 11008
rect 16212 10965 16221 10999
rect 16221 10965 16255 10999
rect 16255 10965 16264 10999
rect 16212 10956 16264 10965
rect 16396 10956 16448 11008
rect 18604 10956 18656 11008
rect 4250 10854 4302 10906
rect 4314 10854 4366 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 11955 10854 12007 10906
rect 12019 10854 12071 10906
rect 12083 10854 12135 10906
rect 12147 10854 12199 10906
rect 12211 10854 12263 10906
rect 19660 10854 19712 10906
rect 19724 10854 19776 10906
rect 19788 10854 19840 10906
rect 19852 10854 19904 10906
rect 19916 10854 19968 10906
rect 27365 10854 27417 10906
rect 27429 10854 27481 10906
rect 27493 10854 27545 10906
rect 27557 10854 27609 10906
rect 27621 10854 27673 10906
rect 9036 10548 9088 10600
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 13820 10752 13872 10804
rect 13912 10752 13964 10804
rect 14188 10752 14240 10804
rect 15200 10752 15252 10804
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 16212 10752 16264 10804
rect 18880 10795 18932 10804
rect 18880 10761 18889 10795
rect 18889 10761 18923 10795
rect 18923 10761 18932 10795
rect 18880 10752 18932 10761
rect 11612 10684 11664 10736
rect 12440 10616 12492 10668
rect 9956 10548 10008 10557
rect 11428 10548 11480 10600
rect 13268 10616 13320 10668
rect 9404 10412 9456 10464
rect 11336 10412 11388 10464
rect 13176 10591 13228 10600
rect 13176 10557 13185 10591
rect 13185 10557 13219 10591
rect 13219 10557 13228 10591
rect 13176 10548 13228 10557
rect 14096 10684 14148 10736
rect 13728 10616 13780 10668
rect 13820 10591 13872 10600
rect 13820 10557 13829 10591
rect 13829 10557 13863 10591
rect 13863 10557 13872 10591
rect 13820 10548 13872 10557
rect 15384 10616 15436 10668
rect 15476 10616 15528 10668
rect 14004 10480 14056 10532
rect 15108 10548 15160 10600
rect 16764 10616 16816 10668
rect 16672 10548 16724 10600
rect 17868 10616 17920 10668
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 12348 10412 12400 10464
rect 12716 10455 12768 10464
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 12900 10412 12952 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 13360 10412 13412 10464
rect 14280 10455 14332 10464
rect 14280 10421 14289 10455
rect 14289 10421 14323 10455
rect 14323 10421 14332 10455
rect 14280 10412 14332 10421
rect 14372 10412 14424 10464
rect 16488 10455 16540 10464
rect 16488 10421 16497 10455
rect 16497 10421 16531 10455
rect 16531 10421 16540 10455
rect 16488 10412 16540 10421
rect 16580 10412 16632 10464
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 18236 10480 18288 10532
rect 18604 10548 18656 10600
rect 20536 10548 20588 10600
rect 19064 10480 19116 10532
rect 17316 10455 17368 10464
rect 17316 10421 17325 10455
rect 17325 10421 17359 10455
rect 17359 10421 17368 10455
rect 17316 10412 17368 10421
rect 17500 10412 17552 10464
rect 17592 10455 17644 10464
rect 17592 10421 17601 10455
rect 17601 10421 17635 10455
rect 17635 10421 17644 10455
rect 17592 10412 17644 10421
rect 18144 10455 18196 10464
rect 18144 10421 18153 10455
rect 18153 10421 18187 10455
rect 18187 10421 18196 10455
rect 18144 10412 18196 10421
rect 19524 10412 19576 10464
rect 19616 10455 19668 10464
rect 19616 10421 19625 10455
rect 19625 10421 19659 10455
rect 19659 10421 19668 10455
rect 19616 10412 19668 10421
rect 20168 10412 20220 10464
rect 8102 10310 8154 10362
rect 8166 10310 8218 10362
rect 8230 10310 8282 10362
rect 8294 10310 8346 10362
rect 8358 10310 8410 10362
rect 15807 10310 15859 10362
rect 15871 10310 15923 10362
rect 15935 10310 15987 10362
rect 15999 10310 16051 10362
rect 16063 10310 16115 10362
rect 23512 10310 23564 10362
rect 23576 10310 23628 10362
rect 23640 10310 23692 10362
rect 23704 10310 23756 10362
rect 23768 10310 23820 10362
rect 31217 10310 31269 10362
rect 31281 10310 31333 10362
rect 31345 10310 31397 10362
rect 31409 10310 31461 10362
rect 31473 10310 31525 10362
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 10508 10208 10560 10260
rect 10600 10208 10652 10260
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 10416 10140 10468 10192
rect 8208 9868 8260 9920
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10968 10208 11020 10260
rect 11152 10208 11204 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 11704 10208 11756 10260
rect 12624 10208 12676 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 12992 10208 13044 10260
rect 13084 10208 13136 10260
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 13268 10208 13320 10260
rect 13820 10208 13872 10260
rect 14280 10208 14332 10260
rect 9864 10004 9916 10056
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 10692 10004 10744 10056
rect 11612 10004 11664 10056
rect 12532 10072 12584 10124
rect 12900 10004 12952 10056
rect 15660 10072 15712 10124
rect 16580 10208 16632 10260
rect 19616 10208 19668 10260
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17316 10072 17368 10124
rect 20168 10208 20220 10260
rect 9496 9936 9548 9988
rect 10232 9936 10284 9988
rect 10508 9936 10560 9988
rect 10968 9936 11020 9988
rect 9680 9868 9732 9920
rect 10048 9868 10100 9920
rect 10600 9868 10652 9920
rect 11428 9868 11480 9920
rect 11612 9911 11664 9920
rect 11612 9877 11621 9911
rect 11621 9877 11655 9911
rect 11655 9877 11664 9911
rect 11612 9868 11664 9877
rect 12440 9868 12492 9920
rect 13544 9868 13596 9920
rect 17868 10004 17920 10056
rect 18420 10072 18472 10124
rect 31668 10140 31720 10192
rect 17776 9936 17828 9988
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 16396 9868 16448 9877
rect 17960 9911 18012 9920
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 19432 9868 19484 9920
rect 4250 9766 4302 9818
rect 4314 9766 4366 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 11955 9766 12007 9818
rect 12019 9766 12071 9818
rect 12083 9766 12135 9818
rect 12147 9766 12199 9818
rect 12211 9766 12263 9818
rect 19660 9766 19712 9818
rect 19724 9766 19776 9818
rect 19788 9766 19840 9818
rect 19852 9766 19904 9818
rect 19916 9766 19968 9818
rect 27365 9766 27417 9818
rect 27429 9766 27481 9818
rect 27493 9766 27545 9818
rect 27557 9766 27609 9818
rect 27621 9766 27673 9818
rect 9772 9664 9824 9716
rect 10692 9664 10744 9716
rect 11244 9664 11296 9716
rect 16396 9707 16448 9716
rect 16396 9673 16405 9707
rect 16405 9673 16439 9707
rect 16439 9673 16448 9707
rect 16396 9664 16448 9673
rect 17592 9664 17644 9716
rect 18420 9664 18472 9716
rect 19524 9664 19576 9716
rect 10140 9596 10192 9648
rect 16580 9596 16632 9648
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9220 9392 9272 9444
rect 9404 9503 9456 9512
rect 9404 9469 9438 9503
rect 9438 9469 9456 9503
rect 11520 9528 11572 9580
rect 9404 9460 9456 9469
rect 8852 9324 8904 9376
rect 11336 9460 11388 9512
rect 11612 9460 11664 9512
rect 15292 9528 15344 9580
rect 18512 9596 18564 9648
rect 19064 9596 19116 9648
rect 13728 9460 13780 9512
rect 14004 9460 14056 9512
rect 14372 9460 14424 9512
rect 17868 9528 17920 9580
rect 16488 9503 16540 9512
rect 16488 9469 16497 9503
rect 16497 9469 16531 9503
rect 16531 9469 16540 9503
rect 16488 9460 16540 9469
rect 17132 9460 17184 9512
rect 13268 9435 13320 9444
rect 13268 9401 13277 9435
rect 13277 9401 13311 9435
rect 13311 9401 13320 9435
rect 13268 9392 13320 9401
rect 17960 9392 18012 9444
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 12440 9324 12492 9376
rect 15384 9367 15436 9376
rect 15384 9333 15393 9367
rect 15393 9333 15427 9367
rect 15427 9333 15436 9367
rect 15384 9324 15436 9333
rect 17224 9324 17276 9376
rect 17500 9324 17552 9376
rect 17684 9324 17736 9376
rect 18972 9324 19024 9376
rect 8102 9222 8154 9274
rect 8166 9222 8218 9274
rect 8230 9222 8282 9274
rect 8294 9222 8346 9274
rect 8358 9222 8410 9274
rect 15807 9222 15859 9274
rect 15871 9222 15923 9274
rect 15935 9222 15987 9274
rect 15999 9222 16051 9274
rect 16063 9222 16115 9274
rect 23512 9222 23564 9274
rect 23576 9222 23628 9274
rect 23640 9222 23692 9274
rect 23704 9222 23756 9274
rect 23768 9222 23820 9274
rect 31217 9222 31269 9274
rect 31281 9222 31333 9274
rect 31345 9222 31397 9274
rect 31409 9222 31461 9274
rect 31473 9222 31525 9274
rect 9312 9120 9364 9172
rect 10784 9120 10836 9172
rect 10876 9120 10928 9172
rect 11520 9120 11572 9172
rect 11888 9120 11940 9172
rect 13268 9120 13320 9172
rect 15660 9120 15712 9172
rect 16304 9120 16356 9172
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 15384 9052 15436 9104
rect 19432 9052 19484 9104
rect 28264 9120 28316 9172
rect 8760 8984 8812 9036
rect 8852 9027 8904 9036
rect 8852 8993 8861 9027
rect 8861 8993 8895 9027
rect 8895 8993 8904 9027
rect 8852 8984 8904 8993
rect 8944 9027 8996 9036
rect 8944 8993 8953 9027
rect 8953 8993 8987 9027
rect 8987 8993 8996 9027
rect 8944 8984 8996 8993
rect 9128 8984 9180 9036
rect 9312 9027 9364 9036
rect 9312 8993 9346 9027
rect 9346 8993 9364 9027
rect 9312 8984 9364 8993
rect 9680 8984 9732 9036
rect 10508 8984 10560 9036
rect 10692 8984 10744 9036
rect 8300 8916 8352 8968
rect 11520 8984 11572 9036
rect 11704 8984 11756 9036
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 8760 8780 8812 8832
rect 11244 8848 11296 8900
rect 13912 9027 13964 9036
rect 13912 8993 13921 9027
rect 13921 8993 13955 9027
rect 13955 8993 13964 9027
rect 13912 8984 13964 8993
rect 15660 8984 15712 9036
rect 15752 8984 15804 9036
rect 12532 8916 12584 8968
rect 13636 8916 13688 8968
rect 16856 8984 16908 9036
rect 18328 8984 18380 9036
rect 19524 8984 19576 9036
rect 20352 9027 20404 9036
rect 20352 8993 20361 9027
rect 20361 8993 20395 9027
rect 20395 8993 20404 9027
rect 20352 8984 20404 8993
rect 20536 8984 20588 9036
rect 20904 8984 20956 9036
rect 16580 8916 16632 8968
rect 17868 8916 17920 8968
rect 20444 8916 20496 8968
rect 9680 8780 9732 8832
rect 9772 8780 9824 8832
rect 11060 8780 11112 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 11520 8780 11572 8832
rect 11704 8823 11756 8832
rect 11704 8789 11713 8823
rect 11713 8789 11747 8823
rect 11747 8789 11756 8823
rect 11704 8780 11756 8789
rect 13084 8848 13136 8900
rect 12624 8780 12676 8832
rect 14004 8848 14056 8900
rect 28264 8848 28316 8900
rect 13268 8780 13320 8832
rect 14648 8780 14700 8832
rect 17040 8780 17092 8832
rect 17960 8780 18012 8832
rect 19984 8780 20036 8832
rect 20536 8780 20588 8832
rect 21364 8823 21416 8832
rect 21364 8789 21373 8823
rect 21373 8789 21407 8823
rect 21407 8789 21416 8823
rect 21364 8780 21416 8789
rect 4250 8678 4302 8730
rect 4314 8678 4366 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 11955 8678 12007 8730
rect 12019 8678 12071 8730
rect 12083 8678 12135 8730
rect 12147 8678 12199 8730
rect 12211 8678 12263 8730
rect 19660 8678 19712 8730
rect 19724 8678 19776 8730
rect 19788 8678 19840 8730
rect 19852 8678 19904 8730
rect 19916 8678 19968 8730
rect 27365 8678 27417 8730
rect 27429 8678 27481 8730
rect 27493 8678 27545 8730
rect 27557 8678 27609 8730
rect 27621 8678 27673 8730
rect 8024 8576 8076 8628
rect 9312 8576 9364 8628
rect 9864 8576 9916 8628
rect 11152 8576 11204 8628
rect 11612 8576 11664 8628
rect 13084 8576 13136 8628
rect 13820 8576 13872 8628
rect 17132 8619 17184 8628
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17132 8576 17184 8585
rect 18972 8576 19024 8628
rect 20352 8576 20404 8628
rect 8852 8440 8904 8492
rect 8392 8372 8444 8424
rect 8024 8304 8076 8356
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 10784 8508 10836 8560
rect 11704 8508 11756 8560
rect 12808 8508 12860 8560
rect 13268 8551 13320 8560
rect 13268 8517 13277 8551
rect 13277 8517 13311 8551
rect 13311 8517 13320 8551
rect 13268 8508 13320 8517
rect 17684 8551 17736 8560
rect 17684 8517 17693 8551
rect 17693 8517 17727 8551
rect 17727 8517 17736 8551
rect 17684 8508 17736 8517
rect 18052 8508 18104 8560
rect 18144 8508 18196 8560
rect 9404 8440 9456 8492
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 8300 8236 8352 8288
rect 9036 8236 9088 8288
rect 9496 8372 9548 8424
rect 10140 8440 10192 8492
rect 10876 8440 10928 8492
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 10232 8372 10284 8424
rect 10324 8415 10376 8424
rect 10324 8381 10333 8415
rect 10333 8381 10367 8415
rect 10367 8381 10376 8415
rect 10324 8372 10376 8381
rect 10508 8372 10560 8424
rect 10600 8372 10652 8424
rect 11520 8440 11572 8492
rect 11612 8440 11664 8492
rect 9404 8347 9456 8356
rect 9404 8313 9413 8347
rect 9413 8313 9447 8347
rect 9447 8313 9456 8347
rect 9404 8304 9456 8313
rect 10968 8304 11020 8356
rect 9772 8236 9824 8288
rect 10416 8236 10468 8288
rect 10876 8236 10928 8288
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 11796 8236 11848 8288
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 12072 8236 12124 8288
rect 12624 8236 12676 8288
rect 12900 8236 12952 8288
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 15016 8440 15068 8492
rect 15292 8440 15344 8492
rect 16856 8440 16908 8492
rect 18328 8440 18380 8492
rect 19984 8440 20036 8492
rect 14280 8304 14332 8356
rect 14372 8236 14424 8288
rect 16212 8372 16264 8424
rect 16580 8372 16632 8424
rect 16948 8391 16957 8424
rect 16957 8391 16991 8424
rect 16991 8391 17000 8424
rect 16948 8372 17000 8391
rect 17132 8304 17184 8356
rect 17224 8304 17276 8356
rect 17776 8415 17828 8424
rect 17776 8381 17785 8415
rect 17785 8381 17819 8415
rect 17819 8381 17828 8415
rect 17776 8372 17828 8381
rect 17868 8415 17920 8424
rect 17868 8381 17877 8415
rect 17877 8381 17911 8415
rect 17911 8381 17920 8415
rect 17868 8372 17920 8381
rect 18236 8372 18288 8424
rect 17408 8304 17460 8356
rect 19432 8304 19484 8356
rect 20260 8347 20312 8356
rect 20260 8313 20269 8347
rect 20269 8313 20303 8347
rect 20303 8313 20312 8347
rect 20260 8304 20312 8313
rect 15200 8279 15252 8288
rect 15200 8245 15209 8279
rect 15209 8245 15243 8279
rect 15243 8245 15252 8279
rect 15200 8236 15252 8245
rect 15660 8236 15712 8288
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 16580 8279 16632 8288
rect 16580 8245 16589 8279
rect 16589 8245 16623 8279
rect 16623 8245 16632 8279
rect 16580 8236 16632 8245
rect 16672 8236 16724 8288
rect 19340 8236 19392 8288
rect 20812 8279 20864 8288
rect 20812 8245 20821 8279
rect 20821 8245 20855 8279
rect 20855 8245 20864 8279
rect 20812 8236 20864 8245
rect 8102 8134 8154 8186
rect 8166 8134 8218 8186
rect 8230 8134 8282 8186
rect 8294 8134 8346 8186
rect 8358 8134 8410 8186
rect 15807 8134 15859 8186
rect 15871 8134 15923 8186
rect 15935 8134 15987 8186
rect 15999 8134 16051 8186
rect 16063 8134 16115 8186
rect 23512 8134 23564 8186
rect 23576 8134 23628 8186
rect 23640 8134 23692 8186
rect 23704 8134 23756 8186
rect 23768 8134 23820 8186
rect 31217 8134 31269 8186
rect 31281 8134 31333 8186
rect 31345 8134 31397 8186
rect 31409 8134 31461 8186
rect 31473 8134 31525 8186
rect 8484 8032 8536 8084
rect 9036 8032 9088 8084
rect 8852 7964 8904 8016
rect 9588 7964 9640 8016
rect 9772 7964 9824 8016
rect 10692 7964 10744 8016
rect 10876 7964 10928 8016
rect 11152 8075 11204 8084
rect 11152 8041 11161 8075
rect 11161 8041 11195 8075
rect 11195 8041 11204 8075
rect 11152 8032 11204 8041
rect 11244 8032 11296 8084
rect 11428 8032 11480 8084
rect 11888 8032 11940 8084
rect 12072 8032 12124 8084
rect 9956 7896 10008 7948
rect 10508 7896 10560 7948
rect 10968 7896 11020 7948
rect 13452 8032 13504 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 14648 8075 14700 8084
rect 14648 8041 14657 8075
rect 14657 8041 14691 8075
rect 14691 8041 14700 8075
rect 14648 8032 14700 8041
rect 12900 7964 12952 8016
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 10324 7828 10376 7880
rect 11428 7828 11480 7880
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 12440 7828 12492 7880
rect 12072 7760 12124 7812
rect 12256 7760 12308 7812
rect 12532 7760 12584 7812
rect 9772 7692 9824 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 10876 7692 10928 7744
rect 10968 7692 11020 7744
rect 11612 7735 11664 7744
rect 11612 7701 11621 7735
rect 11621 7701 11655 7735
rect 11655 7701 11664 7735
rect 11612 7692 11664 7701
rect 12348 7692 12400 7744
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 13820 8007 13872 8016
rect 13820 7973 13829 8007
rect 13829 7973 13863 8007
rect 13863 7973 13872 8007
rect 13820 7964 13872 7973
rect 14004 7964 14056 8016
rect 14096 7896 14148 7948
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 14372 7896 14424 7948
rect 15568 8032 15620 8084
rect 15660 8032 15712 8084
rect 16304 8032 16356 8084
rect 16580 8032 16632 8084
rect 15108 7896 15160 7948
rect 15200 7828 15252 7880
rect 15476 7828 15528 7880
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 17224 8032 17276 8084
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 16672 7828 16724 7880
rect 17960 7828 18012 7880
rect 20352 7939 20404 7948
rect 20352 7905 20361 7939
rect 20361 7905 20395 7939
rect 20395 7905 20404 7939
rect 20352 7896 20404 7905
rect 14004 7760 14056 7812
rect 15384 7692 15436 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 16580 7760 16632 7812
rect 15476 7692 15528 7701
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 18236 7735 18288 7744
rect 18236 7701 18245 7735
rect 18245 7701 18279 7735
rect 18279 7701 18288 7735
rect 18236 7692 18288 7701
rect 20812 7760 20864 7812
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 4250 7590 4302 7642
rect 4314 7590 4366 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 11955 7590 12007 7642
rect 12019 7590 12071 7642
rect 12083 7590 12135 7642
rect 12147 7590 12199 7642
rect 12211 7590 12263 7642
rect 19660 7590 19712 7642
rect 19724 7590 19776 7642
rect 19788 7590 19840 7642
rect 19852 7590 19904 7642
rect 19916 7590 19968 7642
rect 27365 7590 27417 7642
rect 27429 7590 27481 7642
rect 27493 7590 27545 7642
rect 27557 7590 27609 7642
rect 27621 7590 27673 7642
rect 11152 7488 11204 7540
rect 11244 7488 11296 7540
rect 12716 7488 12768 7540
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 14188 7488 14240 7540
rect 15108 7488 15160 7540
rect 16672 7488 16724 7540
rect 18236 7488 18288 7540
rect 19340 7488 19392 7540
rect 19432 7488 19484 7540
rect 20352 7488 20404 7540
rect 9128 7420 9180 7472
rect 10968 7420 11020 7472
rect 12440 7420 12492 7472
rect 13360 7420 13412 7472
rect 9956 7352 10008 7404
rect 13544 7395 13596 7404
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 9956 7216 10008 7268
rect 10232 7148 10284 7200
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 11060 7284 11112 7336
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 15016 7352 15068 7404
rect 16948 7420 17000 7472
rect 10600 7216 10652 7268
rect 12624 7284 12676 7336
rect 12808 7284 12860 7336
rect 14096 7284 14148 7336
rect 11336 7216 11388 7268
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 13820 7259 13872 7268
rect 13820 7225 13854 7259
rect 13854 7225 13872 7259
rect 13820 7216 13872 7225
rect 17132 7284 17184 7336
rect 17316 7284 17368 7336
rect 19064 7420 19116 7472
rect 12624 7191 12676 7200
rect 12624 7157 12633 7191
rect 12633 7157 12667 7191
rect 12667 7157 12676 7191
rect 12624 7148 12676 7157
rect 13728 7148 13780 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 15384 7148 15436 7200
rect 15660 7259 15712 7268
rect 15660 7225 15694 7259
rect 15694 7225 15712 7259
rect 15660 7216 15712 7225
rect 16672 7216 16724 7268
rect 17040 7191 17092 7200
rect 17040 7157 17049 7191
rect 17049 7157 17083 7191
rect 17083 7157 17092 7191
rect 17040 7148 17092 7157
rect 17224 7148 17276 7200
rect 18144 7216 18196 7268
rect 19432 7284 19484 7336
rect 20628 7352 20680 7404
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 18880 7191 18932 7200
rect 18880 7157 18889 7191
rect 18889 7157 18923 7191
rect 18923 7157 18932 7191
rect 18880 7148 18932 7157
rect 8102 7046 8154 7098
rect 8166 7046 8218 7098
rect 8230 7046 8282 7098
rect 8294 7046 8346 7098
rect 8358 7046 8410 7098
rect 15807 7046 15859 7098
rect 15871 7046 15923 7098
rect 15935 7046 15987 7098
rect 15999 7046 16051 7098
rect 16063 7046 16115 7098
rect 23512 7046 23564 7098
rect 23576 7046 23628 7098
rect 23640 7046 23692 7098
rect 23704 7046 23756 7098
rect 23768 7046 23820 7098
rect 31217 7046 31269 7098
rect 31281 7046 31333 7098
rect 31345 7046 31397 7098
rect 31409 7046 31461 7098
rect 31473 7046 31525 7098
rect 9864 6944 9916 6996
rect 11244 6944 11296 6996
rect 11428 6944 11480 6996
rect 11704 6944 11756 6996
rect 11888 6944 11940 6996
rect 8576 6808 8628 6860
rect 9680 6808 9732 6860
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 10416 6808 10468 6860
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 10784 6808 10836 6860
rect 11980 6808 12032 6860
rect 12532 6876 12584 6928
rect 12900 6944 12952 6996
rect 13452 6944 13504 6996
rect 14004 6944 14056 6996
rect 14096 6944 14148 6996
rect 14372 6944 14424 6996
rect 14464 6987 14516 6996
rect 14464 6953 14473 6987
rect 14473 6953 14507 6987
rect 14507 6953 14516 6987
rect 14464 6944 14516 6953
rect 15108 6944 15160 6996
rect 15200 6944 15252 6996
rect 16304 6944 16356 6996
rect 16580 6944 16632 6996
rect 16672 6944 16724 6996
rect 13544 6876 13596 6928
rect 8668 6672 8720 6724
rect 9864 6672 9916 6724
rect 10876 6672 10928 6724
rect 11520 6672 11572 6724
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 10968 6604 11020 6656
rect 12164 6715 12216 6724
rect 12164 6681 12173 6715
rect 12173 6681 12207 6715
rect 12207 6681 12216 6715
rect 12164 6672 12216 6681
rect 11704 6604 11756 6656
rect 13176 6808 13228 6860
rect 13636 6808 13688 6860
rect 14004 6851 14056 6860
rect 14004 6817 14013 6851
rect 14013 6817 14047 6851
rect 14047 6817 14056 6851
rect 14004 6808 14056 6817
rect 14924 6876 14976 6928
rect 15384 6876 15436 6928
rect 15568 6876 15620 6928
rect 14280 6740 14332 6792
rect 16948 6876 17000 6928
rect 17500 6876 17552 6928
rect 17224 6851 17276 6860
rect 17224 6817 17233 6851
rect 17233 6817 17267 6851
rect 17267 6817 17276 6851
rect 17224 6808 17276 6817
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 19432 6944 19484 6996
rect 19524 6944 19576 6996
rect 18144 6876 18196 6928
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 20260 6808 20312 6860
rect 21364 6808 21416 6860
rect 14556 6672 14608 6724
rect 15476 6672 15528 6724
rect 12532 6604 12584 6656
rect 15108 6604 15160 6656
rect 20444 6740 20496 6792
rect 20536 6740 20588 6792
rect 18328 6604 18380 6656
rect 4250 6502 4302 6554
rect 4314 6502 4366 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 11955 6502 12007 6554
rect 12019 6502 12071 6554
rect 12083 6502 12135 6554
rect 12147 6502 12199 6554
rect 12211 6502 12263 6554
rect 19660 6502 19712 6554
rect 19724 6502 19776 6554
rect 19788 6502 19840 6554
rect 19852 6502 19904 6554
rect 19916 6502 19968 6554
rect 27365 6502 27417 6554
rect 27429 6502 27481 6554
rect 27493 6502 27545 6554
rect 27557 6502 27609 6554
rect 27621 6502 27673 6554
rect 10140 6400 10192 6452
rect 10416 6400 10468 6452
rect 10508 6400 10560 6452
rect 11152 6400 11204 6452
rect 11704 6400 11756 6452
rect 12716 6400 12768 6452
rect 13360 6400 13412 6452
rect 14372 6400 14424 6452
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 15660 6400 15712 6452
rect 10600 6332 10652 6384
rect 11428 6332 11480 6384
rect 12348 6332 12400 6384
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 11520 6264 11572 6316
rect 11704 6264 11756 6316
rect 13452 6332 13504 6384
rect 13544 6332 13596 6384
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 10692 6060 10744 6112
rect 12992 6128 13044 6180
rect 13728 6196 13780 6248
rect 14188 6196 14240 6248
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 12164 6060 12216 6112
rect 12624 6103 12676 6112
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 8102 5958 8154 6010
rect 8166 5958 8218 6010
rect 8230 5958 8282 6010
rect 8294 5958 8346 6010
rect 8358 5958 8410 6010
rect 15807 5958 15859 6010
rect 15871 5958 15923 6010
rect 15935 5958 15987 6010
rect 15999 5958 16051 6010
rect 16063 5958 16115 6010
rect 23512 5958 23564 6010
rect 23576 5958 23628 6010
rect 23640 5958 23692 6010
rect 23704 5958 23756 6010
rect 23768 5958 23820 6010
rect 31217 5958 31269 6010
rect 31281 5958 31333 6010
rect 31345 5958 31397 6010
rect 31409 5958 31461 6010
rect 31473 5958 31525 6010
rect 8760 5856 8812 5908
rect 10784 5856 10836 5908
rect 11060 5856 11112 5908
rect 12348 5856 12400 5908
rect 12624 5856 12676 5908
rect 12900 5856 12952 5908
rect 13820 5856 13872 5908
rect 14188 5856 14240 5908
rect 9772 5788 9824 5840
rect 11336 5831 11388 5840
rect 11336 5797 11345 5831
rect 11345 5797 11379 5831
rect 11379 5797 11388 5831
rect 11336 5788 11388 5797
rect 9404 5652 9456 5704
rect 12532 5720 12584 5772
rect 13084 5763 13136 5772
rect 13084 5729 13093 5763
rect 13093 5729 13127 5763
rect 13127 5729 13136 5763
rect 13084 5720 13136 5729
rect 8944 5584 8996 5636
rect 12072 5584 12124 5636
rect 8024 5516 8076 5568
rect 12164 5516 12216 5568
rect 4250 5414 4302 5466
rect 4314 5414 4366 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 11955 5414 12007 5466
rect 12019 5414 12071 5466
rect 12083 5414 12135 5466
rect 12147 5414 12199 5466
rect 12211 5414 12263 5466
rect 19660 5414 19712 5466
rect 19724 5414 19776 5466
rect 19788 5414 19840 5466
rect 19852 5414 19904 5466
rect 19916 5414 19968 5466
rect 27365 5414 27417 5466
rect 27429 5414 27481 5466
rect 27493 5414 27545 5466
rect 27557 5414 27609 5466
rect 27621 5414 27673 5466
rect 8102 4870 8154 4922
rect 8166 4870 8218 4922
rect 8230 4870 8282 4922
rect 8294 4870 8346 4922
rect 8358 4870 8410 4922
rect 15807 4870 15859 4922
rect 15871 4870 15923 4922
rect 15935 4870 15987 4922
rect 15999 4870 16051 4922
rect 16063 4870 16115 4922
rect 23512 4870 23564 4922
rect 23576 4870 23628 4922
rect 23640 4870 23692 4922
rect 23704 4870 23756 4922
rect 23768 4870 23820 4922
rect 31217 4870 31269 4922
rect 31281 4870 31333 4922
rect 31345 4870 31397 4922
rect 31409 4870 31461 4922
rect 31473 4870 31525 4922
rect 4250 4326 4302 4378
rect 4314 4326 4366 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 11955 4326 12007 4378
rect 12019 4326 12071 4378
rect 12083 4326 12135 4378
rect 12147 4326 12199 4378
rect 12211 4326 12263 4378
rect 19660 4326 19712 4378
rect 19724 4326 19776 4378
rect 19788 4326 19840 4378
rect 19852 4326 19904 4378
rect 19916 4326 19968 4378
rect 27365 4326 27417 4378
rect 27429 4326 27481 4378
rect 27493 4326 27545 4378
rect 27557 4326 27609 4378
rect 27621 4326 27673 4378
rect 14188 4088 14240 4140
rect 15292 4088 15344 4140
rect 8102 3782 8154 3834
rect 8166 3782 8218 3834
rect 8230 3782 8282 3834
rect 8294 3782 8346 3834
rect 8358 3782 8410 3834
rect 15807 3782 15859 3834
rect 15871 3782 15923 3834
rect 15935 3782 15987 3834
rect 15999 3782 16051 3834
rect 16063 3782 16115 3834
rect 23512 3782 23564 3834
rect 23576 3782 23628 3834
rect 23640 3782 23692 3834
rect 23704 3782 23756 3834
rect 23768 3782 23820 3834
rect 31217 3782 31269 3834
rect 31281 3782 31333 3834
rect 31345 3782 31397 3834
rect 31409 3782 31461 3834
rect 31473 3782 31525 3834
rect 9680 3476 9732 3528
rect 13912 3476 13964 3528
rect 4250 3238 4302 3290
rect 4314 3238 4366 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 11955 3238 12007 3290
rect 12019 3238 12071 3290
rect 12083 3238 12135 3290
rect 12147 3238 12199 3290
rect 12211 3238 12263 3290
rect 19660 3238 19712 3290
rect 19724 3238 19776 3290
rect 19788 3238 19840 3290
rect 19852 3238 19904 3290
rect 19916 3238 19968 3290
rect 27365 3238 27417 3290
rect 27429 3238 27481 3290
rect 27493 3238 27545 3290
rect 27557 3238 27609 3290
rect 27621 3238 27673 3290
rect 8102 2694 8154 2746
rect 8166 2694 8218 2746
rect 8230 2694 8282 2746
rect 8294 2694 8346 2746
rect 8358 2694 8410 2746
rect 15807 2694 15859 2746
rect 15871 2694 15923 2746
rect 15935 2694 15987 2746
rect 15999 2694 16051 2746
rect 16063 2694 16115 2746
rect 23512 2694 23564 2746
rect 23576 2694 23628 2746
rect 23640 2694 23692 2746
rect 23704 2694 23756 2746
rect 23768 2694 23820 2746
rect 31217 2694 31269 2746
rect 31281 2694 31333 2746
rect 31345 2694 31397 2746
rect 31409 2694 31461 2746
rect 31473 2694 31525 2746
rect 4250 2150 4302 2202
rect 4314 2150 4366 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 11955 2150 12007 2202
rect 12019 2150 12071 2202
rect 12083 2150 12135 2202
rect 12147 2150 12199 2202
rect 12211 2150 12263 2202
rect 19660 2150 19712 2202
rect 19724 2150 19776 2202
rect 19788 2150 19840 2202
rect 19852 2150 19904 2202
rect 19916 2150 19968 2202
rect 27365 2150 27417 2202
rect 27429 2150 27481 2202
rect 27493 2150 27545 2202
rect 27557 2150 27609 2202
rect 27621 2150 27673 2202
rect 8102 1606 8154 1658
rect 8166 1606 8218 1658
rect 8230 1606 8282 1658
rect 8294 1606 8346 1658
rect 8358 1606 8410 1658
rect 15807 1606 15859 1658
rect 15871 1606 15923 1658
rect 15935 1606 15987 1658
rect 15999 1606 16051 1658
rect 16063 1606 16115 1658
rect 23512 1606 23564 1658
rect 23576 1606 23628 1658
rect 23640 1606 23692 1658
rect 23704 1606 23756 1658
rect 23768 1606 23820 1658
rect 31217 1606 31269 1658
rect 31281 1606 31333 1658
rect 31345 1606 31397 1658
rect 31409 1606 31461 1658
rect 31473 1606 31525 1658
rect 4250 1062 4302 1114
rect 4314 1062 4366 1114
rect 4378 1062 4430 1114
rect 4442 1062 4494 1114
rect 4506 1062 4558 1114
rect 11955 1062 12007 1114
rect 12019 1062 12071 1114
rect 12083 1062 12135 1114
rect 12147 1062 12199 1114
rect 12211 1062 12263 1114
rect 19660 1062 19712 1114
rect 19724 1062 19776 1114
rect 19788 1062 19840 1114
rect 19852 1062 19904 1114
rect 19916 1062 19968 1114
rect 27365 1062 27417 1114
rect 27429 1062 27481 1114
rect 27493 1062 27545 1114
rect 27557 1062 27609 1114
rect 27621 1062 27673 1114
rect 8102 518 8154 570
rect 8166 518 8218 570
rect 8230 518 8282 570
rect 8294 518 8346 570
rect 8358 518 8410 570
rect 15807 518 15859 570
rect 15871 518 15923 570
rect 15935 518 15987 570
rect 15999 518 16051 570
rect 16063 518 16115 570
rect 23512 518 23564 570
rect 23576 518 23628 570
rect 23640 518 23692 570
rect 23704 518 23756 570
rect 23768 518 23820 570
rect 31217 518 31269 570
rect 31281 518 31333 570
rect 31345 518 31397 570
rect 31409 518 31461 570
rect 31473 518 31525 570
<< metal2 >>
rect 12898 19600 12954 20000
rect 13542 19600 13598 20000
rect 18050 19600 18106 20000
rect 18694 19600 18750 20000
rect 19338 19600 19394 20000
rect 19982 19600 20038 20000
rect 8102 19068 8410 19077
rect 8102 19066 8108 19068
rect 8164 19066 8188 19068
rect 8244 19066 8268 19068
rect 8324 19066 8348 19068
rect 8404 19066 8410 19068
rect 8164 19014 8166 19066
rect 8346 19014 8348 19066
rect 8102 19012 8108 19014
rect 8164 19012 8188 19014
rect 8244 19012 8268 19014
rect 8324 19012 8348 19014
rect 8404 19012 8410 19014
rect 8102 19003 8410 19012
rect 4250 18524 4558 18533
rect 4250 18522 4256 18524
rect 4312 18522 4336 18524
rect 4392 18522 4416 18524
rect 4472 18522 4496 18524
rect 4552 18522 4558 18524
rect 4312 18470 4314 18522
rect 4494 18470 4496 18522
rect 4250 18468 4256 18470
rect 4312 18468 4336 18470
rect 4392 18468 4416 18470
rect 4472 18468 4496 18470
rect 4552 18468 4558 18470
rect 4250 18459 4558 18468
rect 11955 18524 12263 18533
rect 11955 18522 11961 18524
rect 12017 18522 12041 18524
rect 12097 18522 12121 18524
rect 12177 18522 12201 18524
rect 12257 18522 12263 18524
rect 12017 18470 12019 18522
rect 12199 18470 12201 18522
rect 11955 18468 11961 18470
rect 12017 18468 12041 18470
rect 12097 18468 12121 18470
rect 12177 18468 12201 18470
rect 12257 18468 12263 18470
rect 11955 18459 12263 18468
rect 8102 17980 8410 17989
rect 8102 17978 8108 17980
rect 8164 17978 8188 17980
rect 8244 17978 8268 17980
rect 8324 17978 8348 17980
rect 8404 17978 8410 17980
rect 8164 17926 8166 17978
rect 8346 17926 8348 17978
rect 8102 17924 8108 17926
rect 8164 17924 8188 17926
rect 8244 17924 8268 17926
rect 8324 17924 8348 17926
rect 8404 17924 8410 17926
rect 8102 17915 8410 17924
rect 4250 17436 4558 17445
rect 4250 17434 4256 17436
rect 4312 17434 4336 17436
rect 4392 17434 4416 17436
rect 4472 17434 4496 17436
rect 4552 17434 4558 17436
rect 4312 17382 4314 17434
rect 4494 17382 4496 17434
rect 4250 17380 4256 17382
rect 4312 17380 4336 17382
rect 4392 17380 4416 17382
rect 4472 17380 4496 17382
rect 4552 17380 4558 17382
rect 4250 17371 4558 17380
rect 11955 17436 12263 17445
rect 11955 17434 11961 17436
rect 12017 17434 12041 17436
rect 12097 17434 12121 17436
rect 12177 17434 12201 17436
rect 12257 17434 12263 17436
rect 12017 17382 12019 17434
rect 12199 17382 12201 17434
rect 11955 17380 11961 17382
rect 12017 17380 12041 17382
rect 12097 17380 12121 17382
rect 12177 17380 12201 17382
rect 12257 17380 12263 17382
rect 11955 17371 12263 17380
rect 8102 16892 8410 16901
rect 8102 16890 8108 16892
rect 8164 16890 8188 16892
rect 8244 16890 8268 16892
rect 8324 16890 8348 16892
rect 8404 16890 8410 16892
rect 8164 16838 8166 16890
rect 8346 16838 8348 16890
rect 8102 16836 8108 16838
rect 8164 16836 8188 16838
rect 8244 16836 8268 16838
rect 8324 16836 8348 16838
rect 8404 16836 8410 16838
rect 8102 16827 8410 16836
rect 12912 16574 12940 19600
rect 13556 18970 13584 19600
rect 15807 19068 16115 19077
rect 15807 19066 15813 19068
rect 15869 19066 15893 19068
rect 15949 19066 15973 19068
rect 16029 19066 16053 19068
rect 16109 19066 16115 19068
rect 15869 19014 15871 19066
rect 16051 19014 16053 19066
rect 15807 19012 15813 19014
rect 15869 19012 15893 19014
rect 15949 19012 15973 19014
rect 16029 19012 16053 19014
rect 16109 19012 16115 19014
rect 15807 19003 16115 19012
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 12912 16546 13032 16574
rect 4250 16348 4558 16357
rect 4250 16346 4256 16348
rect 4312 16346 4336 16348
rect 4392 16346 4416 16348
rect 4472 16346 4496 16348
rect 4552 16346 4558 16348
rect 4312 16294 4314 16346
rect 4494 16294 4496 16346
rect 4250 16292 4256 16294
rect 4312 16292 4336 16294
rect 4392 16292 4416 16294
rect 4472 16292 4496 16294
rect 4552 16292 4558 16294
rect 4250 16283 4558 16292
rect 11955 16348 12263 16357
rect 11955 16346 11961 16348
rect 12017 16346 12041 16348
rect 12097 16346 12121 16348
rect 12177 16346 12201 16348
rect 12257 16346 12263 16348
rect 12017 16294 12019 16346
rect 12199 16294 12201 16346
rect 11955 16292 11961 16294
rect 12017 16292 12041 16294
rect 12097 16292 12121 16294
rect 12177 16292 12201 16294
rect 12257 16292 12263 16294
rect 11955 16283 12263 16292
rect 8102 15804 8410 15813
rect 8102 15802 8108 15804
rect 8164 15802 8188 15804
rect 8244 15802 8268 15804
rect 8324 15802 8348 15804
rect 8404 15802 8410 15804
rect 8164 15750 8166 15802
rect 8346 15750 8348 15802
rect 8102 15748 8108 15750
rect 8164 15748 8188 15750
rect 8244 15748 8268 15750
rect 8324 15748 8348 15750
rect 8404 15748 8410 15750
rect 8102 15739 8410 15748
rect 4250 15260 4558 15269
rect 4250 15258 4256 15260
rect 4312 15258 4336 15260
rect 4392 15258 4416 15260
rect 4472 15258 4496 15260
rect 4552 15258 4558 15260
rect 4312 15206 4314 15258
rect 4494 15206 4496 15258
rect 4250 15204 4256 15206
rect 4312 15204 4336 15206
rect 4392 15204 4416 15206
rect 4472 15204 4496 15206
rect 4552 15204 4558 15206
rect 4250 15195 4558 15204
rect 11955 15260 12263 15269
rect 11955 15258 11961 15260
rect 12017 15258 12041 15260
rect 12097 15258 12121 15260
rect 12177 15258 12201 15260
rect 12257 15258 12263 15260
rect 12017 15206 12019 15258
rect 12199 15206 12201 15258
rect 11955 15204 11961 15206
rect 12017 15204 12041 15206
rect 12097 15204 12121 15206
rect 12177 15204 12201 15206
rect 12257 15204 12263 15206
rect 11955 15195 12263 15204
rect 8102 14716 8410 14725
rect 8102 14714 8108 14716
rect 8164 14714 8188 14716
rect 8244 14714 8268 14716
rect 8324 14714 8348 14716
rect 8404 14714 8410 14716
rect 8164 14662 8166 14714
rect 8346 14662 8348 14714
rect 8102 14660 8108 14662
rect 8164 14660 8188 14662
rect 8244 14660 8268 14662
rect 8324 14660 8348 14662
rect 8404 14660 8410 14662
rect 8102 14651 8410 14660
rect 4250 14172 4558 14181
rect 4250 14170 4256 14172
rect 4312 14170 4336 14172
rect 4392 14170 4416 14172
rect 4472 14170 4496 14172
rect 4552 14170 4558 14172
rect 4312 14118 4314 14170
rect 4494 14118 4496 14170
rect 4250 14116 4256 14118
rect 4312 14116 4336 14118
rect 4392 14116 4416 14118
rect 4472 14116 4496 14118
rect 4552 14116 4558 14118
rect 4250 14107 4558 14116
rect 11955 14172 12263 14181
rect 11955 14170 11961 14172
rect 12017 14170 12041 14172
rect 12097 14170 12121 14172
rect 12177 14170 12201 14172
rect 12257 14170 12263 14172
rect 12017 14118 12019 14170
rect 12199 14118 12201 14170
rect 11955 14116 11961 14118
rect 12017 14116 12041 14118
rect 12097 14116 12121 14118
rect 12177 14116 12201 14118
rect 12257 14116 12263 14118
rect 11955 14107 12263 14116
rect 8102 13628 8410 13637
rect 8102 13626 8108 13628
rect 8164 13626 8188 13628
rect 8244 13626 8268 13628
rect 8324 13626 8348 13628
rect 8404 13626 8410 13628
rect 8164 13574 8166 13626
rect 8346 13574 8348 13626
rect 8102 13572 8108 13574
rect 8164 13572 8188 13574
rect 8244 13572 8268 13574
rect 8324 13572 8348 13574
rect 8404 13572 8410 13574
rect 8102 13563 8410 13572
rect 4250 13084 4558 13093
rect 4250 13082 4256 13084
rect 4312 13082 4336 13084
rect 4392 13082 4416 13084
rect 4472 13082 4496 13084
rect 4552 13082 4558 13084
rect 4312 13030 4314 13082
rect 4494 13030 4496 13082
rect 4250 13028 4256 13030
rect 4312 13028 4336 13030
rect 4392 13028 4416 13030
rect 4472 13028 4496 13030
rect 4552 13028 4558 13030
rect 4250 13019 4558 13028
rect 11955 13084 12263 13093
rect 11955 13082 11961 13084
rect 12017 13082 12041 13084
rect 12097 13082 12121 13084
rect 12177 13082 12201 13084
rect 12257 13082 12263 13084
rect 12017 13030 12019 13082
rect 12199 13030 12201 13082
rect 11955 13028 11961 13030
rect 12017 13028 12041 13030
rect 12097 13028 12121 13030
rect 12177 13028 12201 13030
rect 12257 13028 12263 13030
rect 11955 13019 12263 13028
rect 8102 12540 8410 12549
rect 8102 12538 8108 12540
rect 8164 12538 8188 12540
rect 8244 12538 8268 12540
rect 8324 12538 8348 12540
rect 8404 12538 8410 12540
rect 8164 12486 8166 12538
rect 8346 12486 8348 12538
rect 8102 12484 8108 12486
rect 8164 12484 8188 12486
rect 8244 12484 8268 12486
rect 8324 12484 8348 12486
rect 8404 12484 8410 12486
rect 8102 12475 8410 12484
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 4250 11996 4558 12005
rect 4250 11994 4256 11996
rect 4312 11994 4336 11996
rect 4392 11994 4416 11996
rect 4472 11994 4496 11996
rect 4552 11994 4558 11996
rect 4312 11942 4314 11994
rect 4494 11942 4496 11994
rect 4250 11940 4256 11942
rect 4312 11940 4336 11942
rect 4392 11940 4416 11942
rect 4472 11940 4496 11942
rect 4552 11940 4558 11942
rect 4250 11931 4558 11940
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8102 11452 8410 11461
rect 8102 11450 8108 11452
rect 8164 11450 8188 11452
rect 8244 11450 8268 11452
rect 8324 11450 8348 11452
rect 8404 11450 8410 11452
rect 8164 11398 8166 11450
rect 8346 11398 8348 11450
rect 8102 11396 8108 11398
rect 8164 11396 8188 11398
rect 8244 11396 8268 11398
rect 8324 11396 8348 11398
rect 8404 11396 8410 11398
rect 8102 11387 8410 11396
rect 4250 10908 4558 10917
rect 4250 10906 4256 10908
rect 4312 10906 4336 10908
rect 4392 10906 4416 10908
rect 4472 10906 4496 10908
rect 4552 10906 4558 10908
rect 4312 10854 4314 10906
rect 4494 10854 4496 10906
rect 4250 10852 4256 10854
rect 4312 10852 4336 10854
rect 4392 10852 4416 10854
rect 4472 10852 4496 10854
rect 4552 10852 4558 10854
rect 4250 10843 4558 10852
rect 8102 10364 8410 10373
rect 8102 10362 8108 10364
rect 8164 10362 8188 10364
rect 8244 10362 8268 10364
rect 8324 10362 8348 10364
rect 8404 10362 8410 10364
rect 8164 10310 8166 10362
rect 8346 10310 8348 10362
rect 8102 10308 8108 10310
rect 8164 10308 8188 10310
rect 8244 10308 8268 10310
rect 8324 10308 8348 10310
rect 8404 10308 8410 10310
rect 8102 10299 8410 10308
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 4250 9820 4558 9829
rect 4250 9818 4256 9820
rect 4312 9818 4336 9820
rect 4392 9818 4416 9820
rect 4472 9818 4496 9820
rect 4552 9818 4558 9820
rect 4312 9766 4314 9818
rect 4494 9766 4496 9818
rect 4250 9764 4256 9766
rect 4312 9764 4336 9766
rect 4392 9764 4416 9766
rect 4472 9764 4496 9766
rect 4552 9764 4558 9766
rect 4250 9755 4558 9764
rect 8220 9518 8248 9862
rect 8956 9586 8984 11698
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9048 10266 9076 10542
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8102 9276 8410 9285
rect 8102 9274 8108 9276
rect 8164 9274 8188 9276
rect 8244 9274 8268 9276
rect 8324 9274 8348 9276
rect 8404 9274 8410 9276
rect 8164 9222 8166 9274
rect 8346 9222 8348 9274
rect 8102 9220 8108 9222
rect 8164 9220 8188 9222
rect 8244 9220 8268 9222
rect 8324 9220 8348 9222
rect 8404 9220 8410 9222
rect 8102 9211 8410 9220
rect 8206 9072 8262 9081
rect 8772 9042 8800 9454
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8864 9042 8892 9318
rect 9140 9042 9168 9454
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9232 9058 9260 9386
rect 9324 9178 9352 11018
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 9518 9444 10406
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9508 9994 9536 10066
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9600 9761 9628 10066
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9586 9752 9642 9761
rect 9586 9687 9642 9696
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9232 9042 9352 9058
rect 9692 9042 9720 9862
rect 9784 9722 9812 10066
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 8206 9007 8208 9016
rect 8260 9007 8262 9016
rect 8760 9036 8812 9042
rect 8208 8978 8260 8984
rect 8760 8978 8812 8984
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 9128 9036 9180 9042
rect 9232 9036 9364 9042
rect 9232 9030 9312 9036
rect 9128 8978 9180 8984
rect 9312 8978 9364 8984
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 4250 8732 4558 8741
rect 4250 8730 4256 8732
rect 4312 8730 4336 8732
rect 4392 8730 4416 8732
rect 4472 8730 4496 8732
rect 4552 8730 4558 8732
rect 4312 8678 4314 8730
rect 4494 8678 4496 8730
rect 4250 8676 4256 8678
rect 4312 8676 4336 8678
rect 4392 8676 4416 8678
rect 4472 8676 4496 8678
rect 4552 8676 4558 8678
rect 4250 8667 4558 8676
rect 8036 8634 8064 8774
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 4250 7644 4558 7653
rect 4250 7642 4256 7644
rect 4312 7642 4336 7644
rect 4392 7642 4416 7644
rect 4472 7642 4496 7644
rect 4552 7642 4558 7644
rect 4312 7590 4314 7642
rect 4494 7590 4496 7642
rect 4250 7588 4256 7590
rect 4312 7588 4336 7590
rect 4392 7588 4416 7590
rect 4472 7588 4496 7590
rect 4552 7588 4558 7590
rect 4250 7579 4558 7588
rect 4250 6556 4558 6565
rect 4250 6554 4256 6556
rect 4312 6554 4336 6556
rect 4392 6554 4416 6556
rect 4472 6554 4496 6556
rect 4552 6554 4558 6556
rect 4312 6502 4314 6554
rect 4494 6502 4496 6554
rect 4250 6500 4256 6502
rect 4312 6500 4336 6502
rect 4392 6500 4416 6502
rect 4472 6500 4496 6502
rect 4552 6500 4558 6502
rect 4250 6491 4558 6500
rect 8036 5574 8064 8298
rect 8312 8294 8340 8910
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8392 8424 8444 8430
rect 8668 8424 8720 8430
rect 8444 8384 8524 8412
rect 8392 8366 8444 8372
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8102 8188 8410 8197
rect 8102 8186 8108 8188
rect 8164 8186 8188 8188
rect 8244 8186 8268 8188
rect 8324 8186 8348 8188
rect 8404 8186 8410 8188
rect 8164 8134 8166 8186
rect 8346 8134 8348 8186
rect 8102 8132 8108 8134
rect 8164 8132 8188 8134
rect 8244 8132 8268 8134
rect 8324 8132 8348 8134
rect 8404 8132 8410 8134
rect 8102 8123 8410 8132
rect 8496 8090 8524 8384
rect 8668 8366 8720 8372
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8102 7100 8410 7109
rect 8102 7098 8108 7100
rect 8164 7098 8188 7100
rect 8244 7098 8268 7100
rect 8324 7098 8348 7100
rect 8404 7098 8410 7100
rect 8164 7046 8166 7098
rect 8346 7046 8348 7098
rect 8102 7044 8108 7046
rect 8164 7044 8188 7046
rect 8244 7044 8268 7046
rect 8324 7044 8348 7046
rect 8404 7044 8410 7046
rect 8102 7035 8410 7044
rect 8588 6866 8616 8298
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8680 6730 8708 8366
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8102 6012 8410 6021
rect 8102 6010 8108 6012
rect 8164 6010 8188 6012
rect 8244 6010 8268 6012
rect 8324 6010 8348 6012
rect 8404 6010 8410 6012
rect 8164 5958 8166 6010
rect 8346 5958 8348 6010
rect 8102 5956 8108 5958
rect 8164 5956 8188 5958
rect 8244 5956 8268 5958
rect 8324 5956 8348 5958
rect 8404 5956 8410 5958
rect 8102 5947 8410 5956
rect 8772 5914 8800 8774
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8864 8022 8892 8434
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8956 5642 8984 8978
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8090 9076 8230
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9140 7886 9168 8978
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9312 8628 9364 8634
rect 9364 8588 9536 8616
rect 9312 8570 9364 8576
rect 9402 8528 9458 8537
rect 9402 8463 9404 8472
rect 9456 8463 9458 8472
rect 9404 8434 9456 8440
rect 9508 8430 9536 8588
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7478 9168 7822
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9416 5710 9444 8298
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9600 6746 9628 7958
rect 9692 6866 9720 8774
rect 9784 8430 9812 8774
rect 9876 8634 9904 9998
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9968 8430 9996 10542
rect 10520 10266 10548 11154
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10612 10266 10640 11018
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10266 10732 10950
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 8022 9812 8230
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9600 6718 9720 6746
rect 9692 6633 9720 6718
rect 9678 6624 9734 6633
rect 9678 6559 9734 6568
rect 9784 5846 9812 7686
rect 9968 7410 9996 7890
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 7002 9904 7278
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9876 6361 9904 6666
rect 9862 6352 9918 6361
rect 9968 6338 9996 7210
rect 10060 6769 10088 9862
rect 10140 9648 10192 9654
rect 10138 9616 10140 9625
rect 10192 9616 10194 9625
rect 10138 9551 10194 9560
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10152 7177 10180 8434
rect 10244 8430 10272 9930
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10244 7342 10272 8366
rect 10336 7886 10364 8366
rect 10428 8294 10456 10134
rect 10520 9994 10548 10202
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8430 10548 8978
rect 10612 8430 10640 9862
rect 10704 9722 10732 9998
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9178 10824 11494
rect 10888 11286 10916 11630
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10888 9178 10916 11222
rect 10980 10266 11008 12106
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11164 10266 11192 11494
rect 11256 11218 11284 11494
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9994 11008 10066
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11256 9722 11284 11154
rect 11440 10606 11468 11630
rect 11624 10742 11652 12378
rect 12268 12322 12296 12378
rect 12268 12306 12388 12322
rect 11704 12300 11756 12306
rect 12268 12300 12400 12306
rect 12268 12294 12348 12300
rect 11704 12242 11756 12248
rect 12348 12242 12400 12248
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 11716 11354 11744 12242
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 11808 11694 11836 12038
rect 11955 11996 12263 12005
rect 11955 11994 11961 11996
rect 12017 11994 12041 11996
rect 12097 11994 12121 11996
rect 12177 11994 12201 11996
rect 12257 11994 12263 11996
rect 12017 11942 12019 11994
rect 12199 11942 12201 11994
rect 11955 11940 11961 11942
rect 12017 11940 12041 11942
rect 12097 11940 12121 11942
rect 12177 11940 12201 11942
rect 12257 11940 12263 11942
rect 11955 11931 12263 11940
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10266 11376 10406
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10520 7954 10548 8366
rect 10704 8022 10732 8978
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10692 8016 10744 8022
rect 10612 7976 10692 8004
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10324 7880 10376 7886
rect 10376 7840 10456 7868
rect 10324 7822 10376 7828
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10232 7200 10284 7206
rect 10138 7168 10194 7177
rect 10232 7142 10284 7148
rect 10138 7103 10194 7112
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10046 6760 10102 6769
rect 10046 6695 10102 6704
rect 10152 6458 10180 6802
rect 10244 6497 10272 7142
rect 10428 6866 10456 7840
rect 10612 7274 10640 7976
rect 10692 7958 10744 7964
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10598 7168 10654 7177
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10230 6488 10286 6497
rect 10140 6452 10192 6458
rect 10428 6458 10456 6598
rect 10520 6458 10548 7142
rect 10598 7103 10654 7112
rect 10612 6866 10640 7103
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10230 6423 10286 6432
rect 10416 6452 10468 6458
rect 10140 6394 10192 6400
rect 10416 6394 10468 6400
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10600 6384 10652 6390
rect 9968 6332 10600 6338
rect 9968 6326 10652 6332
rect 9968 6310 10640 6326
rect 9862 6287 9918 6296
rect 10704 6118 10732 7686
rect 10796 7206 10824 8502
rect 10888 8498 10916 9114
rect 11150 8936 11206 8945
rect 11150 8871 11206 8880
rect 11244 8900 11296 8906
rect 11164 8838 11192 8871
rect 11244 8842 11296 8848
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10876 8288 10928 8294
rect 10980 8265 11008 8298
rect 10876 8230 10928 8236
rect 10966 8256 11022 8265
rect 10888 8022 10916 8230
rect 10966 8191 11022 8200
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10980 7750 11008 7890
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11072 7698 11100 8774
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 8401 11192 8570
rect 11150 8392 11206 8401
rect 11150 8327 11206 8336
rect 11150 8120 11206 8129
rect 11256 8090 11284 8842
rect 11150 8055 11152 8064
rect 11204 8055 11206 8064
rect 11244 8084 11296 8090
rect 11152 8026 11204 8032
rect 11244 8026 11296 8032
rect 11348 7970 11376 9454
rect 11440 8090 11468 9862
rect 11532 9586 11560 10066
rect 11624 10062 11652 10678
rect 11716 10266 11744 11290
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 9178 11560 9522
rect 11624 9518 11652 9862
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11532 9042 11560 9114
rect 11808 9081 11836 11494
rect 12176 11354 12204 11630
rect 12360 11354 12388 12038
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 11955 10908 12263 10917
rect 11955 10906 11961 10908
rect 12017 10906 12041 10908
rect 12097 10906 12121 10908
rect 12177 10906 12201 10908
rect 12257 10906 12263 10908
rect 12017 10854 12019 10906
rect 12199 10854 12201 10906
rect 11955 10852 11961 10854
rect 12017 10852 12041 10854
rect 12097 10852 12121 10854
rect 12177 10852 12201 10854
rect 12257 10852 12263 10854
rect 11955 10843 12263 10852
rect 12360 10470 12388 10950
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 11900 10305 11928 10406
rect 11886 10296 11942 10305
rect 11886 10231 11942 10240
rect 11955 9820 12263 9829
rect 11955 9818 11961 9820
rect 12017 9818 12041 9820
rect 12097 9818 12121 9820
rect 12177 9818 12201 9820
rect 12257 9818 12263 9820
rect 12017 9766 12019 9818
rect 12199 9766 12201 9818
rect 11955 9764 11961 9766
rect 12017 9764 12041 9766
rect 12097 9764 12121 9766
rect 12177 9764 12201 9766
rect 12257 9764 12263 9766
rect 11955 9755 12263 9764
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11794 9072 11850 9081
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11704 9036 11756 9042
rect 11794 9007 11850 9016
rect 11704 8978 11756 8984
rect 11716 8922 11744 8978
rect 11624 8894 11744 8922
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8498 11560 8774
rect 11624 8634 11652 8894
rect 11704 8832 11756 8838
rect 11900 8786 11928 9114
rect 11704 8774 11756 8780
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11716 8566 11744 8774
rect 11808 8758 11928 8786
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11624 7993 11652 8434
rect 11808 8378 11836 8758
rect 11955 8732 12263 8741
rect 11955 8730 11961 8732
rect 12017 8730 12041 8732
rect 12097 8730 12121 8732
rect 12177 8730 12201 8732
rect 12257 8730 12263 8732
rect 12017 8678 12019 8730
rect 12199 8678 12201 8730
rect 11955 8676 11961 8678
rect 12017 8676 12041 8678
rect 12097 8676 12121 8678
rect 12177 8676 12201 8678
rect 12257 8676 12263 8678
rect 11955 8667 12263 8676
rect 11716 8350 11836 8378
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12162 8392 12218 8401
rect 11610 7984 11666 7993
rect 11348 7942 11560 7970
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 10888 7342 10916 7686
rect 11072 7670 11284 7698
rect 11256 7546 11284 7670
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10980 7342 11008 7414
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10966 7032 11022 7041
rect 10966 6967 11022 6976
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10796 5914 10824 6802
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10888 6361 10916 6666
rect 10980 6662 11008 6967
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10874 6352 10930 6361
rect 10874 6287 10930 6296
rect 11072 5914 11100 7278
rect 11164 6458 11192 7482
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11256 6322 11284 6938
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11348 5846 11376 7210
rect 11440 7002 11468 7822
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11440 6390 11468 6938
rect 11532 6730 11560 7942
rect 11610 7919 11666 7928
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11518 6624 11574 6633
rect 11518 6559 11574 6568
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11532 6322 11560 6559
rect 11624 6338 11652 7686
rect 11716 7041 11744 8350
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11808 7562 11836 8230
rect 11900 8090 11928 8230
rect 11992 8129 12020 8366
rect 12218 8350 12296 8378
rect 12162 8327 12218 8336
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11978 8120 12034 8129
rect 11888 8084 11940 8090
rect 12084 8090 12112 8230
rect 11978 8055 12034 8064
rect 12072 8084 12124 8090
rect 11888 8026 11940 8032
rect 12072 8026 12124 8032
rect 12084 7818 12112 8026
rect 12164 7880 12216 7886
rect 12162 7848 12164 7857
rect 12216 7848 12218 7857
rect 12072 7812 12124 7818
rect 12268 7818 12296 8350
rect 12162 7783 12218 7792
rect 12256 7812 12308 7818
rect 12072 7754 12124 7760
rect 12256 7754 12308 7760
rect 12360 7750 12388 10406
rect 12452 9926 12480 10610
rect 12544 10130 12572 11154
rect 12636 10266 12664 12242
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11354 12940 11494
rect 13004 11354 13032 16546
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13096 11098 13124 11494
rect 13556 11354 13584 12038
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13648 11286 13676 18566
rect 15807 17980 16115 17989
rect 15807 17978 15813 17980
rect 15869 17978 15893 17980
rect 15949 17978 15973 17980
rect 16029 17978 16053 17980
rect 16109 17978 16115 17980
rect 15869 17926 15871 17978
rect 16051 17926 16053 17978
rect 15807 17924 15813 17926
rect 15869 17924 15893 17926
rect 15949 17924 15973 17926
rect 16029 17924 16053 17926
rect 16109 17924 16115 17926
rect 15807 17915 16115 17924
rect 15807 16892 16115 16901
rect 15807 16890 15813 16892
rect 15869 16890 15893 16892
rect 15949 16890 15973 16892
rect 16029 16890 16053 16892
rect 16109 16890 16115 16892
rect 15869 16838 15871 16890
rect 16051 16838 16053 16890
rect 15807 16836 15813 16838
rect 15869 16836 15893 16838
rect 15949 16836 15973 16838
rect 16029 16836 16053 16838
rect 16109 16836 16115 16838
rect 15807 16827 16115 16836
rect 18064 16574 18092 19600
rect 18708 16574 18736 19600
rect 19352 16574 19380 19600
rect 19660 18524 19968 18533
rect 19660 18522 19666 18524
rect 19722 18522 19746 18524
rect 19802 18522 19826 18524
rect 19882 18522 19906 18524
rect 19962 18522 19968 18524
rect 19722 18470 19724 18522
rect 19904 18470 19906 18522
rect 19660 18468 19666 18470
rect 19722 18468 19746 18470
rect 19802 18468 19826 18470
rect 19882 18468 19906 18470
rect 19962 18468 19968 18470
rect 19660 18459 19968 18468
rect 19660 17436 19968 17445
rect 19660 17434 19666 17436
rect 19722 17434 19746 17436
rect 19802 17434 19826 17436
rect 19882 17434 19906 17436
rect 19962 17434 19968 17436
rect 19722 17382 19724 17434
rect 19904 17382 19906 17434
rect 19660 17380 19666 17382
rect 19722 17380 19746 17382
rect 19802 17380 19826 17382
rect 19882 17380 19906 17382
rect 19962 17380 19968 17382
rect 19660 17371 19968 17380
rect 18064 16546 18552 16574
rect 18708 16546 18920 16574
rect 19352 16546 19472 16574
rect 15807 15804 16115 15813
rect 15807 15802 15813 15804
rect 15869 15802 15893 15804
rect 15949 15802 15973 15804
rect 16029 15802 16053 15804
rect 16109 15802 16115 15804
rect 15869 15750 15871 15802
rect 16051 15750 16053 15802
rect 15807 15748 15813 15750
rect 15869 15748 15893 15750
rect 15949 15748 15973 15750
rect 16029 15748 16053 15750
rect 16109 15748 16115 15750
rect 15807 15739 16115 15748
rect 15807 14716 16115 14725
rect 15807 14714 15813 14716
rect 15869 14714 15893 14716
rect 15949 14714 15973 14716
rect 16029 14714 16053 14716
rect 16109 14714 16115 14716
rect 15869 14662 15871 14714
rect 16051 14662 16053 14714
rect 15807 14660 15813 14662
rect 15869 14660 15893 14662
rect 15949 14660 15973 14662
rect 16029 14660 16053 14662
rect 16109 14660 16115 14662
rect 15807 14651 16115 14660
rect 15807 13628 16115 13637
rect 15807 13626 15813 13628
rect 15869 13626 15893 13628
rect 15949 13626 15973 13628
rect 16029 13626 16053 13628
rect 16109 13626 16115 13628
rect 15869 13574 15871 13626
rect 16051 13574 16053 13626
rect 15807 13572 15813 13574
rect 15869 13572 15893 13574
rect 15949 13572 15973 13574
rect 16029 13572 16053 13574
rect 16109 13572 16115 13574
rect 15807 13563 16115 13572
rect 15807 12540 16115 12549
rect 15807 12538 15813 12540
rect 15869 12538 15893 12540
rect 15949 12538 15973 12540
rect 16029 12538 16053 12540
rect 16109 12538 16115 12540
rect 15869 12486 15871 12538
rect 16051 12486 16053 12538
rect 15807 12484 15813 12486
rect 15869 12484 15893 12486
rect 15949 12484 15973 12486
rect 16029 12484 16053 12486
rect 16109 12484 16115 12486
rect 15807 12475 16115 12484
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13924 11898 13952 12038
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11354 13768 11630
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 14016 11218 14044 12038
rect 14108 11694 14136 12242
rect 14660 11898 14688 12242
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14108 11354 14136 11630
rect 15028 11354 15056 11766
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 13004 11070 13124 11098
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 14016 11098 14044 11154
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12728 10266 12756 10406
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12912 10062 12940 10406
rect 13004 10266 13032 11070
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10266 13124 10950
rect 13832 10810 13860 11086
rect 14016 11070 14136 11098
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13924 10810 13952 10950
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14108 10742 14136 11070
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10810 14228 10950
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13280 10554 13308 10610
rect 13188 10266 13216 10542
rect 13280 10526 13400 10554
rect 13372 10470 13400 10526
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13280 10266 13308 10406
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 12452 9382 12480 9862
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 13280 9178 13308 9386
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12544 8430 12572 8910
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 13096 8786 13124 8842
rect 13268 8832 13320 8838
rect 12636 8430 12664 8774
rect 13096 8758 13216 8786
rect 13268 8774 13320 8780
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 11955 7644 12263 7653
rect 11955 7642 11961 7644
rect 12017 7642 12041 7644
rect 12097 7642 12121 7644
rect 12177 7642 12201 7644
rect 12257 7642 12263 7644
rect 12017 7590 12019 7642
rect 12199 7590 12201 7642
rect 11955 7588 11961 7590
rect 12017 7588 12041 7590
rect 12097 7588 12121 7590
rect 12177 7588 12201 7590
rect 12257 7588 12263 7590
rect 11955 7579 12263 7588
rect 11808 7534 11928 7562
rect 11702 7032 11758 7041
rect 11900 7002 11928 7534
rect 12452 7478 12480 7822
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 11702 6967 11704 6976
rect 11756 6967 11758 6976
rect 11888 6996 11940 7002
rect 11704 6938 11756 6944
rect 11888 6938 11940 6944
rect 12544 6934 12572 7754
rect 12636 7342 12664 8230
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12532 6928 12584 6934
rect 11886 6896 11942 6905
rect 11942 6866 12020 6882
rect 12532 6870 12584 6876
rect 11942 6860 12032 6866
rect 11942 6854 11980 6860
rect 11886 6831 11942 6840
rect 11980 6802 12032 6808
rect 12162 6760 12218 6769
rect 12636 6746 12664 7142
rect 12162 6695 12164 6704
rect 12216 6695 12218 6704
rect 12452 6718 12664 6746
rect 12164 6666 12216 6672
rect 11704 6656 11756 6662
rect 11702 6624 11704 6633
rect 11756 6624 11758 6633
rect 11702 6559 11758 6568
rect 11955 6556 12263 6565
rect 11955 6554 11961 6556
rect 12017 6554 12041 6556
rect 12097 6554 12121 6556
rect 12177 6554 12201 6556
rect 12257 6554 12263 6556
rect 12017 6502 12019 6554
rect 12199 6502 12201 6554
rect 11955 6500 11961 6502
rect 12017 6500 12041 6502
rect 12097 6500 12121 6502
rect 12177 6500 12201 6502
rect 12257 6500 12263 6502
rect 11702 6488 11758 6497
rect 11955 6491 12263 6500
rect 11702 6423 11704 6432
rect 11756 6423 11758 6432
rect 11704 6394 11756 6400
rect 12348 6384 12400 6390
rect 11624 6322 11744 6338
rect 12348 6326 12400 6332
rect 11520 6316 11572 6322
rect 11624 6316 11756 6322
rect 11624 6310 11704 6316
rect 11520 6258 11572 6264
rect 11704 6258 11756 6264
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 12084 5642 12112 6054
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12176 5574 12204 6054
rect 12360 5914 12388 6326
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 4250 5468 4558 5477
rect 4250 5466 4256 5468
rect 4312 5466 4336 5468
rect 4392 5466 4416 5468
rect 4472 5466 4496 5468
rect 4552 5466 4558 5468
rect 4312 5414 4314 5466
rect 4494 5414 4496 5466
rect 4250 5412 4256 5414
rect 4312 5412 4336 5414
rect 4392 5412 4416 5414
rect 4472 5412 4496 5414
rect 4552 5412 4558 5414
rect 4250 5403 4558 5412
rect 11955 5468 12263 5477
rect 11955 5466 11961 5468
rect 12017 5466 12041 5468
rect 12097 5466 12121 5468
rect 12177 5466 12201 5468
rect 12257 5466 12263 5468
rect 12017 5414 12019 5466
rect 12199 5414 12201 5466
rect 11955 5412 11961 5414
rect 12017 5412 12041 5414
rect 12097 5412 12121 5414
rect 12177 5412 12201 5414
rect 12257 5412 12263 5414
rect 11955 5403 12263 5412
rect 8102 4924 8410 4933
rect 8102 4922 8108 4924
rect 8164 4922 8188 4924
rect 8244 4922 8268 4924
rect 8324 4922 8348 4924
rect 8404 4922 8410 4924
rect 8164 4870 8166 4922
rect 8346 4870 8348 4922
rect 8102 4868 8108 4870
rect 8164 4868 8188 4870
rect 8244 4868 8268 4870
rect 8324 4868 8348 4870
rect 8404 4868 8410 4870
rect 8102 4859 8410 4868
rect 4250 4380 4558 4389
rect 4250 4378 4256 4380
rect 4312 4378 4336 4380
rect 4392 4378 4416 4380
rect 4472 4378 4496 4380
rect 4552 4378 4558 4380
rect 4312 4326 4314 4378
rect 4494 4326 4496 4378
rect 4250 4324 4256 4326
rect 4312 4324 4336 4326
rect 4392 4324 4416 4326
rect 4472 4324 4496 4326
rect 4552 4324 4558 4326
rect 4250 4315 4558 4324
rect 11955 4380 12263 4389
rect 11955 4378 11961 4380
rect 12017 4378 12041 4380
rect 12097 4378 12121 4380
rect 12177 4378 12201 4380
rect 12257 4378 12263 4380
rect 12017 4326 12019 4378
rect 12199 4326 12201 4378
rect 11955 4324 11961 4326
rect 12017 4324 12041 4326
rect 12097 4324 12121 4326
rect 12177 4324 12201 4326
rect 12257 4324 12263 4326
rect 11955 4315 12263 4324
rect 8102 3836 8410 3845
rect 8102 3834 8108 3836
rect 8164 3834 8188 3836
rect 8244 3834 8268 3836
rect 8324 3834 8348 3836
rect 8404 3834 8410 3836
rect 8164 3782 8166 3834
rect 8346 3782 8348 3834
rect 8102 3780 8108 3782
rect 8164 3780 8188 3782
rect 8244 3780 8268 3782
rect 8324 3780 8348 3782
rect 8404 3780 8410 3782
rect 8102 3771 8410 3780
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 4250 3292 4558 3301
rect 4250 3290 4256 3292
rect 4312 3290 4336 3292
rect 4392 3290 4416 3292
rect 4472 3290 4496 3292
rect 4552 3290 4558 3292
rect 4312 3238 4314 3290
rect 4494 3238 4496 3290
rect 4250 3236 4256 3238
rect 4312 3236 4336 3238
rect 4392 3236 4416 3238
rect 4472 3236 4496 3238
rect 4552 3236 4558 3238
rect 4250 3227 4558 3236
rect 8102 2748 8410 2757
rect 8102 2746 8108 2748
rect 8164 2746 8188 2748
rect 8244 2746 8268 2748
rect 8324 2746 8348 2748
rect 8404 2746 8410 2748
rect 8164 2694 8166 2746
rect 8346 2694 8348 2746
rect 8102 2692 8108 2694
rect 8164 2692 8188 2694
rect 8244 2692 8268 2694
rect 8324 2692 8348 2694
rect 8404 2692 8410 2694
rect 8102 2683 8410 2692
rect 4250 2204 4558 2213
rect 4250 2202 4256 2204
rect 4312 2202 4336 2204
rect 4392 2202 4416 2204
rect 4472 2202 4496 2204
rect 4552 2202 4558 2204
rect 4312 2150 4314 2202
rect 4494 2150 4496 2202
rect 4250 2148 4256 2150
rect 4312 2148 4336 2150
rect 4392 2148 4416 2150
rect 4472 2148 4496 2150
rect 4552 2148 4558 2150
rect 4250 2139 4558 2148
rect 8102 1660 8410 1669
rect 8102 1658 8108 1660
rect 8164 1658 8188 1660
rect 8244 1658 8268 1660
rect 8324 1658 8348 1660
rect 8404 1658 8410 1660
rect 8164 1606 8166 1658
rect 8346 1606 8348 1658
rect 8102 1604 8108 1606
rect 8164 1604 8188 1606
rect 8244 1604 8268 1606
rect 8324 1604 8348 1606
rect 8404 1604 8410 1606
rect 8102 1595 8410 1604
rect 4250 1116 4558 1125
rect 4250 1114 4256 1116
rect 4312 1114 4336 1116
rect 4392 1114 4416 1116
rect 4472 1114 4496 1116
rect 4552 1114 4558 1116
rect 4312 1062 4314 1114
rect 4494 1062 4496 1114
rect 4250 1060 4256 1062
rect 4312 1060 4336 1062
rect 4392 1060 4416 1062
rect 4472 1060 4496 1062
rect 4552 1060 4558 1062
rect 4250 1051 4558 1060
rect 8102 572 8410 581
rect 8102 570 8108 572
rect 8164 570 8188 572
rect 8244 570 8268 572
rect 8324 570 8348 572
rect 8404 570 8410 572
rect 8164 518 8166 570
rect 8346 518 8348 570
rect 8102 516 8108 518
rect 8164 516 8188 518
rect 8244 516 8268 518
rect 8324 516 8348 518
rect 8404 516 8410 518
rect 8102 507 8410 516
rect 9692 400 9720 3470
rect 11955 3292 12263 3301
rect 11955 3290 11961 3292
rect 12017 3290 12041 3292
rect 12097 3290 12121 3292
rect 12177 3290 12201 3292
rect 12257 3290 12263 3292
rect 12017 3238 12019 3290
rect 12199 3238 12201 3290
rect 11955 3236 11961 3238
rect 12017 3236 12041 3238
rect 12097 3236 12121 3238
rect 12177 3236 12201 3238
rect 12257 3236 12263 3238
rect 11955 3227 12263 3236
rect 12452 3210 12480 6718
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 5778 12572 6598
rect 12728 6458 12756 7482
rect 12820 7342 12848 8502
rect 13096 8430 13124 8570
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 13082 8256 13138 8265
rect 12912 8022 12940 8230
rect 13082 8191 13138 8200
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12990 7984 13046 7993
rect 12990 7919 13046 7928
rect 12898 7848 12954 7857
rect 12898 7783 12954 7792
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12912 7002 12940 7783
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12806 6896 12862 6905
rect 12806 6831 12862 6840
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12820 6254 12848 6831
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 13004 6186 13032 7919
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12636 5914 12664 6054
rect 12912 5914 12940 6054
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13096 5778 13124 8191
rect 13188 6866 13216 8758
rect 13280 8566 13308 8774
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13556 8498 13584 9862
rect 13740 9518 13768 10610
rect 15120 10606 15148 11154
rect 15212 10810 15240 11562
rect 15396 11558 15424 12038
rect 16316 11898 16344 12242
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 16304 11688 16356 11694
rect 16488 11688 16540 11694
rect 16356 11648 16488 11676
rect 16304 11630 16356 11636
rect 16856 11688 16908 11694
rect 16488 11630 16540 11636
rect 16776 11648 16856 11676
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15396 10674 15424 11494
rect 15488 10810 15516 11630
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 15807 11452 16115 11461
rect 15807 11450 15813 11452
rect 15869 11450 15893 11452
rect 15949 11450 15973 11452
rect 16029 11450 16053 11452
rect 16109 11450 16115 11452
rect 15869 11398 15871 11450
rect 16051 11398 16053 11450
rect 15807 11396 15813 11398
rect 15869 11396 15893 11398
rect 15949 11396 15973 11398
rect 16029 11396 16053 11398
rect 16109 11396 16115 11398
rect 15807 11387 16115 11396
rect 16224 11234 16252 11494
rect 16500 11354 16528 11630
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16224 11206 16436 11234
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15580 10690 15608 11086
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16224 10810 16252 10950
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 15488 10674 15608 10690
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15476 10668 15608 10674
rect 15528 10662 15608 10668
rect 15476 10610 15528 10616
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 13832 10266 13860 10542
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14016 9518 14044 10474
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14292 10266 14320 10406
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14384 9518 14412 10406
rect 15488 9602 15516 10610
rect 15807 10364 16115 10373
rect 15807 10362 15813 10364
rect 15869 10362 15893 10364
rect 15949 10362 15973 10364
rect 16029 10362 16053 10364
rect 16109 10362 16115 10364
rect 15869 10310 15871 10362
rect 16051 10310 16053 10362
rect 15807 10308 15813 10310
rect 15869 10308 15893 10310
rect 15949 10308 15973 10310
rect 16029 10308 16053 10310
rect 16109 10308 16115 10310
rect 15807 10299 16115 10308
rect 16316 10282 16344 11018
rect 16408 11014 16436 11206
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16592 10470 16620 11154
rect 16776 11150 16804 11648
rect 16856 11630 16908 11636
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18432 11218 18460 11630
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16224 10254 16344 10282
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9761 15608 9862
rect 15566 9752 15622 9761
rect 15566 9687 15622 9696
rect 15292 9580 15344 9586
rect 15488 9574 15608 9602
rect 15292 9522 15344 9528
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7546 13308 7686
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13372 6458 13400 7414
rect 13464 7002 13492 8026
rect 13556 7410 13584 8434
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13464 6390 13492 6938
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13556 6390 13584 6870
rect 13648 6866 13676 8910
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13832 8022 13860 8570
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13740 6254 13768 7142
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13832 5914 13860 7210
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13924 3534 13952 8978
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 14016 8022 14044 8842
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14094 8120 14150 8129
rect 14292 8106 14320 8298
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14150 8078 14320 8106
rect 14384 8090 14412 8230
rect 14660 8090 14688 8774
rect 15304 8498 15332 9522
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 9110 15424 9318
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15580 8922 15608 9574
rect 15672 9178 15700 10066
rect 15807 9276 16115 9285
rect 15807 9274 15813 9276
rect 15869 9274 15893 9276
rect 15949 9274 15973 9276
rect 16029 9274 16053 9276
rect 16109 9274 16115 9276
rect 15869 9222 15871 9274
rect 16051 9222 16053 9274
rect 15807 9220 15813 9222
rect 15869 9220 15893 9222
rect 15949 9220 15973 9222
rect 16029 9220 16053 9222
rect 16109 9220 16115 9222
rect 15807 9211 16115 9220
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15672 9042 15700 9114
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15764 8922 15792 8978
rect 15580 8894 15792 8922
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14094 8055 14150 8064
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14016 7002 14044 7754
rect 14108 7342 14136 7890
rect 14200 7546 14228 7890
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14004 6860 14056 6866
rect 14108 6848 14136 6938
rect 14056 6820 14136 6848
rect 14004 6802 14056 6808
rect 14200 6254 14228 7482
rect 14292 6798 14320 8078
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14384 7002 14412 7890
rect 15028 7410 15056 8434
rect 16224 8430 16252 10254
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16316 9178 16344 10066
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16408 9722 16436 9862
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16500 9518 16528 10406
rect 16592 10266 16620 10406
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16684 10146 16712 10542
rect 16592 10118 16712 10146
rect 16592 9654 16620 10118
rect 16776 10010 16804 10610
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17328 10130 17356 10406
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 16684 9982 16804 10010
rect 16684 9674 16712 9982
rect 16580 9648 16632 9654
rect 16684 9646 17080 9674
rect 16580 9590 16632 9596
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16592 8974 16620 9590
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16592 8430 16620 8910
rect 16868 8498 16896 8978
rect 17052 8838 17080 9646
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 15212 7970 15240 8230
rect 15672 8090 15700 8230
rect 15807 8188 16115 8197
rect 15807 8186 15813 8188
rect 15869 8186 15893 8188
rect 15949 8186 15973 8188
rect 16029 8186 16053 8188
rect 16109 8186 16115 8188
rect 15869 8134 15871 8186
rect 16051 8134 16053 8186
rect 15807 8132 15813 8134
rect 15869 8132 15893 8134
rect 15949 8132 15973 8134
rect 16029 8132 16053 8134
rect 16109 8132 16115 8134
rect 15807 8123 16115 8132
rect 16316 8090 16344 8230
rect 16592 8090 16620 8230
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 15108 7948 15160 7954
rect 15212 7942 15332 7970
rect 15108 7890 15160 7896
rect 15120 7546 15148 7890
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14384 6458 14412 6938
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5914 14228 6054
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 12360 3182 12480 3210
rect 11955 2204 12263 2213
rect 11955 2202 11961 2204
rect 12017 2202 12041 2204
rect 12097 2202 12121 2204
rect 12177 2202 12201 2204
rect 12257 2202 12263 2204
rect 12017 2150 12019 2202
rect 12199 2150 12201 2202
rect 11955 2148 11961 2150
rect 12017 2148 12041 2150
rect 12097 2148 12121 2150
rect 12177 2148 12201 2150
rect 12257 2148 12263 2150
rect 11955 2139 12263 2148
rect 11955 1116 12263 1125
rect 11955 1114 11961 1116
rect 12017 1114 12041 1116
rect 12097 1114 12121 1116
rect 12177 1114 12201 1116
rect 12257 1114 12263 1116
rect 12017 1062 12019 1114
rect 12199 1062 12201 1114
rect 11955 1060 11961 1062
rect 12017 1060 12041 1062
rect 12097 1060 12121 1062
rect 12177 1060 12201 1062
rect 12257 1060 12263 1062
rect 11955 1051 12263 1060
rect 12360 898 12388 3182
rect 12268 870 12388 898
rect 12268 400 12296 870
rect 14200 400 14228 4082
rect 14476 2774 14504 6938
rect 14936 6934 14964 7142
rect 15120 7002 15148 7482
rect 15212 7002 15240 7822
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14568 6458 14596 6666
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 15120 6254 15148 6598
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15304 4146 15332 7942
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7750 15516 7822
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15396 7290 15424 7686
rect 15396 7262 15516 7290
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 6934 15424 7142
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15488 6730 15516 7262
rect 15580 6934 15608 8026
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15672 6458 15700 7210
rect 15807 7100 16115 7109
rect 15807 7098 15813 7100
rect 15869 7098 15893 7100
rect 15949 7098 15973 7100
rect 16029 7098 16053 7100
rect 16109 7098 16115 7100
rect 15869 7046 15871 7098
rect 16051 7046 16053 7098
rect 15807 7044 15813 7046
rect 15869 7044 15893 7046
rect 15949 7044 15973 7046
rect 16029 7044 16053 7046
rect 16109 7044 16115 7046
rect 15807 7035 16115 7044
rect 16316 7002 16344 7890
rect 16684 7886 16712 8230
rect 16868 7954 16896 8434
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16592 7002 16620 7754
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7546 16712 7686
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16960 7478 16988 8366
rect 17052 8344 17080 8774
rect 17144 8634 17172 9454
rect 17512 9382 17540 10406
rect 17604 9722 17632 10406
rect 17880 10062 17908 10610
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17236 8362 17264 9318
rect 17696 8566 17724 9318
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17788 8430 17816 9930
rect 17880 9586 17908 9998
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17880 8974 17908 9522
rect 17972 9450 18000 9862
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8430 17908 8910
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17132 8356 17184 8362
rect 17052 8316 17132 8344
rect 17132 8298 17184 8304
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 7002 16712 7210
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16960 6934 16988 7414
rect 17144 7342 17172 8298
rect 17236 8090 17264 8298
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15807 6012 16115 6021
rect 15807 6010 15813 6012
rect 15869 6010 15893 6012
rect 15949 6010 15973 6012
rect 16029 6010 16053 6012
rect 16109 6010 16115 6012
rect 15869 5958 15871 6010
rect 16051 5958 16053 6010
rect 15807 5956 15813 5958
rect 15869 5956 15893 5958
rect 15949 5956 15973 5958
rect 16029 5956 16053 5958
rect 16109 5956 16115 5958
rect 15807 5947 16115 5956
rect 15807 4924 16115 4933
rect 15807 4922 15813 4924
rect 15869 4922 15893 4924
rect 15949 4922 15973 4924
rect 16029 4922 16053 4924
rect 16109 4922 16115 4924
rect 15869 4870 15871 4922
rect 16051 4870 16053 4922
rect 15807 4868 15813 4870
rect 15869 4868 15893 4870
rect 15949 4868 15973 4870
rect 16029 4868 16053 4870
rect 16109 4868 16115 4870
rect 15807 4859 16115 4868
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15474 4040 15530 4049
rect 15474 3975 15530 3984
rect 14384 2746 14504 2774
rect 9678 0 9734 400
rect 12254 0 12310 400
rect 14186 0 14242 400
rect 14384 354 14412 2746
rect 14752 462 14872 490
rect 14752 354 14780 462
rect 14844 400 14872 462
rect 15488 400 15516 3975
rect 15807 3836 16115 3845
rect 15807 3834 15813 3836
rect 15869 3834 15893 3836
rect 15949 3834 15973 3836
rect 16029 3834 16053 3836
rect 16109 3834 16115 3836
rect 15869 3782 15871 3834
rect 16051 3782 16053 3834
rect 15807 3780 15813 3782
rect 15869 3780 15893 3782
rect 15949 3780 15973 3782
rect 16029 3780 16053 3782
rect 16109 3780 16115 3782
rect 15807 3771 16115 3780
rect 15807 2748 16115 2757
rect 15807 2746 15813 2748
rect 15869 2746 15893 2748
rect 15949 2746 15973 2748
rect 16029 2746 16053 2748
rect 16109 2746 16115 2748
rect 15869 2694 15871 2746
rect 16051 2694 16053 2746
rect 15807 2692 15813 2694
rect 15869 2692 15893 2694
rect 15949 2692 15973 2694
rect 16029 2692 16053 2694
rect 16109 2692 16115 2694
rect 15807 2683 16115 2692
rect 15807 1660 16115 1669
rect 15807 1658 15813 1660
rect 15869 1658 15893 1660
rect 15949 1658 15973 1660
rect 16029 1658 16053 1660
rect 16109 1658 16115 1660
rect 15869 1606 15871 1658
rect 16051 1606 16053 1658
rect 15807 1604 15813 1606
rect 15869 1604 15893 1606
rect 15949 1604 15973 1606
rect 16029 1604 16053 1606
rect 16109 1604 16115 1606
rect 15807 1595 16115 1604
rect 15807 572 16115 581
rect 15807 570 15813 572
rect 15869 570 15893 572
rect 15949 570 15973 572
rect 16029 570 16053 572
rect 16109 570 16115 572
rect 15869 518 15871 570
rect 16051 518 16053 570
rect 15807 516 15813 518
rect 15869 516 15893 518
rect 15949 516 15973 518
rect 16029 516 16053 518
rect 16109 516 16115 518
rect 15807 507 16115 516
rect 16776 462 16896 490
rect 16776 400 16804 462
rect 14384 326 14780 354
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16762 0 16818 400
rect 16868 354 16896 462
rect 17052 354 17080 7142
rect 17236 6866 17264 7142
rect 17328 6866 17356 7278
rect 17420 6866 17448 8298
rect 17972 7886 18000 8774
rect 18064 8566 18092 10542
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 8566 18184 10406
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18248 8430 18276 10474
rect 18432 10130 18460 11154
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18432 9722 18460 10066
rect 18420 9716 18472 9722
rect 18340 9664 18420 9674
rect 18340 9658 18472 9664
rect 18340 9646 18460 9658
rect 18524 9654 18552 16546
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18800 11694 18828 12038
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18616 10606 18644 10950
rect 18892 10810 18920 16546
rect 19444 12374 19472 16546
rect 19660 16348 19968 16357
rect 19660 16346 19666 16348
rect 19722 16346 19746 16348
rect 19802 16346 19826 16348
rect 19882 16346 19906 16348
rect 19962 16346 19968 16348
rect 19722 16294 19724 16346
rect 19904 16294 19906 16346
rect 19660 16292 19666 16294
rect 19722 16292 19746 16294
rect 19802 16292 19826 16294
rect 19882 16292 19906 16294
rect 19962 16292 19968 16294
rect 19660 16283 19968 16292
rect 19660 15260 19968 15269
rect 19660 15258 19666 15260
rect 19722 15258 19746 15260
rect 19802 15258 19826 15260
rect 19882 15258 19906 15260
rect 19962 15258 19968 15260
rect 19722 15206 19724 15258
rect 19904 15206 19906 15258
rect 19660 15204 19666 15206
rect 19722 15204 19746 15206
rect 19802 15204 19826 15206
rect 19882 15204 19906 15206
rect 19962 15204 19968 15206
rect 19660 15195 19968 15204
rect 19660 14172 19968 14181
rect 19660 14170 19666 14172
rect 19722 14170 19746 14172
rect 19802 14170 19826 14172
rect 19882 14170 19906 14172
rect 19962 14170 19968 14172
rect 19722 14118 19724 14170
rect 19904 14118 19906 14170
rect 19660 14116 19666 14118
rect 19722 14116 19746 14118
rect 19802 14116 19826 14118
rect 19882 14116 19906 14118
rect 19962 14116 19968 14118
rect 19660 14107 19968 14116
rect 19660 13084 19968 13093
rect 19660 13082 19666 13084
rect 19722 13082 19746 13084
rect 19802 13082 19826 13084
rect 19882 13082 19906 13084
rect 19962 13082 19968 13084
rect 19722 13030 19724 13082
rect 19904 13030 19906 13082
rect 19660 13028 19666 13030
rect 19722 13028 19746 13030
rect 19802 13028 19826 13030
rect 19882 13028 19906 13030
rect 19962 13028 19968 13030
rect 19660 13019 19968 13028
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19660 11996 19968 12005
rect 19660 11994 19666 11996
rect 19722 11994 19746 11996
rect 19802 11994 19826 11996
rect 19882 11994 19906 11996
rect 19962 11994 19968 11996
rect 19722 11942 19724 11994
rect 19904 11942 19906 11994
rect 19660 11940 19666 11942
rect 19722 11940 19746 11942
rect 19802 11940 19826 11942
rect 19882 11940 19906 11942
rect 19962 11940 19968 11942
rect 19660 11931 19968 11940
rect 19996 11336 20024 19600
rect 23512 19068 23820 19077
rect 23512 19066 23518 19068
rect 23574 19066 23598 19068
rect 23654 19066 23678 19068
rect 23734 19066 23758 19068
rect 23814 19066 23820 19068
rect 23574 19014 23576 19066
rect 23756 19014 23758 19066
rect 23512 19012 23518 19014
rect 23574 19012 23598 19014
rect 23654 19012 23678 19014
rect 23734 19012 23758 19014
rect 23814 19012 23820 19014
rect 23512 19003 23820 19012
rect 31217 19068 31525 19077
rect 31217 19066 31223 19068
rect 31279 19066 31303 19068
rect 31359 19066 31383 19068
rect 31439 19066 31463 19068
rect 31519 19066 31525 19068
rect 31279 19014 31281 19066
rect 31461 19014 31463 19066
rect 31217 19012 31223 19014
rect 31279 19012 31303 19014
rect 31359 19012 31383 19014
rect 31439 19012 31463 19014
rect 31519 19012 31525 19014
rect 31217 19003 31525 19012
rect 27365 18524 27673 18533
rect 27365 18522 27371 18524
rect 27427 18522 27451 18524
rect 27507 18522 27531 18524
rect 27587 18522 27611 18524
rect 27667 18522 27673 18524
rect 27427 18470 27429 18522
rect 27609 18470 27611 18522
rect 27365 18468 27371 18470
rect 27427 18468 27451 18470
rect 27507 18468 27531 18470
rect 27587 18468 27611 18470
rect 27667 18468 27673 18470
rect 27365 18459 27673 18468
rect 23512 17980 23820 17989
rect 23512 17978 23518 17980
rect 23574 17978 23598 17980
rect 23654 17978 23678 17980
rect 23734 17978 23758 17980
rect 23814 17978 23820 17980
rect 23574 17926 23576 17978
rect 23756 17926 23758 17978
rect 23512 17924 23518 17926
rect 23574 17924 23598 17926
rect 23654 17924 23678 17926
rect 23734 17924 23758 17926
rect 23814 17924 23820 17926
rect 23512 17915 23820 17924
rect 31217 17980 31525 17989
rect 31217 17978 31223 17980
rect 31279 17978 31303 17980
rect 31359 17978 31383 17980
rect 31439 17978 31463 17980
rect 31519 17978 31525 17980
rect 31279 17926 31281 17978
rect 31461 17926 31463 17978
rect 31217 17924 31223 17926
rect 31279 17924 31303 17926
rect 31359 17924 31383 17926
rect 31439 17924 31463 17926
rect 31519 17924 31525 17926
rect 31217 17915 31525 17924
rect 27365 17436 27673 17445
rect 27365 17434 27371 17436
rect 27427 17434 27451 17436
rect 27507 17434 27531 17436
rect 27587 17434 27611 17436
rect 27667 17434 27673 17436
rect 27427 17382 27429 17434
rect 27609 17382 27611 17434
rect 27365 17380 27371 17382
rect 27427 17380 27451 17382
rect 27507 17380 27531 17382
rect 27587 17380 27611 17382
rect 27667 17380 27673 17382
rect 27365 17371 27673 17380
rect 23512 16892 23820 16901
rect 23512 16890 23518 16892
rect 23574 16890 23598 16892
rect 23654 16890 23678 16892
rect 23734 16890 23758 16892
rect 23814 16890 23820 16892
rect 23574 16838 23576 16890
rect 23756 16838 23758 16890
rect 23512 16836 23518 16838
rect 23574 16836 23598 16838
rect 23654 16836 23678 16838
rect 23734 16836 23758 16838
rect 23814 16836 23820 16838
rect 23512 16827 23820 16836
rect 31217 16892 31525 16901
rect 31217 16890 31223 16892
rect 31279 16890 31303 16892
rect 31359 16890 31383 16892
rect 31439 16890 31463 16892
rect 31519 16890 31525 16892
rect 31279 16838 31281 16890
rect 31461 16838 31463 16890
rect 31217 16836 31223 16838
rect 31279 16836 31303 16838
rect 31359 16836 31383 16838
rect 31439 16836 31463 16838
rect 31519 16836 31525 16838
rect 31217 16827 31525 16836
rect 27365 16348 27673 16357
rect 27365 16346 27371 16348
rect 27427 16346 27451 16348
rect 27507 16346 27531 16348
rect 27587 16346 27611 16348
rect 27667 16346 27673 16348
rect 27427 16294 27429 16346
rect 27609 16294 27611 16346
rect 27365 16292 27371 16294
rect 27427 16292 27451 16294
rect 27507 16292 27531 16294
rect 27587 16292 27611 16294
rect 27667 16292 27673 16294
rect 27365 16283 27673 16292
rect 23512 15804 23820 15813
rect 23512 15802 23518 15804
rect 23574 15802 23598 15804
rect 23654 15802 23678 15804
rect 23734 15802 23758 15804
rect 23814 15802 23820 15804
rect 23574 15750 23576 15802
rect 23756 15750 23758 15802
rect 23512 15748 23518 15750
rect 23574 15748 23598 15750
rect 23654 15748 23678 15750
rect 23734 15748 23758 15750
rect 23814 15748 23820 15750
rect 23512 15739 23820 15748
rect 31217 15804 31525 15813
rect 31217 15802 31223 15804
rect 31279 15802 31303 15804
rect 31359 15802 31383 15804
rect 31439 15802 31463 15804
rect 31519 15802 31525 15804
rect 31279 15750 31281 15802
rect 31461 15750 31463 15802
rect 31217 15748 31223 15750
rect 31279 15748 31303 15750
rect 31359 15748 31383 15750
rect 31439 15748 31463 15750
rect 31519 15748 31525 15750
rect 31217 15739 31525 15748
rect 27365 15260 27673 15269
rect 27365 15258 27371 15260
rect 27427 15258 27451 15260
rect 27507 15258 27531 15260
rect 27587 15258 27611 15260
rect 27667 15258 27673 15260
rect 27427 15206 27429 15258
rect 27609 15206 27611 15258
rect 27365 15204 27371 15206
rect 27427 15204 27451 15206
rect 27507 15204 27531 15206
rect 27587 15204 27611 15206
rect 27667 15204 27673 15206
rect 27365 15195 27673 15204
rect 23512 14716 23820 14725
rect 23512 14714 23518 14716
rect 23574 14714 23598 14716
rect 23654 14714 23678 14716
rect 23734 14714 23758 14716
rect 23814 14714 23820 14716
rect 23574 14662 23576 14714
rect 23756 14662 23758 14714
rect 23512 14660 23518 14662
rect 23574 14660 23598 14662
rect 23654 14660 23678 14662
rect 23734 14660 23758 14662
rect 23814 14660 23820 14662
rect 23512 14651 23820 14660
rect 31217 14716 31525 14725
rect 31217 14714 31223 14716
rect 31279 14714 31303 14716
rect 31359 14714 31383 14716
rect 31439 14714 31463 14716
rect 31519 14714 31525 14716
rect 31279 14662 31281 14714
rect 31461 14662 31463 14714
rect 31217 14660 31223 14662
rect 31279 14660 31303 14662
rect 31359 14660 31383 14662
rect 31439 14660 31463 14662
rect 31519 14660 31525 14662
rect 31217 14651 31525 14660
rect 27365 14172 27673 14181
rect 27365 14170 27371 14172
rect 27427 14170 27451 14172
rect 27507 14170 27531 14172
rect 27587 14170 27611 14172
rect 27667 14170 27673 14172
rect 27427 14118 27429 14170
rect 27609 14118 27611 14170
rect 27365 14116 27371 14118
rect 27427 14116 27451 14118
rect 27507 14116 27531 14118
rect 27587 14116 27611 14118
rect 27667 14116 27673 14118
rect 27365 14107 27673 14116
rect 23512 13628 23820 13637
rect 23512 13626 23518 13628
rect 23574 13626 23598 13628
rect 23654 13626 23678 13628
rect 23734 13626 23758 13628
rect 23814 13626 23820 13628
rect 23574 13574 23576 13626
rect 23756 13574 23758 13626
rect 23512 13572 23518 13574
rect 23574 13572 23598 13574
rect 23654 13572 23678 13574
rect 23734 13572 23758 13574
rect 23814 13572 23820 13574
rect 23512 13563 23820 13572
rect 31217 13628 31525 13637
rect 31217 13626 31223 13628
rect 31279 13626 31303 13628
rect 31359 13626 31383 13628
rect 31439 13626 31463 13628
rect 31519 13626 31525 13628
rect 31279 13574 31281 13626
rect 31461 13574 31463 13626
rect 31217 13572 31223 13574
rect 31279 13572 31303 13574
rect 31359 13572 31383 13574
rect 31439 13572 31463 13574
rect 31519 13572 31525 13574
rect 31217 13563 31525 13572
rect 27365 13084 27673 13093
rect 27365 13082 27371 13084
rect 27427 13082 27451 13084
rect 27507 13082 27531 13084
rect 27587 13082 27611 13084
rect 27667 13082 27673 13084
rect 27427 13030 27429 13082
rect 27609 13030 27611 13082
rect 27365 13028 27371 13030
rect 27427 13028 27451 13030
rect 27507 13028 27531 13030
rect 27587 13028 27611 13030
rect 27667 13028 27673 13030
rect 27365 13019 27673 13028
rect 23512 12540 23820 12549
rect 23512 12538 23518 12540
rect 23574 12538 23598 12540
rect 23654 12538 23678 12540
rect 23734 12538 23758 12540
rect 23814 12538 23820 12540
rect 23574 12486 23576 12538
rect 23756 12486 23758 12538
rect 23512 12484 23518 12486
rect 23574 12484 23598 12486
rect 23654 12484 23678 12486
rect 23734 12484 23758 12486
rect 23814 12484 23820 12486
rect 23512 12475 23820 12484
rect 31217 12540 31525 12549
rect 31217 12538 31223 12540
rect 31279 12538 31303 12540
rect 31359 12538 31383 12540
rect 31439 12538 31463 12540
rect 31519 12538 31525 12540
rect 31279 12486 31281 12538
rect 31461 12486 31463 12538
rect 31217 12484 31223 12486
rect 31279 12484 31303 12486
rect 31359 12484 31383 12486
rect 31439 12484 31463 12486
rect 31519 12484 31525 12486
rect 31217 12475 31525 12484
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20088 11898 20116 12242
rect 27365 11996 27673 12005
rect 27365 11994 27371 11996
rect 27427 11994 27451 11996
rect 27507 11994 27531 11996
rect 27587 11994 27611 11996
rect 27667 11994 27673 11996
rect 27427 11942 27429 11994
rect 27609 11942 27611 11994
rect 27365 11940 27371 11942
rect 27427 11940 27451 11942
rect 27507 11940 27531 11942
rect 27587 11940 27611 11942
rect 27667 11940 27673 11942
rect 27365 11931 27673 11940
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 23512 11452 23820 11461
rect 23512 11450 23518 11452
rect 23574 11450 23598 11452
rect 23654 11450 23678 11452
rect 23734 11450 23758 11452
rect 23814 11450 23820 11452
rect 23574 11398 23576 11450
rect 23756 11398 23758 11450
rect 23512 11396 23518 11398
rect 23574 11396 23598 11398
rect 23654 11396 23678 11398
rect 23734 11396 23758 11398
rect 23814 11396 23820 11398
rect 23512 11387 23820 11396
rect 31217 11452 31525 11461
rect 31217 11450 31223 11452
rect 31279 11450 31303 11452
rect 31359 11450 31383 11452
rect 31439 11450 31463 11452
rect 31519 11450 31525 11452
rect 31279 11398 31281 11450
rect 31461 11398 31463 11450
rect 31217 11396 31223 11398
rect 31279 11396 31303 11398
rect 31359 11396 31383 11398
rect 31439 11396 31463 11398
rect 31519 11396 31525 11398
rect 31217 11387 31525 11396
rect 20076 11348 20128 11354
rect 19996 11308 20076 11336
rect 20076 11290 20128 11296
rect 19660 10908 19968 10917
rect 19660 10906 19666 10908
rect 19722 10906 19746 10908
rect 19802 10906 19826 10908
rect 19882 10906 19906 10908
rect 19962 10906 19968 10908
rect 19722 10854 19724 10906
rect 19904 10854 19906 10906
rect 19660 10852 19666 10854
rect 19722 10852 19746 10854
rect 19802 10852 19826 10854
rect 19882 10852 19906 10854
rect 19962 10852 19968 10854
rect 19660 10843 19968 10852
rect 27365 10908 27673 10917
rect 27365 10906 27371 10908
rect 27427 10906 27451 10908
rect 27507 10906 27531 10908
rect 27587 10906 27611 10908
rect 27667 10906 27673 10908
rect 27427 10854 27429 10906
rect 27609 10854 27611 10906
rect 27365 10852 27371 10854
rect 27427 10852 27451 10854
rect 27507 10852 27531 10854
rect 27587 10852 27611 10854
rect 27667 10852 27673 10854
rect 27365 10843 27673 10852
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 19076 9654 19104 10474
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 18512 9648 18564 9654
rect 18340 9042 18368 9646
rect 18512 9590 18564 9596
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18340 8498 18368 8978
rect 18984 8634 19012 9318
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7546 18276 7686
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 19076 7478 19104 9590
rect 19444 9110 19472 9862
rect 19536 9722 19564 10406
rect 19628 10266 19656 10406
rect 20180 10266 20208 10406
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 19660 9820 19968 9829
rect 19660 9818 19666 9820
rect 19722 9818 19746 9820
rect 19802 9818 19826 9820
rect 19882 9818 19906 9820
rect 19962 9818 19968 9820
rect 19722 9766 19724 9818
rect 19904 9766 19906 9818
rect 19660 9764 19666 9766
rect 19722 9764 19746 9766
rect 19802 9764 19826 9766
rect 19882 9764 19906 9766
rect 19962 9764 19968 9766
rect 19660 9755 19968 9764
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 20548 9518 20576 10542
rect 23512 10364 23820 10373
rect 23512 10362 23518 10364
rect 23574 10362 23598 10364
rect 23654 10362 23678 10364
rect 23734 10362 23758 10364
rect 23814 10362 23820 10364
rect 23574 10310 23576 10362
rect 23756 10310 23758 10362
rect 23512 10308 23518 10310
rect 23574 10308 23598 10310
rect 23654 10308 23678 10310
rect 23734 10308 23758 10310
rect 23814 10308 23820 10310
rect 23512 10299 23820 10308
rect 31217 10364 31525 10373
rect 31217 10362 31223 10364
rect 31279 10362 31303 10364
rect 31359 10362 31383 10364
rect 31439 10362 31463 10364
rect 31519 10362 31525 10364
rect 31279 10310 31281 10362
rect 31461 10310 31463 10362
rect 31217 10308 31223 10310
rect 31279 10308 31303 10310
rect 31359 10308 31383 10310
rect 31439 10308 31463 10310
rect 31519 10308 31525 10310
rect 31217 10299 31525 10308
rect 31666 10296 31722 10305
rect 31666 10231 31722 10240
rect 31680 10198 31708 10231
rect 31668 10192 31720 10198
rect 31668 10134 31720 10140
rect 27365 9820 27673 9829
rect 27365 9818 27371 9820
rect 27427 9818 27451 9820
rect 27507 9818 27531 9820
rect 27587 9818 27611 9820
rect 27667 9818 27673 9820
rect 27427 9766 27429 9818
rect 27609 9766 27611 9818
rect 27365 9764 27371 9766
rect 27427 9764 27451 9766
rect 27507 9764 27531 9766
rect 27587 9764 27611 9766
rect 27667 9764 27673 9766
rect 27365 9755 27673 9764
rect 28262 9616 28318 9625
rect 28262 9551 28318 9560
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 20548 9042 20576 9454
rect 23512 9276 23820 9285
rect 23512 9274 23518 9276
rect 23574 9274 23598 9276
rect 23654 9274 23678 9276
rect 23734 9274 23758 9276
rect 23814 9274 23820 9276
rect 23574 9222 23576 9274
rect 23756 9222 23758 9274
rect 23512 9220 23518 9222
rect 23574 9220 23598 9222
rect 23654 9220 23678 9222
rect 23734 9220 23758 9222
rect 23814 9220 23820 9222
rect 23512 9211 23820 9220
rect 28276 9178 28304 9551
rect 31217 9276 31525 9285
rect 31217 9274 31223 9276
rect 31279 9274 31303 9276
rect 31359 9274 31383 9276
rect 31439 9274 31463 9276
rect 31519 9274 31525 9276
rect 31279 9222 31281 9274
rect 31461 9222 31463 9274
rect 31217 9220 31223 9222
rect 31279 9220 31303 9222
rect 31359 9220 31383 9222
rect 31439 9220 31463 9222
rect 31519 9220 31525 9222
rect 31217 9211 31525 9220
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 7546 19380 8230
rect 19444 7546 19472 8298
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 6934 17540 7142
rect 18156 6934 18184 7210
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18064 6644 18092 6802
rect 18328 6656 18380 6662
rect 18064 6616 18328 6644
rect 18328 6598 18380 6604
rect 18892 2774 18920 7142
rect 19444 7002 19472 7278
rect 19536 7002 19564 8978
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19660 8732 19968 8741
rect 19660 8730 19666 8732
rect 19722 8730 19746 8732
rect 19802 8730 19826 8732
rect 19882 8730 19906 8732
rect 19962 8730 19968 8732
rect 19722 8678 19724 8730
rect 19904 8678 19906 8730
rect 19660 8676 19666 8678
rect 19722 8676 19746 8678
rect 19802 8676 19826 8678
rect 19882 8676 19906 8678
rect 19962 8676 19968 8678
rect 19660 8667 19968 8676
rect 19996 8498 20024 8774
rect 20364 8634 20392 8978
rect 20444 8968 20496 8974
rect 20916 8922 20944 8978
rect 20444 8910 20496 8916
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19660 7644 19968 7653
rect 19660 7642 19666 7644
rect 19722 7642 19746 7644
rect 19802 7642 19826 7644
rect 19882 7642 19906 7644
rect 19962 7642 19968 7644
rect 19722 7590 19724 7642
rect 19904 7590 19906 7642
rect 19660 7588 19666 7590
rect 19722 7588 19746 7590
rect 19802 7588 19826 7590
rect 19882 7588 19906 7590
rect 19962 7588 19968 7590
rect 19660 7579 19968 7588
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19660 6556 19968 6565
rect 19660 6554 19666 6556
rect 19722 6554 19746 6556
rect 19802 6554 19826 6556
rect 19882 6554 19906 6556
rect 19962 6554 19968 6556
rect 19722 6502 19724 6554
rect 19904 6502 19906 6554
rect 19660 6500 19666 6502
rect 19722 6500 19746 6502
rect 19802 6500 19826 6502
rect 19882 6500 19906 6502
rect 19962 6500 19968 6502
rect 19660 6491 19968 6500
rect 19660 5468 19968 5477
rect 19660 5466 19666 5468
rect 19722 5466 19746 5468
rect 19802 5466 19826 5468
rect 19882 5466 19906 5468
rect 19962 5466 19968 5468
rect 19722 5414 19724 5466
rect 19904 5414 19906 5466
rect 19660 5412 19666 5414
rect 19722 5412 19746 5414
rect 19802 5412 19826 5414
rect 19882 5412 19906 5414
rect 19962 5412 19968 5414
rect 19660 5403 19968 5412
rect 19660 4380 19968 4389
rect 19660 4378 19666 4380
rect 19722 4378 19746 4380
rect 19802 4378 19826 4380
rect 19882 4378 19906 4380
rect 19962 4378 19968 4380
rect 19722 4326 19724 4378
rect 19904 4326 19906 4378
rect 19660 4324 19666 4326
rect 19722 4324 19746 4326
rect 19802 4324 19826 4326
rect 19882 4324 19906 4326
rect 19962 4324 19968 4326
rect 19660 4315 19968 4324
rect 19660 3292 19968 3301
rect 19660 3290 19666 3292
rect 19722 3290 19746 3292
rect 19802 3290 19826 3292
rect 19882 3290 19906 3292
rect 19962 3290 19968 3292
rect 19722 3238 19724 3290
rect 19904 3238 19906 3290
rect 19660 3236 19666 3238
rect 19722 3236 19746 3238
rect 19802 3236 19826 3238
rect 19882 3236 19906 3238
rect 19962 3236 19968 3238
rect 19660 3227 19968 3236
rect 18708 2746 18920 2774
rect 18708 400 18736 2746
rect 19660 2204 19968 2213
rect 19660 2202 19666 2204
rect 19722 2202 19746 2204
rect 19802 2202 19826 2204
rect 19882 2202 19906 2204
rect 19962 2202 19968 2204
rect 19722 2150 19724 2202
rect 19904 2150 19906 2202
rect 19660 2148 19666 2150
rect 19722 2148 19746 2150
rect 19802 2148 19826 2150
rect 19882 2148 19906 2150
rect 19962 2148 19968 2150
rect 19660 2139 19968 2148
rect 19660 1116 19968 1125
rect 19660 1114 19666 1116
rect 19722 1114 19746 1116
rect 19802 1114 19826 1116
rect 19882 1114 19906 1116
rect 19962 1114 19968 1116
rect 19722 1062 19724 1114
rect 19904 1062 19906 1114
rect 19660 1060 19666 1062
rect 19722 1060 19746 1062
rect 19802 1060 19826 1062
rect 19882 1060 19906 1062
rect 19962 1060 19968 1062
rect 19660 1051 19968 1060
rect 19996 400 20024 7686
rect 20272 6866 20300 8298
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20364 7546 20392 7890
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20456 6798 20484 8910
rect 20640 8894 20944 8922
rect 28262 8936 28318 8945
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20548 6798 20576 8774
rect 20640 7410 20668 8894
rect 28262 8871 28264 8880
rect 28316 8871 28318 8880
rect 28264 8842 28316 8848
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20824 7818 20852 8230
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 21376 6866 21404 8774
rect 27365 8732 27673 8741
rect 27365 8730 27371 8732
rect 27427 8730 27451 8732
rect 27507 8730 27531 8732
rect 27587 8730 27611 8732
rect 27667 8730 27673 8732
rect 27427 8678 27429 8730
rect 27609 8678 27611 8730
rect 27365 8676 27371 8678
rect 27427 8676 27451 8678
rect 27507 8676 27531 8678
rect 27587 8676 27611 8678
rect 27667 8676 27673 8678
rect 27365 8667 27673 8676
rect 23512 8188 23820 8197
rect 23512 8186 23518 8188
rect 23574 8186 23598 8188
rect 23654 8186 23678 8188
rect 23734 8186 23758 8188
rect 23814 8186 23820 8188
rect 23574 8134 23576 8186
rect 23756 8134 23758 8186
rect 23512 8132 23518 8134
rect 23574 8132 23598 8134
rect 23654 8132 23678 8134
rect 23734 8132 23758 8134
rect 23814 8132 23820 8134
rect 23512 8123 23820 8132
rect 31217 8188 31525 8197
rect 31217 8186 31223 8188
rect 31279 8186 31303 8188
rect 31359 8186 31383 8188
rect 31439 8186 31463 8188
rect 31519 8186 31525 8188
rect 31279 8134 31281 8186
rect 31461 8134 31463 8186
rect 31217 8132 31223 8134
rect 31279 8132 31303 8134
rect 31359 8132 31383 8134
rect 31439 8132 31463 8134
rect 31519 8132 31525 8134
rect 31217 8123 31525 8132
rect 27365 7644 27673 7653
rect 27365 7642 27371 7644
rect 27427 7642 27451 7644
rect 27507 7642 27531 7644
rect 27587 7642 27611 7644
rect 27667 7642 27673 7644
rect 27427 7590 27429 7642
rect 27609 7590 27611 7642
rect 27365 7588 27371 7590
rect 27427 7588 27451 7590
rect 27507 7588 27531 7590
rect 27587 7588 27611 7590
rect 27667 7588 27673 7590
rect 27365 7579 27673 7588
rect 23512 7100 23820 7109
rect 23512 7098 23518 7100
rect 23574 7098 23598 7100
rect 23654 7098 23678 7100
rect 23734 7098 23758 7100
rect 23814 7098 23820 7100
rect 23574 7046 23576 7098
rect 23756 7046 23758 7098
rect 23512 7044 23518 7046
rect 23574 7044 23598 7046
rect 23654 7044 23678 7046
rect 23734 7044 23758 7046
rect 23814 7044 23820 7046
rect 23512 7035 23820 7044
rect 31217 7100 31525 7109
rect 31217 7098 31223 7100
rect 31279 7098 31303 7100
rect 31359 7098 31383 7100
rect 31439 7098 31463 7100
rect 31519 7098 31525 7100
rect 31279 7046 31281 7098
rect 31461 7046 31463 7098
rect 31217 7044 31223 7046
rect 31279 7044 31303 7046
rect 31359 7044 31383 7046
rect 31439 7044 31463 7046
rect 31519 7044 31525 7046
rect 31217 7035 31525 7044
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 27365 6556 27673 6565
rect 27365 6554 27371 6556
rect 27427 6554 27451 6556
rect 27507 6554 27531 6556
rect 27587 6554 27611 6556
rect 27667 6554 27673 6556
rect 27427 6502 27429 6554
rect 27609 6502 27611 6554
rect 27365 6500 27371 6502
rect 27427 6500 27451 6502
rect 27507 6500 27531 6502
rect 27587 6500 27611 6502
rect 27667 6500 27673 6502
rect 27365 6491 27673 6500
rect 23512 6012 23820 6021
rect 23512 6010 23518 6012
rect 23574 6010 23598 6012
rect 23654 6010 23678 6012
rect 23734 6010 23758 6012
rect 23814 6010 23820 6012
rect 23574 5958 23576 6010
rect 23756 5958 23758 6010
rect 23512 5956 23518 5958
rect 23574 5956 23598 5958
rect 23654 5956 23678 5958
rect 23734 5956 23758 5958
rect 23814 5956 23820 5958
rect 23512 5947 23820 5956
rect 31217 6012 31525 6021
rect 31217 6010 31223 6012
rect 31279 6010 31303 6012
rect 31359 6010 31383 6012
rect 31439 6010 31463 6012
rect 31519 6010 31525 6012
rect 31279 5958 31281 6010
rect 31461 5958 31463 6010
rect 31217 5956 31223 5958
rect 31279 5956 31303 5958
rect 31359 5956 31383 5958
rect 31439 5956 31463 5958
rect 31519 5956 31525 5958
rect 31217 5947 31525 5956
rect 27365 5468 27673 5477
rect 27365 5466 27371 5468
rect 27427 5466 27451 5468
rect 27507 5466 27531 5468
rect 27587 5466 27611 5468
rect 27667 5466 27673 5468
rect 27427 5414 27429 5466
rect 27609 5414 27611 5466
rect 27365 5412 27371 5414
rect 27427 5412 27451 5414
rect 27507 5412 27531 5414
rect 27587 5412 27611 5414
rect 27667 5412 27673 5414
rect 27365 5403 27673 5412
rect 23512 4924 23820 4933
rect 23512 4922 23518 4924
rect 23574 4922 23598 4924
rect 23654 4922 23678 4924
rect 23734 4922 23758 4924
rect 23814 4922 23820 4924
rect 23574 4870 23576 4922
rect 23756 4870 23758 4922
rect 23512 4868 23518 4870
rect 23574 4868 23598 4870
rect 23654 4868 23678 4870
rect 23734 4868 23758 4870
rect 23814 4868 23820 4870
rect 23512 4859 23820 4868
rect 31217 4924 31525 4933
rect 31217 4922 31223 4924
rect 31279 4922 31303 4924
rect 31359 4922 31383 4924
rect 31439 4922 31463 4924
rect 31519 4922 31525 4924
rect 31279 4870 31281 4922
rect 31461 4870 31463 4922
rect 31217 4868 31223 4870
rect 31279 4868 31303 4870
rect 31359 4868 31383 4870
rect 31439 4868 31463 4870
rect 31519 4868 31525 4870
rect 31217 4859 31525 4868
rect 27365 4380 27673 4389
rect 27365 4378 27371 4380
rect 27427 4378 27451 4380
rect 27507 4378 27531 4380
rect 27587 4378 27611 4380
rect 27667 4378 27673 4380
rect 27427 4326 27429 4378
rect 27609 4326 27611 4378
rect 27365 4324 27371 4326
rect 27427 4324 27451 4326
rect 27507 4324 27531 4326
rect 27587 4324 27611 4326
rect 27667 4324 27673 4326
rect 27365 4315 27673 4324
rect 23512 3836 23820 3845
rect 23512 3834 23518 3836
rect 23574 3834 23598 3836
rect 23654 3834 23678 3836
rect 23734 3834 23758 3836
rect 23814 3834 23820 3836
rect 23574 3782 23576 3834
rect 23756 3782 23758 3834
rect 23512 3780 23518 3782
rect 23574 3780 23598 3782
rect 23654 3780 23678 3782
rect 23734 3780 23758 3782
rect 23814 3780 23820 3782
rect 23512 3771 23820 3780
rect 31217 3836 31525 3845
rect 31217 3834 31223 3836
rect 31279 3834 31303 3836
rect 31359 3834 31383 3836
rect 31439 3834 31463 3836
rect 31519 3834 31525 3836
rect 31279 3782 31281 3834
rect 31461 3782 31463 3834
rect 31217 3780 31223 3782
rect 31279 3780 31303 3782
rect 31359 3780 31383 3782
rect 31439 3780 31463 3782
rect 31519 3780 31525 3782
rect 31217 3771 31525 3780
rect 27365 3292 27673 3301
rect 27365 3290 27371 3292
rect 27427 3290 27451 3292
rect 27507 3290 27531 3292
rect 27587 3290 27611 3292
rect 27667 3290 27673 3292
rect 27427 3238 27429 3290
rect 27609 3238 27611 3290
rect 27365 3236 27371 3238
rect 27427 3236 27451 3238
rect 27507 3236 27531 3238
rect 27587 3236 27611 3238
rect 27667 3236 27673 3238
rect 27365 3227 27673 3236
rect 23512 2748 23820 2757
rect 23512 2746 23518 2748
rect 23574 2746 23598 2748
rect 23654 2746 23678 2748
rect 23734 2746 23758 2748
rect 23814 2746 23820 2748
rect 23574 2694 23576 2746
rect 23756 2694 23758 2746
rect 23512 2692 23518 2694
rect 23574 2692 23598 2694
rect 23654 2692 23678 2694
rect 23734 2692 23758 2694
rect 23814 2692 23820 2694
rect 23512 2683 23820 2692
rect 31217 2748 31525 2757
rect 31217 2746 31223 2748
rect 31279 2746 31303 2748
rect 31359 2746 31383 2748
rect 31439 2746 31463 2748
rect 31519 2746 31525 2748
rect 31279 2694 31281 2746
rect 31461 2694 31463 2746
rect 31217 2692 31223 2694
rect 31279 2692 31303 2694
rect 31359 2692 31383 2694
rect 31439 2692 31463 2694
rect 31519 2692 31525 2694
rect 31217 2683 31525 2692
rect 27365 2204 27673 2213
rect 27365 2202 27371 2204
rect 27427 2202 27451 2204
rect 27507 2202 27531 2204
rect 27587 2202 27611 2204
rect 27667 2202 27673 2204
rect 27427 2150 27429 2202
rect 27609 2150 27611 2202
rect 27365 2148 27371 2150
rect 27427 2148 27451 2150
rect 27507 2148 27531 2150
rect 27587 2148 27611 2150
rect 27667 2148 27673 2150
rect 27365 2139 27673 2148
rect 23512 1660 23820 1669
rect 23512 1658 23518 1660
rect 23574 1658 23598 1660
rect 23654 1658 23678 1660
rect 23734 1658 23758 1660
rect 23814 1658 23820 1660
rect 23574 1606 23576 1658
rect 23756 1606 23758 1658
rect 23512 1604 23518 1606
rect 23574 1604 23598 1606
rect 23654 1604 23678 1606
rect 23734 1604 23758 1606
rect 23814 1604 23820 1606
rect 23512 1595 23820 1604
rect 31217 1660 31525 1669
rect 31217 1658 31223 1660
rect 31279 1658 31303 1660
rect 31359 1658 31383 1660
rect 31439 1658 31463 1660
rect 31519 1658 31525 1660
rect 31279 1606 31281 1658
rect 31461 1606 31463 1658
rect 31217 1604 31223 1606
rect 31279 1604 31303 1606
rect 31359 1604 31383 1606
rect 31439 1604 31463 1606
rect 31519 1604 31525 1606
rect 31217 1595 31525 1604
rect 27365 1116 27673 1125
rect 27365 1114 27371 1116
rect 27427 1114 27451 1116
rect 27507 1114 27531 1116
rect 27587 1114 27611 1116
rect 27667 1114 27673 1116
rect 27427 1062 27429 1114
rect 27609 1062 27611 1114
rect 27365 1060 27371 1062
rect 27427 1060 27451 1062
rect 27507 1060 27531 1062
rect 27587 1060 27611 1062
rect 27667 1060 27673 1062
rect 27365 1051 27673 1060
rect 23512 572 23820 581
rect 23512 570 23518 572
rect 23574 570 23598 572
rect 23654 570 23678 572
rect 23734 570 23758 572
rect 23814 570 23820 572
rect 23574 518 23576 570
rect 23756 518 23758 570
rect 23512 516 23518 518
rect 23574 516 23598 518
rect 23654 516 23678 518
rect 23734 516 23758 518
rect 23814 516 23820 518
rect 23512 507 23820 516
rect 31217 572 31525 581
rect 31217 570 31223 572
rect 31279 570 31303 572
rect 31359 570 31383 572
rect 31439 570 31463 572
rect 31519 570 31525 572
rect 31279 518 31281 570
rect 31461 518 31463 570
rect 31217 516 31223 518
rect 31279 516 31303 518
rect 31359 516 31383 518
rect 31439 516 31463 518
rect 31519 516 31525 518
rect 31217 507 31525 516
rect 16868 326 17080 354
rect 18694 0 18750 400
rect 19982 0 20038 400
<< via2 >>
rect 8108 19066 8164 19068
rect 8188 19066 8244 19068
rect 8268 19066 8324 19068
rect 8348 19066 8404 19068
rect 8108 19014 8154 19066
rect 8154 19014 8164 19066
rect 8188 19014 8218 19066
rect 8218 19014 8230 19066
rect 8230 19014 8244 19066
rect 8268 19014 8282 19066
rect 8282 19014 8294 19066
rect 8294 19014 8324 19066
rect 8348 19014 8358 19066
rect 8358 19014 8404 19066
rect 8108 19012 8164 19014
rect 8188 19012 8244 19014
rect 8268 19012 8324 19014
rect 8348 19012 8404 19014
rect 4256 18522 4312 18524
rect 4336 18522 4392 18524
rect 4416 18522 4472 18524
rect 4496 18522 4552 18524
rect 4256 18470 4302 18522
rect 4302 18470 4312 18522
rect 4336 18470 4366 18522
rect 4366 18470 4378 18522
rect 4378 18470 4392 18522
rect 4416 18470 4430 18522
rect 4430 18470 4442 18522
rect 4442 18470 4472 18522
rect 4496 18470 4506 18522
rect 4506 18470 4552 18522
rect 4256 18468 4312 18470
rect 4336 18468 4392 18470
rect 4416 18468 4472 18470
rect 4496 18468 4552 18470
rect 11961 18522 12017 18524
rect 12041 18522 12097 18524
rect 12121 18522 12177 18524
rect 12201 18522 12257 18524
rect 11961 18470 12007 18522
rect 12007 18470 12017 18522
rect 12041 18470 12071 18522
rect 12071 18470 12083 18522
rect 12083 18470 12097 18522
rect 12121 18470 12135 18522
rect 12135 18470 12147 18522
rect 12147 18470 12177 18522
rect 12201 18470 12211 18522
rect 12211 18470 12257 18522
rect 11961 18468 12017 18470
rect 12041 18468 12097 18470
rect 12121 18468 12177 18470
rect 12201 18468 12257 18470
rect 8108 17978 8164 17980
rect 8188 17978 8244 17980
rect 8268 17978 8324 17980
rect 8348 17978 8404 17980
rect 8108 17926 8154 17978
rect 8154 17926 8164 17978
rect 8188 17926 8218 17978
rect 8218 17926 8230 17978
rect 8230 17926 8244 17978
rect 8268 17926 8282 17978
rect 8282 17926 8294 17978
rect 8294 17926 8324 17978
rect 8348 17926 8358 17978
rect 8358 17926 8404 17978
rect 8108 17924 8164 17926
rect 8188 17924 8244 17926
rect 8268 17924 8324 17926
rect 8348 17924 8404 17926
rect 4256 17434 4312 17436
rect 4336 17434 4392 17436
rect 4416 17434 4472 17436
rect 4496 17434 4552 17436
rect 4256 17382 4302 17434
rect 4302 17382 4312 17434
rect 4336 17382 4366 17434
rect 4366 17382 4378 17434
rect 4378 17382 4392 17434
rect 4416 17382 4430 17434
rect 4430 17382 4442 17434
rect 4442 17382 4472 17434
rect 4496 17382 4506 17434
rect 4506 17382 4552 17434
rect 4256 17380 4312 17382
rect 4336 17380 4392 17382
rect 4416 17380 4472 17382
rect 4496 17380 4552 17382
rect 11961 17434 12017 17436
rect 12041 17434 12097 17436
rect 12121 17434 12177 17436
rect 12201 17434 12257 17436
rect 11961 17382 12007 17434
rect 12007 17382 12017 17434
rect 12041 17382 12071 17434
rect 12071 17382 12083 17434
rect 12083 17382 12097 17434
rect 12121 17382 12135 17434
rect 12135 17382 12147 17434
rect 12147 17382 12177 17434
rect 12201 17382 12211 17434
rect 12211 17382 12257 17434
rect 11961 17380 12017 17382
rect 12041 17380 12097 17382
rect 12121 17380 12177 17382
rect 12201 17380 12257 17382
rect 8108 16890 8164 16892
rect 8188 16890 8244 16892
rect 8268 16890 8324 16892
rect 8348 16890 8404 16892
rect 8108 16838 8154 16890
rect 8154 16838 8164 16890
rect 8188 16838 8218 16890
rect 8218 16838 8230 16890
rect 8230 16838 8244 16890
rect 8268 16838 8282 16890
rect 8282 16838 8294 16890
rect 8294 16838 8324 16890
rect 8348 16838 8358 16890
rect 8358 16838 8404 16890
rect 8108 16836 8164 16838
rect 8188 16836 8244 16838
rect 8268 16836 8324 16838
rect 8348 16836 8404 16838
rect 15813 19066 15869 19068
rect 15893 19066 15949 19068
rect 15973 19066 16029 19068
rect 16053 19066 16109 19068
rect 15813 19014 15859 19066
rect 15859 19014 15869 19066
rect 15893 19014 15923 19066
rect 15923 19014 15935 19066
rect 15935 19014 15949 19066
rect 15973 19014 15987 19066
rect 15987 19014 15999 19066
rect 15999 19014 16029 19066
rect 16053 19014 16063 19066
rect 16063 19014 16109 19066
rect 15813 19012 15869 19014
rect 15893 19012 15949 19014
rect 15973 19012 16029 19014
rect 16053 19012 16109 19014
rect 4256 16346 4312 16348
rect 4336 16346 4392 16348
rect 4416 16346 4472 16348
rect 4496 16346 4552 16348
rect 4256 16294 4302 16346
rect 4302 16294 4312 16346
rect 4336 16294 4366 16346
rect 4366 16294 4378 16346
rect 4378 16294 4392 16346
rect 4416 16294 4430 16346
rect 4430 16294 4442 16346
rect 4442 16294 4472 16346
rect 4496 16294 4506 16346
rect 4506 16294 4552 16346
rect 4256 16292 4312 16294
rect 4336 16292 4392 16294
rect 4416 16292 4472 16294
rect 4496 16292 4552 16294
rect 11961 16346 12017 16348
rect 12041 16346 12097 16348
rect 12121 16346 12177 16348
rect 12201 16346 12257 16348
rect 11961 16294 12007 16346
rect 12007 16294 12017 16346
rect 12041 16294 12071 16346
rect 12071 16294 12083 16346
rect 12083 16294 12097 16346
rect 12121 16294 12135 16346
rect 12135 16294 12147 16346
rect 12147 16294 12177 16346
rect 12201 16294 12211 16346
rect 12211 16294 12257 16346
rect 11961 16292 12017 16294
rect 12041 16292 12097 16294
rect 12121 16292 12177 16294
rect 12201 16292 12257 16294
rect 8108 15802 8164 15804
rect 8188 15802 8244 15804
rect 8268 15802 8324 15804
rect 8348 15802 8404 15804
rect 8108 15750 8154 15802
rect 8154 15750 8164 15802
rect 8188 15750 8218 15802
rect 8218 15750 8230 15802
rect 8230 15750 8244 15802
rect 8268 15750 8282 15802
rect 8282 15750 8294 15802
rect 8294 15750 8324 15802
rect 8348 15750 8358 15802
rect 8358 15750 8404 15802
rect 8108 15748 8164 15750
rect 8188 15748 8244 15750
rect 8268 15748 8324 15750
rect 8348 15748 8404 15750
rect 4256 15258 4312 15260
rect 4336 15258 4392 15260
rect 4416 15258 4472 15260
rect 4496 15258 4552 15260
rect 4256 15206 4302 15258
rect 4302 15206 4312 15258
rect 4336 15206 4366 15258
rect 4366 15206 4378 15258
rect 4378 15206 4392 15258
rect 4416 15206 4430 15258
rect 4430 15206 4442 15258
rect 4442 15206 4472 15258
rect 4496 15206 4506 15258
rect 4506 15206 4552 15258
rect 4256 15204 4312 15206
rect 4336 15204 4392 15206
rect 4416 15204 4472 15206
rect 4496 15204 4552 15206
rect 11961 15258 12017 15260
rect 12041 15258 12097 15260
rect 12121 15258 12177 15260
rect 12201 15258 12257 15260
rect 11961 15206 12007 15258
rect 12007 15206 12017 15258
rect 12041 15206 12071 15258
rect 12071 15206 12083 15258
rect 12083 15206 12097 15258
rect 12121 15206 12135 15258
rect 12135 15206 12147 15258
rect 12147 15206 12177 15258
rect 12201 15206 12211 15258
rect 12211 15206 12257 15258
rect 11961 15204 12017 15206
rect 12041 15204 12097 15206
rect 12121 15204 12177 15206
rect 12201 15204 12257 15206
rect 8108 14714 8164 14716
rect 8188 14714 8244 14716
rect 8268 14714 8324 14716
rect 8348 14714 8404 14716
rect 8108 14662 8154 14714
rect 8154 14662 8164 14714
rect 8188 14662 8218 14714
rect 8218 14662 8230 14714
rect 8230 14662 8244 14714
rect 8268 14662 8282 14714
rect 8282 14662 8294 14714
rect 8294 14662 8324 14714
rect 8348 14662 8358 14714
rect 8358 14662 8404 14714
rect 8108 14660 8164 14662
rect 8188 14660 8244 14662
rect 8268 14660 8324 14662
rect 8348 14660 8404 14662
rect 4256 14170 4312 14172
rect 4336 14170 4392 14172
rect 4416 14170 4472 14172
rect 4496 14170 4552 14172
rect 4256 14118 4302 14170
rect 4302 14118 4312 14170
rect 4336 14118 4366 14170
rect 4366 14118 4378 14170
rect 4378 14118 4392 14170
rect 4416 14118 4430 14170
rect 4430 14118 4442 14170
rect 4442 14118 4472 14170
rect 4496 14118 4506 14170
rect 4506 14118 4552 14170
rect 4256 14116 4312 14118
rect 4336 14116 4392 14118
rect 4416 14116 4472 14118
rect 4496 14116 4552 14118
rect 11961 14170 12017 14172
rect 12041 14170 12097 14172
rect 12121 14170 12177 14172
rect 12201 14170 12257 14172
rect 11961 14118 12007 14170
rect 12007 14118 12017 14170
rect 12041 14118 12071 14170
rect 12071 14118 12083 14170
rect 12083 14118 12097 14170
rect 12121 14118 12135 14170
rect 12135 14118 12147 14170
rect 12147 14118 12177 14170
rect 12201 14118 12211 14170
rect 12211 14118 12257 14170
rect 11961 14116 12017 14118
rect 12041 14116 12097 14118
rect 12121 14116 12177 14118
rect 12201 14116 12257 14118
rect 8108 13626 8164 13628
rect 8188 13626 8244 13628
rect 8268 13626 8324 13628
rect 8348 13626 8404 13628
rect 8108 13574 8154 13626
rect 8154 13574 8164 13626
rect 8188 13574 8218 13626
rect 8218 13574 8230 13626
rect 8230 13574 8244 13626
rect 8268 13574 8282 13626
rect 8282 13574 8294 13626
rect 8294 13574 8324 13626
rect 8348 13574 8358 13626
rect 8358 13574 8404 13626
rect 8108 13572 8164 13574
rect 8188 13572 8244 13574
rect 8268 13572 8324 13574
rect 8348 13572 8404 13574
rect 4256 13082 4312 13084
rect 4336 13082 4392 13084
rect 4416 13082 4472 13084
rect 4496 13082 4552 13084
rect 4256 13030 4302 13082
rect 4302 13030 4312 13082
rect 4336 13030 4366 13082
rect 4366 13030 4378 13082
rect 4378 13030 4392 13082
rect 4416 13030 4430 13082
rect 4430 13030 4442 13082
rect 4442 13030 4472 13082
rect 4496 13030 4506 13082
rect 4506 13030 4552 13082
rect 4256 13028 4312 13030
rect 4336 13028 4392 13030
rect 4416 13028 4472 13030
rect 4496 13028 4552 13030
rect 11961 13082 12017 13084
rect 12041 13082 12097 13084
rect 12121 13082 12177 13084
rect 12201 13082 12257 13084
rect 11961 13030 12007 13082
rect 12007 13030 12017 13082
rect 12041 13030 12071 13082
rect 12071 13030 12083 13082
rect 12083 13030 12097 13082
rect 12121 13030 12135 13082
rect 12135 13030 12147 13082
rect 12147 13030 12177 13082
rect 12201 13030 12211 13082
rect 12211 13030 12257 13082
rect 11961 13028 12017 13030
rect 12041 13028 12097 13030
rect 12121 13028 12177 13030
rect 12201 13028 12257 13030
rect 8108 12538 8164 12540
rect 8188 12538 8244 12540
rect 8268 12538 8324 12540
rect 8348 12538 8404 12540
rect 8108 12486 8154 12538
rect 8154 12486 8164 12538
rect 8188 12486 8218 12538
rect 8218 12486 8230 12538
rect 8230 12486 8244 12538
rect 8268 12486 8282 12538
rect 8282 12486 8294 12538
rect 8294 12486 8324 12538
rect 8348 12486 8358 12538
rect 8358 12486 8404 12538
rect 8108 12484 8164 12486
rect 8188 12484 8244 12486
rect 8268 12484 8324 12486
rect 8348 12484 8404 12486
rect 4256 11994 4312 11996
rect 4336 11994 4392 11996
rect 4416 11994 4472 11996
rect 4496 11994 4552 11996
rect 4256 11942 4302 11994
rect 4302 11942 4312 11994
rect 4336 11942 4366 11994
rect 4366 11942 4378 11994
rect 4378 11942 4392 11994
rect 4416 11942 4430 11994
rect 4430 11942 4442 11994
rect 4442 11942 4472 11994
rect 4496 11942 4506 11994
rect 4506 11942 4552 11994
rect 4256 11940 4312 11942
rect 4336 11940 4392 11942
rect 4416 11940 4472 11942
rect 4496 11940 4552 11942
rect 8108 11450 8164 11452
rect 8188 11450 8244 11452
rect 8268 11450 8324 11452
rect 8348 11450 8404 11452
rect 8108 11398 8154 11450
rect 8154 11398 8164 11450
rect 8188 11398 8218 11450
rect 8218 11398 8230 11450
rect 8230 11398 8244 11450
rect 8268 11398 8282 11450
rect 8282 11398 8294 11450
rect 8294 11398 8324 11450
rect 8348 11398 8358 11450
rect 8358 11398 8404 11450
rect 8108 11396 8164 11398
rect 8188 11396 8244 11398
rect 8268 11396 8324 11398
rect 8348 11396 8404 11398
rect 4256 10906 4312 10908
rect 4336 10906 4392 10908
rect 4416 10906 4472 10908
rect 4496 10906 4552 10908
rect 4256 10854 4302 10906
rect 4302 10854 4312 10906
rect 4336 10854 4366 10906
rect 4366 10854 4378 10906
rect 4378 10854 4392 10906
rect 4416 10854 4430 10906
rect 4430 10854 4442 10906
rect 4442 10854 4472 10906
rect 4496 10854 4506 10906
rect 4506 10854 4552 10906
rect 4256 10852 4312 10854
rect 4336 10852 4392 10854
rect 4416 10852 4472 10854
rect 4496 10852 4552 10854
rect 8108 10362 8164 10364
rect 8188 10362 8244 10364
rect 8268 10362 8324 10364
rect 8348 10362 8404 10364
rect 8108 10310 8154 10362
rect 8154 10310 8164 10362
rect 8188 10310 8218 10362
rect 8218 10310 8230 10362
rect 8230 10310 8244 10362
rect 8268 10310 8282 10362
rect 8282 10310 8294 10362
rect 8294 10310 8324 10362
rect 8348 10310 8358 10362
rect 8358 10310 8404 10362
rect 8108 10308 8164 10310
rect 8188 10308 8244 10310
rect 8268 10308 8324 10310
rect 8348 10308 8404 10310
rect 4256 9818 4312 9820
rect 4336 9818 4392 9820
rect 4416 9818 4472 9820
rect 4496 9818 4552 9820
rect 4256 9766 4302 9818
rect 4302 9766 4312 9818
rect 4336 9766 4366 9818
rect 4366 9766 4378 9818
rect 4378 9766 4392 9818
rect 4416 9766 4430 9818
rect 4430 9766 4442 9818
rect 4442 9766 4472 9818
rect 4496 9766 4506 9818
rect 4506 9766 4552 9818
rect 4256 9764 4312 9766
rect 4336 9764 4392 9766
rect 4416 9764 4472 9766
rect 4496 9764 4552 9766
rect 8108 9274 8164 9276
rect 8188 9274 8244 9276
rect 8268 9274 8324 9276
rect 8348 9274 8404 9276
rect 8108 9222 8154 9274
rect 8154 9222 8164 9274
rect 8188 9222 8218 9274
rect 8218 9222 8230 9274
rect 8230 9222 8244 9274
rect 8268 9222 8282 9274
rect 8282 9222 8294 9274
rect 8294 9222 8324 9274
rect 8348 9222 8358 9274
rect 8358 9222 8404 9274
rect 8108 9220 8164 9222
rect 8188 9220 8244 9222
rect 8268 9220 8324 9222
rect 8348 9220 8404 9222
rect 8206 9036 8262 9072
rect 9586 9696 9642 9752
rect 8206 9016 8208 9036
rect 8208 9016 8260 9036
rect 8260 9016 8262 9036
rect 4256 8730 4312 8732
rect 4336 8730 4392 8732
rect 4416 8730 4472 8732
rect 4496 8730 4552 8732
rect 4256 8678 4302 8730
rect 4302 8678 4312 8730
rect 4336 8678 4366 8730
rect 4366 8678 4378 8730
rect 4378 8678 4392 8730
rect 4416 8678 4430 8730
rect 4430 8678 4442 8730
rect 4442 8678 4472 8730
rect 4496 8678 4506 8730
rect 4506 8678 4552 8730
rect 4256 8676 4312 8678
rect 4336 8676 4392 8678
rect 4416 8676 4472 8678
rect 4496 8676 4552 8678
rect 4256 7642 4312 7644
rect 4336 7642 4392 7644
rect 4416 7642 4472 7644
rect 4496 7642 4552 7644
rect 4256 7590 4302 7642
rect 4302 7590 4312 7642
rect 4336 7590 4366 7642
rect 4366 7590 4378 7642
rect 4378 7590 4392 7642
rect 4416 7590 4430 7642
rect 4430 7590 4442 7642
rect 4442 7590 4472 7642
rect 4496 7590 4506 7642
rect 4506 7590 4552 7642
rect 4256 7588 4312 7590
rect 4336 7588 4392 7590
rect 4416 7588 4472 7590
rect 4496 7588 4552 7590
rect 4256 6554 4312 6556
rect 4336 6554 4392 6556
rect 4416 6554 4472 6556
rect 4496 6554 4552 6556
rect 4256 6502 4302 6554
rect 4302 6502 4312 6554
rect 4336 6502 4366 6554
rect 4366 6502 4378 6554
rect 4378 6502 4392 6554
rect 4416 6502 4430 6554
rect 4430 6502 4442 6554
rect 4442 6502 4472 6554
rect 4496 6502 4506 6554
rect 4506 6502 4552 6554
rect 4256 6500 4312 6502
rect 4336 6500 4392 6502
rect 4416 6500 4472 6502
rect 4496 6500 4552 6502
rect 8108 8186 8164 8188
rect 8188 8186 8244 8188
rect 8268 8186 8324 8188
rect 8348 8186 8404 8188
rect 8108 8134 8154 8186
rect 8154 8134 8164 8186
rect 8188 8134 8218 8186
rect 8218 8134 8230 8186
rect 8230 8134 8244 8186
rect 8268 8134 8282 8186
rect 8282 8134 8294 8186
rect 8294 8134 8324 8186
rect 8348 8134 8358 8186
rect 8358 8134 8404 8186
rect 8108 8132 8164 8134
rect 8188 8132 8244 8134
rect 8268 8132 8324 8134
rect 8348 8132 8404 8134
rect 8108 7098 8164 7100
rect 8188 7098 8244 7100
rect 8268 7098 8324 7100
rect 8348 7098 8404 7100
rect 8108 7046 8154 7098
rect 8154 7046 8164 7098
rect 8188 7046 8218 7098
rect 8218 7046 8230 7098
rect 8230 7046 8244 7098
rect 8268 7046 8282 7098
rect 8282 7046 8294 7098
rect 8294 7046 8324 7098
rect 8348 7046 8358 7098
rect 8358 7046 8404 7098
rect 8108 7044 8164 7046
rect 8188 7044 8244 7046
rect 8268 7044 8324 7046
rect 8348 7044 8404 7046
rect 8108 6010 8164 6012
rect 8188 6010 8244 6012
rect 8268 6010 8324 6012
rect 8348 6010 8404 6012
rect 8108 5958 8154 6010
rect 8154 5958 8164 6010
rect 8188 5958 8218 6010
rect 8218 5958 8230 6010
rect 8230 5958 8244 6010
rect 8268 5958 8282 6010
rect 8282 5958 8294 6010
rect 8294 5958 8324 6010
rect 8348 5958 8358 6010
rect 8358 5958 8404 6010
rect 8108 5956 8164 5958
rect 8188 5956 8244 5958
rect 8268 5956 8324 5958
rect 8348 5956 8404 5958
rect 9402 8492 9458 8528
rect 9402 8472 9404 8492
rect 9404 8472 9456 8492
rect 9456 8472 9458 8492
rect 9678 6568 9734 6624
rect 9862 6296 9918 6352
rect 10138 9596 10140 9616
rect 10140 9596 10192 9616
rect 10192 9596 10194 9616
rect 10138 9560 10194 9596
rect 11961 11994 12017 11996
rect 12041 11994 12097 11996
rect 12121 11994 12177 11996
rect 12201 11994 12257 11996
rect 11961 11942 12007 11994
rect 12007 11942 12017 11994
rect 12041 11942 12071 11994
rect 12071 11942 12083 11994
rect 12083 11942 12097 11994
rect 12121 11942 12135 11994
rect 12135 11942 12147 11994
rect 12147 11942 12177 11994
rect 12201 11942 12211 11994
rect 12211 11942 12257 11994
rect 11961 11940 12017 11942
rect 12041 11940 12097 11942
rect 12121 11940 12177 11942
rect 12201 11940 12257 11942
rect 10138 7112 10194 7168
rect 10046 6704 10102 6760
rect 10230 6432 10286 6488
rect 10598 7112 10654 7168
rect 11150 8880 11206 8936
rect 10966 8200 11022 8256
rect 11150 8336 11206 8392
rect 11150 8084 11206 8120
rect 11150 8064 11152 8084
rect 11152 8064 11204 8084
rect 11204 8064 11206 8084
rect 11961 10906 12017 10908
rect 12041 10906 12097 10908
rect 12121 10906 12177 10908
rect 12201 10906 12257 10908
rect 11961 10854 12007 10906
rect 12007 10854 12017 10906
rect 12041 10854 12071 10906
rect 12071 10854 12083 10906
rect 12083 10854 12097 10906
rect 12121 10854 12135 10906
rect 12135 10854 12147 10906
rect 12147 10854 12177 10906
rect 12201 10854 12211 10906
rect 12211 10854 12257 10906
rect 11961 10852 12017 10854
rect 12041 10852 12097 10854
rect 12121 10852 12177 10854
rect 12201 10852 12257 10854
rect 11886 10240 11942 10296
rect 11961 9818 12017 9820
rect 12041 9818 12097 9820
rect 12121 9818 12177 9820
rect 12201 9818 12257 9820
rect 11961 9766 12007 9818
rect 12007 9766 12017 9818
rect 12041 9766 12071 9818
rect 12071 9766 12083 9818
rect 12083 9766 12097 9818
rect 12121 9766 12135 9818
rect 12135 9766 12147 9818
rect 12147 9766 12177 9818
rect 12201 9766 12211 9818
rect 12211 9766 12257 9818
rect 11961 9764 12017 9766
rect 12041 9764 12097 9766
rect 12121 9764 12177 9766
rect 12201 9764 12257 9766
rect 11794 9016 11850 9072
rect 11961 8730 12017 8732
rect 12041 8730 12097 8732
rect 12121 8730 12177 8732
rect 12201 8730 12257 8732
rect 11961 8678 12007 8730
rect 12007 8678 12017 8730
rect 12041 8678 12071 8730
rect 12071 8678 12083 8730
rect 12083 8678 12097 8730
rect 12121 8678 12135 8730
rect 12135 8678 12147 8730
rect 12147 8678 12177 8730
rect 12201 8678 12211 8730
rect 12211 8678 12257 8730
rect 11961 8676 12017 8678
rect 12041 8676 12097 8678
rect 12121 8676 12177 8678
rect 12201 8676 12257 8678
rect 10966 6976 11022 7032
rect 10874 6296 10930 6352
rect 11610 7928 11666 7984
rect 11518 6568 11574 6624
rect 12162 8336 12218 8392
rect 11978 8064 12034 8120
rect 12162 7828 12164 7848
rect 12164 7828 12216 7848
rect 12216 7828 12218 7848
rect 12162 7792 12218 7828
rect 15813 17978 15869 17980
rect 15893 17978 15949 17980
rect 15973 17978 16029 17980
rect 16053 17978 16109 17980
rect 15813 17926 15859 17978
rect 15859 17926 15869 17978
rect 15893 17926 15923 17978
rect 15923 17926 15935 17978
rect 15935 17926 15949 17978
rect 15973 17926 15987 17978
rect 15987 17926 15999 17978
rect 15999 17926 16029 17978
rect 16053 17926 16063 17978
rect 16063 17926 16109 17978
rect 15813 17924 15869 17926
rect 15893 17924 15949 17926
rect 15973 17924 16029 17926
rect 16053 17924 16109 17926
rect 15813 16890 15869 16892
rect 15893 16890 15949 16892
rect 15973 16890 16029 16892
rect 16053 16890 16109 16892
rect 15813 16838 15859 16890
rect 15859 16838 15869 16890
rect 15893 16838 15923 16890
rect 15923 16838 15935 16890
rect 15935 16838 15949 16890
rect 15973 16838 15987 16890
rect 15987 16838 15999 16890
rect 15999 16838 16029 16890
rect 16053 16838 16063 16890
rect 16063 16838 16109 16890
rect 15813 16836 15869 16838
rect 15893 16836 15949 16838
rect 15973 16836 16029 16838
rect 16053 16836 16109 16838
rect 19666 18522 19722 18524
rect 19746 18522 19802 18524
rect 19826 18522 19882 18524
rect 19906 18522 19962 18524
rect 19666 18470 19712 18522
rect 19712 18470 19722 18522
rect 19746 18470 19776 18522
rect 19776 18470 19788 18522
rect 19788 18470 19802 18522
rect 19826 18470 19840 18522
rect 19840 18470 19852 18522
rect 19852 18470 19882 18522
rect 19906 18470 19916 18522
rect 19916 18470 19962 18522
rect 19666 18468 19722 18470
rect 19746 18468 19802 18470
rect 19826 18468 19882 18470
rect 19906 18468 19962 18470
rect 19666 17434 19722 17436
rect 19746 17434 19802 17436
rect 19826 17434 19882 17436
rect 19906 17434 19962 17436
rect 19666 17382 19712 17434
rect 19712 17382 19722 17434
rect 19746 17382 19776 17434
rect 19776 17382 19788 17434
rect 19788 17382 19802 17434
rect 19826 17382 19840 17434
rect 19840 17382 19852 17434
rect 19852 17382 19882 17434
rect 19906 17382 19916 17434
rect 19916 17382 19962 17434
rect 19666 17380 19722 17382
rect 19746 17380 19802 17382
rect 19826 17380 19882 17382
rect 19906 17380 19962 17382
rect 15813 15802 15869 15804
rect 15893 15802 15949 15804
rect 15973 15802 16029 15804
rect 16053 15802 16109 15804
rect 15813 15750 15859 15802
rect 15859 15750 15869 15802
rect 15893 15750 15923 15802
rect 15923 15750 15935 15802
rect 15935 15750 15949 15802
rect 15973 15750 15987 15802
rect 15987 15750 15999 15802
rect 15999 15750 16029 15802
rect 16053 15750 16063 15802
rect 16063 15750 16109 15802
rect 15813 15748 15869 15750
rect 15893 15748 15949 15750
rect 15973 15748 16029 15750
rect 16053 15748 16109 15750
rect 15813 14714 15869 14716
rect 15893 14714 15949 14716
rect 15973 14714 16029 14716
rect 16053 14714 16109 14716
rect 15813 14662 15859 14714
rect 15859 14662 15869 14714
rect 15893 14662 15923 14714
rect 15923 14662 15935 14714
rect 15935 14662 15949 14714
rect 15973 14662 15987 14714
rect 15987 14662 15999 14714
rect 15999 14662 16029 14714
rect 16053 14662 16063 14714
rect 16063 14662 16109 14714
rect 15813 14660 15869 14662
rect 15893 14660 15949 14662
rect 15973 14660 16029 14662
rect 16053 14660 16109 14662
rect 15813 13626 15869 13628
rect 15893 13626 15949 13628
rect 15973 13626 16029 13628
rect 16053 13626 16109 13628
rect 15813 13574 15859 13626
rect 15859 13574 15869 13626
rect 15893 13574 15923 13626
rect 15923 13574 15935 13626
rect 15935 13574 15949 13626
rect 15973 13574 15987 13626
rect 15987 13574 15999 13626
rect 15999 13574 16029 13626
rect 16053 13574 16063 13626
rect 16063 13574 16109 13626
rect 15813 13572 15869 13574
rect 15893 13572 15949 13574
rect 15973 13572 16029 13574
rect 16053 13572 16109 13574
rect 15813 12538 15869 12540
rect 15893 12538 15949 12540
rect 15973 12538 16029 12540
rect 16053 12538 16109 12540
rect 15813 12486 15859 12538
rect 15859 12486 15869 12538
rect 15893 12486 15923 12538
rect 15923 12486 15935 12538
rect 15935 12486 15949 12538
rect 15973 12486 15987 12538
rect 15987 12486 15999 12538
rect 15999 12486 16029 12538
rect 16053 12486 16063 12538
rect 16063 12486 16109 12538
rect 15813 12484 15869 12486
rect 15893 12484 15949 12486
rect 15973 12484 16029 12486
rect 16053 12484 16109 12486
rect 11961 7642 12017 7644
rect 12041 7642 12097 7644
rect 12121 7642 12177 7644
rect 12201 7642 12257 7644
rect 11961 7590 12007 7642
rect 12007 7590 12017 7642
rect 12041 7590 12071 7642
rect 12071 7590 12083 7642
rect 12083 7590 12097 7642
rect 12121 7590 12135 7642
rect 12135 7590 12147 7642
rect 12147 7590 12177 7642
rect 12201 7590 12211 7642
rect 12211 7590 12257 7642
rect 11961 7588 12017 7590
rect 12041 7588 12097 7590
rect 12121 7588 12177 7590
rect 12201 7588 12257 7590
rect 11702 6996 11758 7032
rect 11702 6976 11704 6996
rect 11704 6976 11756 6996
rect 11756 6976 11758 6996
rect 11886 6840 11942 6896
rect 12162 6724 12218 6760
rect 12162 6704 12164 6724
rect 12164 6704 12216 6724
rect 12216 6704 12218 6724
rect 11702 6604 11704 6624
rect 11704 6604 11756 6624
rect 11756 6604 11758 6624
rect 11702 6568 11758 6604
rect 11961 6554 12017 6556
rect 12041 6554 12097 6556
rect 12121 6554 12177 6556
rect 12201 6554 12257 6556
rect 11961 6502 12007 6554
rect 12007 6502 12017 6554
rect 12041 6502 12071 6554
rect 12071 6502 12083 6554
rect 12083 6502 12097 6554
rect 12121 6502 12135 6554
rect 12135 6502 12147 6554
rect 12147 6502 12177 6554
rect 12201 6502 12211 6554
rect 12211 6502 12257 6554
rect 11961 6500 12017 6502
rect 12041 6500 12097 6502
rect 12121 6500 12177 6502
rect 12201 6500 12257 6502
rect 11702 6452 11758 6488
rect 11702 6432 11704 6452
rect 11704 6432 11756 6452
rect 11756 6432 11758 6452
rect 4256 5466 4312 5468
rect 4336 5466 4392 5468
rect 4416 5466 4472 5468
rect 4496 5466 4552 5468
rect 4256 5414 4302 5466
rect 4302 5414 4312 5466
rect 4336 5414 4366 5466
rect 4366 5414 4378 5466
rect 4378 5414 4392 5466
rect 4416 5414 4430 5466
rect 4430 5414 4442 5466
rect 4442 5414 4472 5466
rect 4496 5414 4506 5466
rect 4506 5414 4552 5466
rect 4256 5412 4312 5414
rect 4336 5412 4392 5414
rect 4416 5412 4472 5414
rect 4496 5412 4552 5414
rect 11961 5466 12017 5468
rect 12041 5466 12097 5468
rect 12121 5466 12177 5468
rect 12201 5466 12257 5468
rect 11961 5414 12007 5466
rect 12007 5414 12017 5466
rect 12041 5414 12071 5466
rect 12071 5414 12083 5466
rect 12083 5414 12097 5466
rect 12121 5414 12135 5466
rect 12135 5414 12147 5466
rect 12147 5414 12177 5466
rect 12201 5414 12211 5466
rect 12211 5414 12257 5466
rect 11961 5412 12017 5414
rect 12041 5412 12097 5414
rect 12121 5412 12177 5414
rect 12201 5412 12257 5414
rect 8108 4922 8164 4924
rect 8188 4922 8244 4924
rect 8268 4922 8324 4924
rect 8348 4922 8404 4924
rect 8108 4870 8154 4922
rect 8154 4870 8164 4922
rect 8188 4870 8218 4922
rect 8218 4870 8230 4922
rect 8230 4870 8244 4922
rect 8268 4870 8282 4922
rect 8282 4870 8294 4922
rect 8294 4870 8324 4922
rect 8348 4870 8358 4922
rect 8358 4870 8404 4922
rect 8108 4868 8164 4870
rect 8188 4868 8244 4870
rect 8268 4868 8324 4870
rect 8348 4868 8404 4870
rect 4256 4378 4312 4380
rect 4336 4378 4392 4380
rect 4416 4378 4472 4380
rect 4496 4378 4552 4380
rect 4256 4326 4302 4378
rect 4302 4326 4312 4378
rect 4336 4326 4366 4378
rect 4366 4326 4378 4378
rect 4378 4326 4392 4378
rect 4416 4326 4430 4378
rect 4430 4326 4442 4378
rect 4442 4326 4472 4378
rect 4496 4326 4506 4378
rect 4506 4326 4552 4378
rect 4256 4324 4312 4326
rect 4336 4324 4392 4326
rect 4416 4324 4472 4326
rect 4496 4324 4552 4326
rect 11961 4378 12017 4380
rect 12041 4378 12097 4380
rect 12121 4378 12177 4380
rect 12201 4378 12257 4380
rect 11961 4326 12007 4378
rect 12007 4326 12017 4378
rect 12041 4326 12071 4378
rect 12071 4326 12083 4378
rect 12083 4326 12097 4378
rect 12121 4326 12135 4378
rect 12135 4326 12147 4378
rect 12147 4326 12177 4378
rect 12201 4326 12211 4378
rect 12211 4326 12257 4378
rect 11961 4324 12017 4326
rect 12041 4324 12097 4326
rect 12121 4324 12177 4326
rect 12201 4324 12257 4326
rect 8108 3834 8164 3836
rect 8188 3834 8244 3836
rect 8268 3834 8324 3836
rect 8348 3834 8404 3836
rect 8108 3782 8154 3834
rect 8154 3782 8164 3834
rect 8188 3782 8218 3834
rect 8218 3782 8230 3834
rect 8230 3782 8244 3834
rect 8268 3782 8282 3834
rect 8282 3782 8294 3834
rect 8294 3782 8324 3834
rect 8348 3782 8358 3834
rect 8358 3782 8404 3834
rect 8108 3780 8164 3782
rect 8188 3780 8244 3782
rect 8268 3780 8324 3782
rect 8348 3780 8404 3782
rect 4256 3290 4312 3292
rect 4336 3290 4392 3292
rect 4416 3290 4472 3292
rect 4496 3290 4552 3292
rect 4256 3238 4302 3290
rect 4302 3238 4312 3290
rect 4336 3238 4366 3290
rect 4366 3238 4378 3290
rect 4378 3238 4392 3290
rect 4416 3238 4430 3290
rect 4430 3238 4442 3290
rect 4442 3238 4472 3290
rect 4496 3238 4506 3290
rect 4506 3238 4552 3290
rect 4256 3236 4312 3238
rect 4336 3236 4392 3238
rect 4416 3236 4472 3238
rect 4496 3236 4552 3238
rect 8108 2746 8164 2748
rect 8188 2746 8244 2748
rect 8268 2746 8324 2748
rect 8348 2746 8404 2748
rect 8108 2694 8154 2746
rect 8154 2694 8164 2746
rect 8188 2694 8218 2746
rect 8218 2694 8230 2746
rect 8230 2694 8244 2746
rect 8268 2694 8282 2746
rect 8282 2694 8294 2746
rect 8294 2694 8324 2746
rect 8348 2694 8358 2746
rect 8358 2694 8404 2746
rect 8108 2692 8164 2694
rect 8188 2692 8244 2694
rect 8268 2692 8324 2694
rect 8348 2692 8404 2694
rect 4256 2202 4312 2204
rect 4336 2202 4392 2204
rect 4416 2202 4472 2204
rect 4496 2202 4552 2204
rect 4256 2150 4302 2202
rect 4302 2150 4312 2202
rect 4336 2150 4366 2202
rect 4366 2150 4378 2202
rect 4378 2150 4392 2202
rect 4416 2150 4430 2202
rect 4430 2150 4442 2202
rect 4442 2150 4472 2202
rect 4496 2150 4506 2202
rect 4506 2150 4552 2202
rect 4256 2148 4312 2150
rect 4336 2148 4392 2150
rect 4416 2148 4472 2150
rect 4496 2148 4552 2150
rect 8108 1658 8164 1660
rect 8188 1658 8244 1660
rect 8268 1658 8324 1660
rect 8348 1658 8404 1660
rect 8108 1606 8154 1658
rect 8154 1606 8164 1658
rect 8188 1606 8218 1658
rect 8218 1606 8230 1658
rect 8230 1606 8244 1658
rect 8268 1606 8282 1658
rect 8282 1606 8294 1658
rect 8294 1606 8324 1658
rect 8348 1606 8358 1658
rect 8358 1606 8404 1658
rect 8108 1604 8164 1606
rect 8188 1604 8244 1606
rect 8268 1604 8324 1606
rect 8348 1604 8404 1606
rect 4256 1114 4312 1116
rect 4336 1114 4392 1116
rect 4416 1114 4472 1116
rect 4496 1114 4552 1116
rect 4256 1062 4302 1114
rect 4302 1062 4312 1114
rect 4336 1062 4366 1114
rect 4366 1062 4378 1114
rect 4378 1062 4392 1114
rect 4416 1062 4430 1114
rect 4430 1062 4442 1114
rect 4442 1062 4472 1114
rect 4496 1062 4506 1114
rect 4506 1062 4552 1114
rect 4256 1060 4312 1062
rect 4336 1060 4392 1062
rect 4416 1060 4472 1062
rect 4496 1060 4552 1062
rect 8108 570 8164 572
rect 8188 570 8244 572
rect 8268 570 8324 572
rect 8348 570 8404 572
rect 8108 518 8154 570
rect 8154 518 8164 570
rect 8188 518 8218 570
rect 8218 518 8230 570
rect 8230 518 8244 570
rect 8268 518 8282 570
rect 8282 518 8294 570
rect 8294 518 8324 570
rect 8348 518 8358 570
rect 8358 518 8404 570
rect 8108 516 8164 518
rect 8188 516 8244 518
rect 8268 516 8324 518
rect 8348 516 8404 518
rect 11961 3290 12017 3292
rect 12041 3290 12097 3292
rect 12121 3290 12177 3292
rect 12201 3290 12257 3292
rect 11961 3238 12007 3290
rect 12007 3238 12017 3290
rect 12041 3238 12071 3290
rect 12071 3238 12083 3290
rect 12083 3238 12097 3290
rect 12121 3238 12135 3290
rect 12135 3238 12147 3290
rect 12147 3238 12177 3290
rect 12201 3238 12211 3290
rect 12211 3238 12257 3290
rect 11961 3236 12017 3238
rect 12041 3236 12097 3238
rect 12121 3236 12177 3238
rect 12201 3236 12257 3238
rect 13082 8200 13138 8256
rect 12990 7928 13046 7984
rect 12898 7792 12954 7848
rect 12806 6840 12862 6896
rect 15813 11450 15869 11452
rect 15893 11450 15949 11452
rect 15973 11450 16029 11452
rect 16053 11450 16109 11452
rect 15813 11398 15859 11450
rect 15859 11398 15869 11450
rect 15893 11398 15923 11450
rect 15923 11398 15935 11450
rect 15935 11398 15949 11450
rect 15973 11398 15987 11450
rect 15987 11398 15999 11450
rect 15999 11398 16029 11450
rect 16053 11398 16063 11450
rect 16063 11398 16109 11450
rect 15813 11396 15869 11398
rect 15893 11396 15949 11398
rect 15973 11396 16029 11398
rect 16053 11396 16109 11398
rect 15813 10362 15869 10364
rect 15893 10362 15949 10364
rect 15973 10362 16029 10364
rect 16053 10362 16109 10364
rect 15813 10310 15859 10362
rect 15859 10310 15869 10362
rect 15893 10310 15923 10362
rect 15923 10310 15935 10362
rect 15935 10310 15949 10362
rect 15973 10310 15987 10362
rect 15987 10310 15999 10362
rect 15999 10310 16029 10362
rect 16053 10310 16063 10362
rect 16063 10310 16109 10362
rect 15813 10308 15869 10310
rect 15893 10308 15949 10310
rect 15973 10308 16029 10310
rect 16053 10308 16109 10310
rect 15566 9696 15622 9752
rect 14094 8064 14150 8120
rect 15813 9274 15869 9276
rect 15893 9274 15949 9276
rect 15973 9274 16029 9276
rect 16053 9274 16109 9276
rect 15813 9222 15859 9274
rect 15859 9222 15869 9274
rect 15893 9222 15923 9274
rect 15923 9222 15935 9274
rect 15935 9222 15949 9274
rect 15973 9222 15987 9274
rect 15987 9222 15999 9274
rect 15999 9222 16029 9274
rect 16053 9222 16063 9274
rect 16063 9222 16109 9274
rect 15813 9220 15869 9222
rect 15893 9220 15949 9222
rect 15973 9220 16029 9222
rect 16053 9220 16109 9222
rect 15813 8186 15869 8188
rect 15893 8186 15949 8188
rect 15973 8186 16029 8188
rect 16053 8186 16109 8188
rect 15813 8134 15859 8186
rect 15859 8134 15869 8186
rect 15893 8134 15923 8186
rect 15923 8134 15935 8186
rect 15935 8134 15949 8186
rect 15973 8134 15987 8186
rect 15987 8134 15999 8186
rect 15999 8134 16029 8186
rect 16053 8134 16063 8186
rect 16063 8134 16109 8186
rect 15813 8132 15869 8134
rect 15893 8132 15949 8134
rect 15973 8132 16029 8134
rect 16053 8132 16109 8134
rect 11961 2202 12017 2204
rect 12041 2202 12097 2204
rect 12121 2202 12177 2204
rect 12201 2202 12257 2204
rect 11961 2150 12007 2202
rect 12007 2150 12017 2202
rect 12041 2150 12071 2202
rect 12071 2150 12083 2202
rect 12083 2150 12097 2202
rect 12121 2150 12135 2202
rect 12135 2150 12147 2202
rect 12147 2150 12177 2202
rect 12201 2150 12211 2202
rect 12211 2150 12257 2202
rect 11961 2148 12017 2150
rect 12041 2148 12097 2150
rect 12121 2148 12177 2150
rect 12201 2148 12257 2150
rect 11961 1114 12017 1116
rect 12041 1114 12097 1116
rect 12121 1114 12177 1116
rect 12201 1114 12257 1116
rect 11961 1062 12007 1114
rect 12007 1062 12017 1114
rect 12041 1062 12071 1114
rect 12071 1062 12083 1114
rect 12083 1062 12097 1114
rect 12121 1062 12135 1114
rect 12135 1062 12147 1114
rect 12147 1062 12177 1114
rect 12201 1062 12211 1114
rect 12211 1062 12257 1114
rect 11961 1060 12017 1062
rect 12041 1060 12097 1062
rect 12121 1060 12177 1062
rect 12201 1060 12257 1062
rect 15813 7098 15869 7100
rect 15893 7098 15949 7100
rect 15973 7098 16029 7100
rect 16053 7098 16109 7100
rect 15813 7046 15859 7098
rect 15859 7046 15869 7098
rect 15893 7046 15923 7098
rect 15923 7046 15935 7098
rect 15935 7046 15949 7098
rect 15973 7046 15987 7098
rect 15987 7046 15999 7098
rect 15999 7046 16029 7098
rect 16053 7046 16063 7098
rect 16063 7046 16109 7098
rect 15813 7044 15869 7046
rect 15893 7044 15949 7046
rect 15973 7044 16029 7046
rect 16053 7044 16109 7046
rect 15813 6010 15869 6012
rect 15893 6010 15949 6012
rect 15973 6010 16029 6012
rect 16053 6010 16109 6012
rect 15813 5958 15859 6010
rect 15859 5958 15869 6010
rect 15893 5958 15923 6010
rect 15923 5958 15935 6010
rect 15935 5958 15949 6010
rect 15973 5958 15987 6010
rect 15987 5958 15999 6010
rect 15999 5958 16029 6010
rect 16053 5958 16063 6010
rect 16063 5958 16109 6010
rect 15813 5956 15869 5958
rect 15893 5956 15949 5958
rect 15973 5956 16029 5958
rect 16053 5956 16109 5958
rect 15813 4922 15869 4924
rect 15893 4922 15949 4924
rect 15973 4922 16029 4924
rect 16053 4922 16109 4924
rect 15813 4870 15859 4922
rect 15859 4870 15869 4922
rect 15893 4870 15923 4922
rect 15923 4870 15935 4922
rect 15935 4870 15949 4922
rect 15973 4870 15987 4922
rect 15987 4870 15999 4922
rect 15999 4870 16029 4922
rect 16053 4870 16063 4922
rect 16063 4870 16109 4922
rect 15813 4868 15869 4870
rect 15893 4868 15949 4870
rect 15973 4868 16029 4870
rect 16053 4868 16109 4870
rect 15474 3984 15530 4040
rect 15813 3834 15869 3836
rect 15893 3834 15949 3836
rect 15973 3834 16029 3836
rect 16053 3834 16109 3836
rect 15813 3782 15859 3834
rect 15859 3782 15869 3834
rect 15893 3782 15923 3834
rect 15923 3782 15935 3834
rect 15935 3782 15949 3834
rect 15973 3782 15987 3834
rect 15987 3782 15999 3834
rect 15999 3782 16029 3834
rect 16053 3782 16063 3834
rect 16063 3782 16109 3834
rect 15813 3780 15869 3782
rect 15893 3780 15949 3782
rect 15973 3780 16029 3782
rect 16053 3780 16109 3782
rect 15813 2746 15869 2748
rect 15893 2746 15949 2748
rect 15973 2746 16029 2748
rect 16053 2746 16109 2748
rect 15813 2694 15859 2746
rect 15859 2694 15869 2746
rect 15893 2694 15923 2746
rect 15923 2694 15935 2746
rect 15935 2694 15949 2746
rect 15973 2694 15987 2746
rect 15987 2694 15999 2746
rect 15999 2694 16029 2746
rect 16053 2694 16063 2746
rect 16063 2694 16109 2746
rect 15813 2692 15869 2694
rect 15893 2692 15949 2694
rect 15973 2692 16029 2694
rect 16053 2692 16109 2694
rect 15813 1658 15869 1660
rect 15893 1658 15949 1660
rect 15973 1658 16029 1660
rect 16053 1658 16109 1660
rect 15813 1606 15859 1658
rect 15859 1606 15869 1658
rect 15893 1606 15923 1658
rect 15923 1606 15935 1658
rect 15935 1606 15949 1658
rect 15973 1606 15987 1658
rect 15987 1606 15999 1658
rect 15999 1606 16029 1658
rect 16053 1606 16063 1658
rect 16063 1606 16109 1658
rect 15813 1604 15869 1606
rect 15893 1604 15949 1606
rect 15973 1604 16029 1606
rect 16053 1604 16109 1606
rect 15813 570 15869 572
rect 15893 570 15949 572
rect 15973 570 16029 572
rect 16053 570 16109 572
rect 15813 518 15859 570
rect 15859 518 15869 570
rect 15893 518 15923 570
rect 15923 518 15935 570
rect 15935 518 15949 570
rect 15973 518 15987 570
rect 15987 518 15999 570
rect 15999 518 16029 570
rect 16053 518 16063 570
rect 16063 518 16109 570
rect 15813 516 15869 518
rect 15893 516 15949 518
rect 15973 516 16029 518
rect 16053 516 16109 518
rect 19666 16346 19722 16348
rect 19746 16346 19802 16348
rect 19826 16346 19882 16348
rect 19906 16346 19962 16348
rect 19666 16294 19712 16346
rect 19712 16294 19722 16346
rect 19746 16294 19776 16346
rect 19776 16294 19788 16346
rect 19788 16294 19802 16346
rect 19826 16294 19840 16346
rect 19840 16294 19852 16346
rect 19852 16294 19882 16346
rect 19906 16294 19916 16346
rect 19916 16294 19962 16346
rect 19666 16292 19722 16294
rect 19746 16292 19802 16294
rect 19826 16292 19882 16294
rect 19906 16292 19962 16294
rect 19666 15258 19722 15260
rect 19746 15258 19802 15260
rect 19826 15258 19882 15260
rect 19906 15258 19962 15260
rect 19666 15206 19712 15258
rect 19712 15206 19722 15258
rect 19746 15206 19776 15258
rect 19776 15206 19788 15258
rect 19788 15206 19802 15258
rect 19826 15206 19840 15258
rect 19840 15206 19852 15258
rect 19852 15206 19882 15258
rect 19906 15206 19916 15258
rect 19916 15206 19962 15258
rect 19666 15204 19722 15206
rect 19746 15204 19802 15206
rect 19826 15204 19882 15206
rect 19906 15204 19962 15206
rect 19666 14170 19722 14172
rect 19746 14170 19802 14172
rect 19826 14170 19882 14172
rect 19906 14170 19962 14172
rect 19666 14118 19712 14170
rect 19712 14118 19722 14170
rect 19746 14118 19776 14170
rect 19776 14118 19788 14170
rect 19788 14118 19802 14170
rect 19826 14118 19840 14170
rect 19840 14118 19852 14170
rect 19852 14118 19882 14170
rect 19906 14118 19916 14170
rect 19916 14118 19962 14170
rect 19666 14116 19722 14118
rect 19746 14116 19802 14118
rect 19826 14116 19882 14118
rect 19906 14116 19962 14118
rect 19666 13082 19722 13084
rect 19746 13082 19802 13084
rect 19826 13082 19882 13084
rect 19906 13082 19962 13084
rect 19666 13030 19712 13082
rect 19712 13030 19722 13082
rect 19746 13030 19776 13082
rect 19776 13030 19788 13082
rect 19788 13030 19802 13082
rect 19826 13030 19840 13082
rect 19840 13030 19852 13082
rect 19852 13030 19882 13082
rect 19906 13030 19916 13082
rect 19916 13030 19962 13082
rect 19666 13028 19722 13030
rect 19746 13028 19802 13030
rect 19826 13028 19882 13030
rect 19906 13028 19962 13030
rect 19666 11994 19722 11996
rect 19746 11994 19802 11996
rect 19826 11994 19882 11996
rect 19906 11994 19962 11996
rect 19666 11942 19712 11994
rect 19712 11942 19722 11994
rect 19746 11942 19776 11994
rect 19776 11942 19788 11994
rect 19788 11942 19802 11994
rect 19826 11942 19840 11994
rect 19840 11942 19852 11994
rect 19852 11942 19882 11994
rect 19906 11942 19916 11994
rect 19916 11942 19962 11994
rect 19666 11940 19722 11942
rect 19746 11940 19802 11942
rect 19826 11940 19882 11942
rect 19906 11940 19962 11942
rect 23518 19066 23574 19068
rect 23598 19066 23654 19068
rect 23678 19066 23734 19068
rect 23758 19066 23814 19068
rect 23518 19014 23564 19066
rect 23564 19014 23574 19066
rect 23598 19014 23628 19066
rect 23628 19014 23640 19066
rect 23640 19014 23654 19066
rect 23678 19014 23692 19066
rect 23692 19014 23704 19066
rect 23704 19014 23734 19066
rect 23758 19014 23768 19066
rect 23768 19014 23814 19066
rect 23518 19012 23574 19014
rect 23598 19012 23654 19014
rect 23678 19012 23734 19014
rect 23758 19012 23814 19014
rect 31223 19066 31279 19068
rect 31303 19066 31359 19068
rect 31383 19066 31439 19068
rect 31463 19066 31519 19068
rect 31223 19014 31269 19066
rect 31269 19014 31279 19066
rect 31303 19014 31333 19066
rect 31333 19014 31345 19066
rect 31345 19014 31359 19066
rect 31383 19014 31397 19066
rect 31397 19014 31409 19066
rect 31409 19014 31439 19066
rect 31463 19014 31473 19066
rect 31473 19014 31519 19066
rect 31223 19012 31279 19014
rect 31303 19012 31359 19014
rect 31383 19012 31439 19014
rect 31463 19012 31519 19014
rect 27371 18522 27427 18524
rect 27451 18522 27507 18524
rect 27531 18522 27587 18524
rect 27611 18522 27667 18524
rect 27371 18470 27417 18522
rect 27417 18470 27427 18522
rect 27451 18470 27481 18522
rect 27481 18470 27493 18522
rect 27493 18470 27507 18522
rect 27531 18470 27545 18522
rect 27545 18470 27557 18522
rect 27557 18470 27587 18522
rect 27611 18470 27621 18522
rect 27621 18470 27667 18522
rect 27371 18468 27427 18470
rect 27451 18468 27507 18470
rect 27531 18468 27587 18470
rect 27611 18468 27667 18470
rect 23518 17978 23574 17980
rect 23598 17978 23654 17980
rect 23678 17978 23734 17980
rect 23758 17978 23814 17980
rect 23518 17926 23564 17978
rect 23564 17926 23574 17978
rect 23598 17926 23628 17978
rect 23628 17926 23640 17978
rect 23640 17926 23654 17978
rect 23678 17926 23692 17978
rect 23692 17926 23704 17978
rect 23704 17926 23734 17978
rect 23758 17926 23768 17978
rect 23768 17926 23814 17978
rect 23518 17924 23574 17926
rect 23598 17924 23654 17926
rect 23678 17924 23734 17926
rect 23758 17924 23814 17926
rect 31223 17978 31279 17980
rect 31303 17978 31359 17980
rect 31383 17978 31439 17980
rect 31463 17978 31519 17980
rect 31223 17926 31269 17978
rect 31269 17926 31279 17978
rect 31303 17926 31333 17978
rect 31333 17926 31345 17978
rect 31345 17926 31359 17978
rect 31383 17926 31397 17978
rect 31397 17926 31409 17978
rect 31409 17926 31439 17978
rect 31463 17926 31473 17978
rect 31473 17926 31519 17978
rect 31223 17924 31279 17926
rect 31303 17924 31359 17926
rect 31383 17924 31439 17926
rect 31463 17924 31519 17926
rect 27371 17434 27427 17436
rect 27451 17434 27507 17436
rect 27531 17434 27587 17436
rect 27611 17434 27667 17436
rect 27371 17382 27417 17434
rect 27417 17382 27427 17434
rect 27451 17382 27481 17434
rect 27481 17382 27493 17434
rect 27493 17382 27507 17434
rect 27531 17382 27545 17434
rect 27545 17382 27557 17434
rect 27557 17382 27587 17434
rect 27611 17382 27621 17434
rect 27621 17382 27667 17434
rect 27371 17380 27427 17382
rect 27451 17380 27507 17382
rect 27531 17380 27587 17382
rect 27611 17380 27667 17382
rect 23518 16890 23574 16892
rect 23598 16890 23654 16892
rect 23678 16890 23734 16892
rect 23758 16890 23814 16892
rect 23518 16838 23564 16890
rect 23564 16838 23574 16890
rect 23598 16838 23628 16890
rect 23628 16838 23640 16890
rect 23640 16838 23654 16890
rect 23678 16838 23692 16890
rect 23692 16838 23704 16890
rect 23704 16838 23734 16890
rect 23758 16838 23768 16890
rect 23768 16838 23814 16890
rect 23518 16836 23574 16838
rect 23598 16836 23654 16838
rect 23678 16836 23734 16838
rect 23758 16836 23814 16838
rect 31223 16890 31279 16892
rect 31303 16890 31359 16892
rect 31383 16890 31439 16892
rect 31463 16890 31519 16892
rect 31223 16838 31269 16890
rect 31269 16838 31279 16890
rect 31303 16838 31333 16890
rect 31333 16838 31345 16890
rect 31345 16838 31359 16890
rect 31383 16838 31397 16890
rect 31397 16838 31409 16890
rect 31409 16838 31439 16890
rect 31463 16838 31473 16890
rect 31473 16838 31519 16890
rect 31223 16836 31279 16838
rect 31303 16836 31359 16838
rect 31383 16836 31439 16838
rect 31463 16836 31519 16838
rect 27371 16346 27427 16348
rect 27451 16346 27507 16348
rect 27531 16346 27587 16348
rect 27611 16346 27667 16348
rect 27371 16294 27417 16346
rect 27417 16294 27427 16346
rect 27451 16294 27481 16346
rect 27481 16294 27493 16346
rect 27493 16294 27507 16346
rect 27531 16294 27545 16346
rect 27545 16294 27557 16346
rect 27557 16294 27587 16346
rect 27611 16294 27621 16346
rect 27621 16294 27667 16346
rect 27371 16292 27427 16294
rect 27451 16292 27507 16294
rect 27531 16292 27587 16294
rect 27611 16292 27667 16294
rect 23518 15802 23574 15804
rect 23598 15802 23654 15804
rect 23678 15802 23734 15804
rect 23758 15802 23814 15804
rect 23518 15750 23564 15802
rect 23564 15750 23574 15802
rect 23598 15750 23628 15802
rect 23628 15750 23640 15802
rect 23640 15750 23654 15802
rect 23678 15750 23692 15802
rect 23692 15750 23704 15802
rect 23704 15750 23734 15802
rect 23758 15750 23768 15802
rect 23768 15750 23814 15802
rect 23518 15748 23574 15750
rect 23598 15748 23654 15750
rect 23678 15748 23734 15750
rect 23758 15748 23814 15750
rect 31223 15802 31279 15804
rect 31303 15802 31359 15804
rect 31383 15802 31439 15804
rect 31463 15802 31519 15804
rect 31223 15750 31269 15802
rect 31269 15750 31279 15802
rect 31303 15750 31333 15802
rect 31333 15750 31345 15802
rect 31345 15750 31359 15802
rect 31383 15750 31397 15802
rect 31397 15750 31409 15802
rect 31409 15750 31439 15802
rect 31463 15750 31473 15802
rect 31473 15750 31519 15802
rect 31223 15748 31279 15750
rect 31303 15748 31359 15750
rect 31383 15748 31439 15750
rect 31463 15748 31519 15750
rect 27371 15258 27427 15260
rect 27451 15258 27507 15260
rect 27531 15258 27587 15260
rect 27611 15258 27667 15260
rect 27371 15206 27417 15258
rect 27417 15206 27427 15258
rect 27451 15206 27481 15258
rect 27481 15206 27493 15258
rect 27493 15206 27507 15258
rect 27531 15206 27545 15258
rect 27545 15206 27557 15258
rect 27557 15206 27587 15258
rect 27611 15206 27621 15258
rect 27621 15206 27667 15258
rect 27371 15204 27427 15206
rect 27451 15204 27507 15206
rect 27531 15204 27587 15206
rect 27611 15204 27667 15206
rect 23518 14714 23574 14716
rect 23598 14714 23654 14716
rect 23678 14714 23734 14716
rect 23758 14714 23814 14716
rect 23518 14662 23564 14714
rect 23564 14662 23574 14714
rect 23598 14662 23628 14714
rect 23628 14662 23640 14714
rect 23640 14662 23654 14714
rect 23678 14662 23692 14714
rect 23692 14662 23704 14714
rect 23704 14662 23734 14714
rect 23758 14662 23768 14714
rect 23768 14662 23814 14714
rect 23518 14660 23574 14662
rect 23598 14660 23654 14662
rect 23678 14660 23734 14662
rect 23758 14660 23814 14662
rect 31223 14714 31279 14716
rect 31303 14714 31359 14716
rect 31383 14714 31439 14716
rect 31463 14714 31519 14716
rect 31223 14662 31269 14714
rect 31269 14662 31279 14714
rect 31303 14662 31333 14714
rect 31333 14662 31345 14714
rect 31345 14662 31359 14714
rect 31383 14662 31397 14714
rect 31397 14662 31409 14714
rect 31409 14662 31439 14714
rect 31463 14662 31473 14714
rect 31473 14662 31519 14714
rect 31223 14660 31279 14662
rect 31303 14660 31359 14662
rect 31383 14660 31439 14662
rect 31463 14660 31519 14662
rect 27371 14170 27427 14172
rect 27451 14170 27507 14172
rect 27531 14170 27587 14172
rect 27611 14170 27667 14172
rect 27371 14118 27417 14170
rect 27417 14118 27427 14170
rect 27451 14118 27481 14170
rect 27481 14118 27493 14170
rect 27493 14118 27507 14170
rect 27531 14118 27545 14170
rect 27545 14118 27557 14170
rect 27557 14118 27587 14170
rect 27611 14118 27621 14170
rect 27621 14118 27667 14170
rect 27371 14116 27427 14118
rect 27451 14116 27507 14118
rect 27531 14116 27587 14118
rect 27611 14116 27667 14118
rect 23518 13626 23574 13628
rect 23598 13626 23654 13628
rect 23678 13626 23734 13628
rect 23758 13626 23814 13628
rect 23518 13574 23564 13626
rect 23564 13574 23574 13626
rect 23598 13574 23628 13626
rect 23628 13574 23640 13626
rect 23640 13574 23654 13626
rect 23678 13574 23692 13626
rect 23692 13574 23704 13626
rect 23704 13574 23734 13626
rect 23758 13574 23768 13626
rect 23768 13574 23814 13626
rect 23518 13572 23574 13574
rect 23598 13572 23654 13574
rect 23678 13572 23734 13574
rect 23758 13572 23814 13574
rect 31223 13626 31279 13628
rect 31303 13626 31359 13628
rect 31383 13626 31439 13628
rect 31463 13626 31519 13628
rect 31223 13574 31269 13626
rect 31269 13574 31279 13626
rect 31303 13574 31333 13626
rect 31333 13574 31345 13626
rect 31345 13574 31359 13626
rect 31383 13574 31397 13626
rect 31397 13574 31409 13626
rect 31409 13574 31439 13626
rect 31463 13574 31473 13626
rect 31473 13574 31519 13626
rect 31223 13572 31279 13574
rect 31303 13572 31359 13574
rect 31383 13572 31439 13574
rect 31463 13572 31519 13574
rect 27371 13082 27427 13084
rect 27451 13082 27507 13084
rect 27531 13082 27587 13084
rect 27611 13082 27667 13084
rect 27371 13030 27417 13082
rect 27417 13030 27427 13082
rect 27451 13030 27481 13082
rect 27481 13030 27493 13082
rect 27493 13030 27507 13082
rect 27531 13030 27545 13082
rect 27545 13030 27557 13082
rect 27557 13030 27587 13082
rect 27611 13030 27621 13082
rect 27621 13030 27667 13082
rect 27371 13028 27427 13030
rect 27451 13028 27507 13030
rect 27531 13028 27587 13030
rect 27611 13028 27667 13030
rect 23518 12538 23574 12540
rect 23598 12538 23654 12540
rect 23678 12538 23734 12540
rect 23758 12538 23814 12540
rect 23518 12486 23564 12538
rect 23564 12486 23574 12538
rect 23598 12486 23628 12538
rect 23628 12486 23640 12538
rect 23640 12486 23654 12538
rect 23678 12486 23692 12538
rect 23692 12486 23704 12538
rect 23704 12486 23734 12538
rect 23758 12486 23768 12538
rect 23768 12486 23814 12538
rect 23518 12484 23574 12486
rect 23598 12484 23654 12486
rect 23678 12484 23734 12486
rect 23758 12484 23814 12486
rect 31223 12538 31279 12540
rect 31303 12538 31359 12540
rect 31383 12538 31439 12540
rect 31463 12538 31519 12540
rect 31223 12486 31269 12538
rect 31269 12486 31279 12538
rect 31303 12486 31333 12538
rect 31333 12486 31345 12538
rect 31345 12486 31359 12538
rect 31383 12486 31397 12538
rect 31397 12486 31409 12538
rect 31409 12486 31439 12538
rect 31463 12486 31473 12538
rect 31473 12486 31519 12538
rect 31223 12484 31279 12486
rect 31303 12484 31359 12486
rect 31383 12484 31439 12486
rect 31463 12484 31519 12486
rect 27371 11994 27427 11996
rect 27451 11994 27507 11996
rect 27531 11994 27587 11996
rect 27611 11994 27667 11996
rect 27371 11942 27417 11994
rect 27417 11942 27427 11994
rect 27451 11942 27481 11994
rect 27481 11942 27493 11994
rect 27493 11942 27507 11994
rect 27531 11942 27545 11994
rect 27545 11942 27557 11994
rect 27557 11942 27587 11994
rect 27611 11942 27621 11994
rect 27621 11942 27667 11994
rect 27371 11940 27427 11942
rect 27451 11940 27507 11942
rect 27531 11940 27587 11942
rect 27611 11940 27667 11942
rect 23518 11450 23574 11452
rect 23598 11450 23654 11452
rect 23678 11450 23734 11452
rect 23758 11450 23814 11452
rect 23518 11398 23564 11450
rect 23564 11398 23574 11450
rect 23598 11398 23628 11450
rect 23628 11398 23640 11450
rect 23640 11398 23654 11450
rect 23678 11398 23692 11450
rect 23692 11398 23704 11450
rect 23704 11398 23734 11450
rect 23758 11398 23768 11450
rect 23768 11398 23814 11450
rect 23518 11396 23574 11398
rect 23598 11396 23654 11398
rect 23678 11396 23734 11398
rect 23758 11396 23814 11398
rect 31223 11450 31279 11452
rect 31303 11450 31359 11452
rect 31383 11450 31439 11452
rect 31463 11450 31519 11452
rect 31223 11398 31269 11450
rect 31269 11398 31279 11450
rect 31303 11398 31333 11450
rect 31333 11398 31345 11450
rect 31345 11398 31359 11450
rect 31383 11398 31397 11450
rect 31397 11398 31409 11450
rect 31409 11398 31439 11450
rect 31463 11398 31473 11450
rect 31473 11398 31519 11450
rect 31223 11396 31279 11398
rect 31303 11396 31359 11398
rect 31383 11396 31439 11398
rect 31463 11396 31519 11398
rect 19666 10906 19722 10908
rect 19746 10906 19802 10908
rect 19826 10906 19882 10908
rect 19906 10906 19962 10908
rect 19666 10854 19712 10906
rect 19712 10854 19722 10906
rect 19746 10854 19776 10906
rect 19776 10854 19788 10906
rect 19788 10854 19802 10906
rect 19826 10854 19840 10906
rect 19840 10854 19852 10906
rect 19852 10854 19882 10906
rect 19906 10854 19916 10906
rect 19916 10854 19962 10906
rect 19666 10852 19722 10854
rect 19746 10852 19802 10854
rect 19826 10852 19882 10854
rect 19906 10852 19962 10854
rect 27371 10906 27427 10908
rect 27451 10906 27507 10908
rect 27531 10906 27587 10908
rect 27611 10906 27667 10908
rect 27371 10854 27417 10906
rect 27417 10854 27427 10906
rect 27451 10854 27481 10906
rect 27481 10854 27493 10906
rect 27493 10854 27507 10906
rect 27531 10854 27545 10906
rect 27545 10854 27557 10906
rect 27557 10854 27587 10906
rect 27611 10854 27621 10906
rect 27621 10854 27667 10906
rect 27371 10852 27427 10854
rect 27451 10852 27507 10854
rect 27531 10852 27587 10854
rect 27611 10852 27667 10854
rect 19666 9818 19722 9820
rect 19746 9818 19802 9820
rect 19826 9818 19882 9820
rect 19906 9818 19962 9820
rect 19666 9766 19712 9818
rect 19712 9766 19722 9818
rect 19746 9766 19776 9818
rect 19776 9766 19788 9818
rect 19788 9766 19802 9818
rect 19826 9766 19840 9818
rect 19840 9766 19852 9818
rect 19852 9766 19882 9818
rect 19906 9766 19916 9818
rect 19916 9766 19962 9818
rect 19666 9764 19722 9766
rect 19746 9764 19802 9766
rect 19826 9764 19882 9766
rect 19906 9764 19962 9766
rect 23518 10362 23574 10364
rect 23598 10362 23654 10364
rect 23678 10362 23734 10364
rect 23758 10362 23814 10364
rect 23518 10310 23564 10362
rect 23564 10310 23574 10362
rect 23598 10310 23628 10362
rect 23628 10310 23640 10362
rect 23640 10310 23654 10362
rect 23678 10310 23692 10362
rect 23692 10310 23704 10362
rect 23704 10310 23734 10362
rect 23758 10310 23768 10362
rect 23768 10310 23814 10362
rect 23518 10308 23574 10310
rect 23598 10308 23654 10310
rect 23678 10308 23734 10310
rect 23758 10308 23814 10310
rect 31223 10362 31279 10364
rect 31303 10362 31359 10364
rect 31383 10362 31439 10364
rect 31463 10362 31519 10364
rect 31223 10310 31269 10362
rect 31269 10310 31279 10362
rect 31303 10310 31333 10362
rect 31333 10310 31345 10362
rect 31345 10310 31359 10362
rect 31383 10310 31397 10362
rect 31397 10310 31409 10362
rect 31409 10310 31439 10362
rect 31463 10310 31473 10362
rect 31473 10310 31519 10362
rect 31223 10308 31279 10310
rect 31303 10308 31359 10310
rect 31383 10308 31439 10310
rect 31463 10308 31519 10310
rect 31666 10240 31722 10296
rect 27371 9818 27427 9820
rect 27451 9818 27507 9820
rect 27531 9818 27587 9820
rect 27611 9818 27667 9820
rect 27371 9766 27417 9818
rect 27417 9766 27427 9818
rect 27451 9766 27481 9818
rect 27481 9766 27493 9818
rect 27493 9766 27507 9818
rect 27531 9766 27545 9818
rect 27545 9766 27557 9818
rect 27557 9766 27587 9818
rect 27611 9766 27621 9818
rect 27621 9766 27667 9818
rect 27371 9764 27427 9766
rect 27451 9764 27507 9766
rect 27531 9764 27587 9766
rect 27611 9764 27667 9766
rect 28262 9560 28318 9616
rect 23518 9274 23574 9276
rect 23598 9274 23654 9276
rect 23678 9274 23734 9276
rect 23758 9274 23814 9276
rect 23518 9222 23564 9274
rect 23564 9222 23574 9274
rect 23598 9222 23628 9274
rect 23628 9222 23640 9274
rect 23640 9222 23654 9274
rect 23678 9222 23692 9274
rect 23692 9222 23704 9274
rect 23704 9222 23734 9274
rect 23758 9222 23768 9274
rect 23768 9222 23814 9274
rect 23518 9220 23574 9222
rect 23598 9220 23654 9222
rect 23678 9220 23734 9222
rect 23758 9220 23814 9222
rect 31223 9274 31279 9276
rect 31303 9274 31359 9276
rect 31383 9274 31439 9276
rect 31463 9274 31519 9276
rect 31223 9222 31269 9274
rect 31269 9222 31279 9274
rect 31303 9222 31333 9274
rect 31333 9222 31345 9274
rect 31345 9222 31359 9274
rect 31383 9222 31397 9274
rect 31397 9222 31409 9274
rect 31409 9222 31439 9274
rect 31463 9222 31473 9274
rect 31473 9222 31519 9274
rect 31223 9220 31279 9222
rect 31303 9220 31359 9222
rect 31383 9220 31439 9222
rect 31463 9220 31519 9222
rect 19666 8730 19722 8732
rect 19746 8730 19802 8732
rect 19826 8730 19882 8732
rect 19906 8730 19962 8732
rect 19666 8678 19712 8730
rect 19712 8678 19722 8730
rect 19746 8678 19776 8730
rect 19776 8678 19788 8730
rect 19788 8678 19802 8730
rect 19826 8678 19840 8730
rect 19840 8678 19852 8730
rect 19852 8678 19882 8730
rect 19906 8678 19916 8730
rect 19916 8678 19962 8730
rect 19666 8676 19722 8678
rect 19746 8676 19802 8678
rect 19826 8676 19882 8678
rect 19906 8676 19962 8678
rect 19666 7642 19722 7644
rect 19746 7642 19802 7644
rect 19826 7642 19882 7644
rect 19906 7642 19962 7644
rect 19666 7590 19712 7642
rect 19712 7590 19722 7642
rect 19746 7590 19776 7642
rect 19776 7590 19788 7642
rect 19788 7590 19802 7642
rect 19826 7590 19840 7642
rect 19840 7590 19852 7642
rect 19852 7590 19882 7642
rect 19906 7590 19916 7642
rect 19916 7590 19962 7642
rect 19666 7588 19722 7590
rect 19746 7588 19802 7590
rect 19826 7588 19882 7590
rect 19906 7588 19962 7590
rect 19666 6554 19722 6556
rect 19746 6554 19802 6556
rect 19826 6554 19882 6556
rect 19906 6554 19962 6556
rect 19666 6502 19712 6554
rect 19712 6502 19722 6554
rect 19746 6502 19776 6554
rect 19776 6502 19788 6554
rect 19788 6502 19802 6554
rect 19826 6502 19840 6554
rect 19840 6502 19852 6554
rect 19852 6502 19882 6554
rect 19906 6502 19916 6554
rect 19916 6502 19962 6554
rect 19666 6500 19722 6502
rect 19746 6500 19802 6502
rect 19826 6500 19882 6502
rect 19906 6500 19962 6502
rect 19666 5466 19722 5468
rect 19746 5466 19802 5468
rect 19826 5466 19882 5468
rect 19906 5466 19962 5468
rect 19666 5414 19712 5466
rect 19712 5414 19722 5466
rect 19746 5414 19776 5466
rect 19776 5414 19788 5466
rect 19788 5414 19802 5466
rect 19826 5414 19840 5466
rect 19840 5414 19852 5466
rect 19852 5414 19882 5466
rect 19906 5414 19916 5466
rect 19916 5414 19962 5466
rect 19666 5412 19722 5414
rect 19746 5412 19802 5414
rect 19826 5412 19882 5414
rect 19906 5412 19962 5414
rect 19666 4378 19722 4380
rect 19746 4378 19802 4380
rect 19826 4378 19882 4380
rect 19906 4378 19962 4380
rect 19666 4326 19712 4378
rect 19712 4326 19722 4378
rect 19746 4326 19776 4378
rect 19776 4326 19788 4378
rect 19788 4326 19802 4378
rect 19826 4326 19840 4378
rect 19840 4326 19852 4378
rect 19852 4326 19882 4378
rect 19906 4326 19916 4378
rect 19916 4326 19962 4378
rect 19666 4324 19722 4326
rect 19746 4324 19802 4326
rect 19826 4324 19882 4326
rect 19906 4324 19962 4326
rect 19666 3290 19722 3292
rect 19746 3290 19802 3292
rect 19826 3290 19882 3292
rect 19906 3290 19962 3292
rect 19666 3238 19712 3290
rect 19712 3238 19722 3290
rect 19746 3238 19776 3290
rect 19776 3238 19788 3290
rect 19788 3238 19802 3290
rect 19826 3238 19840 3290
rect 19840 3238 19852 3290
rect 19852 3238 19882 3290
rect 19906 3238 19916 3290
rect 19916 3238 19962 3290
rect 19666 3236 19722 3238
rect 19746 3236 19802 3238
rect 19826 3236 19882 3238
rect 19906 3236 19962 3238
rect 19666 2202 19722 2204
rect 19746 2202 19802 2204
rect 19826 2202 19882 2204
rect 19906 2202 19962 2204
rect 19666 2150 19712 2202
rect 19712 2150 19722 2202
rect 19746 2150 19776 2202
rect 19776 2150 19788 2202
rect 19788 2150 19802 2202
rect 19826 2150 19840 2202
rect 19840 2150 19852 2202
rect 19852 2150 19882 2202
rect 19906 2150 19916 2202
rect 19916 2150 19962 2202
rect 19666 2148 19722 2150
rect 19746 2148 19802 2150
rect 19826 2148 19882 2150
rect 19906 2148 19962 2150
rect 19666 1114 19722 1116
rect 19746 1114 19802 1116
rect 19826 1114 19882 1116
rect 19906 1114 19962 1116
rect 19666 1062 19712 1114
rect 19712 1062 19722 1114
rect 19746 1062 19776 1114
rect 19776 1062 19788 1114
rect 19788 1062 19802 1114
rect 19826 1062 19840 1114
rect 19840 1062 19852 1114
rect 19852 1062 19882 1114
rect 19906 1062 19916 1114
rect 19916 1062 19962 1114
rect 19666 1060 19722 1062
rect 19746 1060 19802 1062
rect 19826 1060 19882 1062
rect 19906 1060 19962 1062
rect 28262 8900 28318 8936
rect 28262 8880 28264 8900
rect 28264 8880 28316 8900
rect 28316 8880 28318 8900
rect 27371 8730 27427 8732
rect 27451 8730 27507 8732
rect 27531 8730 27587 8732
rect 27611 8730 27667 8732
rect 27371 8678 27417 8730
rect 27417 8678 27427 8730
rect 27451 8678 27481 8730
rect 27481 8678 27493 8730
rect 27493 8678 27507 8730
rect 27531 8678 27545 8730
rect 27545 8678 27557 8730
rect 27557 8678 27587 8730
rect 27611 8678 27621 8730
rect 27621 8678 27667 8730
rect 27371 8676 27427 8678
rect 27451 8676 27507 8678
rect 27531 8676 27587 8678
rect 27611 8676 27667 8678
rect 23518 8186 23574 8188
rect 23598 8186 23654 8188
rect 23678 8186 23734 8188
rect 23758 8186 23814 8188
rect 23518 8134 23564 8186
rect 23564 8134 23574 8186
rect 23598 8134 23628 8186
rect 23628 8134 23640 8186
rect 23640 8134 23654 8186
rect 23678 8134 23692 8186
rect 23692 8134 23704 8186
rect 23704 8134 23734 8186
rect 23758 8134 23768 8186
rect 23768 8134 23814 8186
rect 23518 8132 23574 8134
rect 23598 8132 23654 8134
rect 23678 8132 23734 8134
rect 23758 8132 23814 8134
rect 31223 8186 31279 8188
rect 31303 8186 31359 8188
rect 31383 8186 31439 8188
rect 31463 8186 31519 8188
rect 31223 8134 31269 8186
rect 31269 8134 31279 8186
rect 31303 8134 31333 8186
rect 31333 8134 31345 8186
rect 31345 8134 31359 8186
rect 31383 8134 31397 8186
rect 31397 8134 31409 8186
rect 31409 8134 31439 8186
rect 31463 8134 31473 8186
rect 31473 8134 31519 8186
rect 31223 8132 31279 8134
rect 31303 8132 31359 8134
rect 31383 8132 31439 8134
rect 31463 8132 31519 8134
rect 27371 7642 27427 7644
rect 27451 7642 27507 7644
rect 27531 7642 27587 7644
rect 27611 7642 27667 7644
rect 27371 7590 27417 7642
rect 27417 7590 27427 7642
rect 27451 7590 27481 7642
rect 27481 7590 27493 7642
rect 27493 7590 27507 7642
rect 27531 7590 27545 7642
rect 27545 7590 27557 7642
rect 27557 7590 27587 7642
rect 27611 7590 27621 7642
rect 27621 7590 27667 7642
rect 27371 7588 27427 7590
rect 27451 7588 27507 7590
rect 27531 7588 27587 7590
rect 27611 7588 27667 7590
rect 23518 7098 23574 7100
rect 23598 7098 23654 7100
rect 23678 7098 23734 7100
rect 23758 7098 23814 7100
rect 23518 7046 23564 7098
rect 23564 7046 23574 7098
rect 23598 7046 23628 7098
rect 23628 7046 23640 7098
rect 23640 7046 23654 7098
rect 23678 7046 23692 7098
rect 23692 7046 23704 7098
rect 23704 7046 23734 7098
rect 23758 7046 23768 7098
rect 23768 7046 23814 7098
rect 23518 7044 23574 7046
rect 23598 7044 23654 7046
rect 23678 7044 23734 7046
rect 23758 7044 23814 7046
rect 31223 7098 31279 7100
rect 31303 7098 31359 7100
rect 31383 7098 31439 7100
rect 31463 7098 31519 7100
rect 31223 7046 31269 7098
rect 31269 7046 31279 7098
rect 31303 7046 31333 7098
rect 31333 7046 31345 7098
rect 31345 7046 31359 7098
rect 31383 7046 31397 7098
rect 31397 7046 31409 7098
rect 31409 7046 31439 7098
rect 31463 7046 31473 7098
rect 31473 7046 31519 7098
rect 31223 7044 31279 7046
rect 31303 7044 31359 7046
rect 31383 7044 31439 7046
rect 31463 7044 31519 7046
rect 27371 6554 27427 6556
rect 27451 6554 27507 6556
rect 27531 6554 27587 6556
rect 27611 6554 27667 6556
rect 27371 6502 27417 6554
rect 27417 6502 27427 6554
rect 27451 6502 27481 6554
rect 27481 6502 27493 6554
rect 27493 6502 27507 6554
rect 27531 6502 27545 6554
rect 27545 6502 27557 6554
rect 27557 6502 27587 6554
rect 27611 6502 27621 6554
rect 27621 6502 27667 6554
rect 27371 6500 27427 6502
rect 27451 6500 27507 6502
rect 27531 6500 27587 6502
rect 27611 6500 27667 6502
rect 23518 6010 23574 6012
rect 23598 6010 23654 6012
rect 23678 6010 23734 6012
rect 23758 6010 23814 6012
rect 23518 5958 23564 6010
rect 23564 5958 23574 6010
rect 23598 5958 23628 6010
rect 23628 5958 23640 6010
rect 23640 5958 23654 6010
rect 23678 5958 23692 6010
rect 23692 5958 23704 6010
rect 23704 5958 23734 6010
rect 23758 5958 23768 6010
rect 23768 5958 23814 6010
rect 23518 5956 23574 5958
rect 23598 5956 23654 5958
rect 23678 5956 23734 5958
rect 23758 5956 23814 5958
rect 31223 6010 31279 6012
rect 31303 6010 31359 6012
rect 31383 6010 31439 6012
rect 31463 6010 31519 6012
rect 31223 5958 31269 6010
rect 31269 5958 31279 6010
rect 31303 5958 31333 6010
rect 31333 5958 31345 6010
rect 31345 5958 31359 6010
rect 31383 5958 31397 6010
rect 31397 5958 31409 6010
rect 31409 5958 31439 6010
rect 31463 5958 31473 6010
rect 31473 5958 31519 6010
rect 31223 5956 31279 5958
rect 31303 5956 31359 5958
rect 31383 5956 31439 5958
rect 31463 5956 31519 5958
rect 27371 5466 27427 5468
rect 27451 5466 27507 5468
rect 27531 5466 27587 5468
rect 27611 5466 27667 5468
rect 27371 5414 27417 5466
rect 27417 5414 27427 5466
rect 27451 5414 27481 5466
rect 27481 5414 27493 5466
rect 27493 5414 27507 5466
rect 27531 5414 27545 5466
rect 27545 5414 27557 5466
rect 27557 5414 27587 5466
rect 27611 5414 27621 5466
rect 27621 5414 27667 5466
rect 27371 5412 27427 5414
rect 27451 5412 27507 5414
rect 27531 5412 27587 5414
rect 27611 5412 27667 5414
rect 23518 4922 23574 4924
rect 23598 4922 23654 4924
rect 23678 4922 23734 4924
rect 23758 4922 23814 4924
rect 23518 4870 23564 4922
rect 23564 4870 23574 4922
rect 23598 4870 23628 4922
rect 23628 4870 23640 4922
rect 23640 4870 23654 4922
rect 23678 4870 23692 4922
rect 23692 4870 23704 4922
rect 23704 4870 23734 4922
rect 23758 4870 23768 4922
rect 23768 4870 23814 4922
rect 23518 4868 23574 4870
rect 23598 4868 23654 4870
rect 23678 4868 23734 4870
rect 23758 4868 23814 4870
rect 31223 4922 31279 4924
rect 31303 4922 31359 4924
rect 31383 4922 31439 4924
rect 31463 4922 31519 4924
rect 31223 4870 31269 4922
rect 31269 4870 31279 4922
rect 31303 4870 31333 4922
rect 31333 4870 31345 4922
rect 31345 4870 31359 4922
rect 31383 4870 31397 4922
rect 31397 4870 31409 4922
rect 31409 4870 31439 4922
rect 31463 4870 31473 4922
rect 31473 4870 31519 4922
rect 31223 4868 31279 4870
rect 31303 4868 31359 4870
rect 31383 4868 31439 4870
rect 31463 4868 31519 4870
rect 27371 4378 27427 4380
rect 27451 4378 27507 4380
rect 27531 4378 27587 4380
rect 27611 4378 27667 4380
rect 27371 4326 27417 4378
rect 27417 4326 27427 4378
rect 27451 4326 27481 4378
rect 27481 4326 27493 4378
rect 27493 4326 27507 4378
rect 27531 4326 27545 4378
rect 27545 4326 27557 4378
rect 27557 4326 27587 4378
rect 27611 4326 27621 4378
rect 27621 4326 27667 4378
rect 27371 4324 27427 4326
rect 27451 4324 27507 4326
rect 27531 4324 27587 4326
rect 27611 4324 27667 4326
rect 23518 3834 23574 3836
rect 23598 3834 23654 3836
rect 23678 3834 23734 3836
rect 23758 3834 23814 3836
rect 23518 3782 23564 3834
rect 23564 3782 23574 3834
rect 23598 3782 23628 3834
rect 23628 3782 23640 3834
rect 23640 3782 23654 3834
rect 23678 3782 23692 3834
rect 23692 3782 23704 3834
rect 23704 3782 23734 3834
rect 23758 3782 23768 3834
rect 23768 3782 23814 3834
rect 23518 3780 23574 3782
rect 23598 3780 23654 3782
rect 23678 3780 23734 3782
rect 23758 3780 23814 3782
rect 31223 3834 31279 3836
rect 31303 3834 31359 3836
rect 31383 3834 31439 3836
rect 31463 3834 31519 3836
rect 31223 3782 31269 3834
rect 31269 3782 31279 3834
rect 31303 3782 31333 3834
rect 31333 3782 31345 3834
rect 31345 3782 31359 3834
rect 31383 3782 31397 3834
rect 31397 3782 31409 3834
rect 31409 3782 31439 3834
rect 31463 3782 31473 3834
rect 31473 3782 31519 3834
rect 31223 3780 31279 3782
rect 31303 3780 31359 3782
rect 31383 3780 31439 3782
rect 31463 3780 31519 3782
rect 27371 3290 27427 3292
rect 27451 3290 27507 3292
rect 27531 3290 27587 3292
rect 27611 3290 27667 3292
rect 27371 3238 27417 3290
rect 27417 3238 27427 3290
rect 27451 3238 27481 3290
rect 27481 3238 27493 3290
rect 27493 3238 27507 3290
rect 27531 3238 27545 3290
rect 27545 3238 27557 3290
rect 27557 3238 27587 3290
rect 27611 3238 27621 3290
rect 27621 3238 27667 3290
rect 27371 3236 27427 3238
rect 27451 3236 27507 3238
rect 27531 3236 27587 3238
rect 27611 3236 27667 3238
rect 23518 2746 23574 2748
rect 23598 2746 23654 2748
rect 23678 2746 23734 2748
rect 23758 2746 23814 2748
rect 23518 2694 23564 2746
rect 23564 2694 23574 2746
rect 23598 2694 23628 2746
rect 23628 2694 23640 2746
rect 23640 2694 23654 2746
rect 23678 2694 23692 2746
rect 23692 2694 23704 2746
rect 23704 2694 23734 2746
rect 23758 2694 23768 2746
rect 23768 2694 23814 2746
rect 23518 2692 23574 2694
rect 23598 2692 23654 2694
rect 23678 2692 23734 2694
rect 23758 2692 23814 2694
rect 31223 2746 31279 2748
rect 31303 2746 31359 2748
rect 31383 2746 31439 2748
rect 31463 2746 31519 2748
rect 31223 2694 31269 2746
rect 31269 2694 31279 2746
rect 31303 2694 31333 2746
rect 31333 2694 31345 2746
rect 31345 2694 31359 2746
rect 31383 2694 31397 2746
rect 31397 2694 31409 2746
rect 31409 2694 31439 2746
rect 31463 2694 31473 2746
rect 31473 2694 31519 2746
rect 31223 2692 31279 2694
rect 31303 2692 31359 2694
rect 31383 2692 31439 2694
rect 31463 2692 31519 2694
rect 27371 2202 27427 2204
rect 27451 2202 27507 2204
rect 27531 2202 27587 2204
rect 27611 2202 27667 2204
rect 27371 2150 27417 2202
rect 27417 2150 27427 2202
rect 27451 2150 27481 2202
rect 27481 2150 27493 2202
rect 27493 2150 27507 2202
rect 27531 2150 27545 2202
rect 27545 2150 27557 2202
rect 27557 2150 27587 2202
rect 27611 2150 27621 2202
rect 27621 2150 27667 2202
rect 27371 2148 27427 2150
rect 27451 2148 27507 2150
rect 27531 2148 27587 2150
rect 27611 2148 27667 2150
rect 23518 1658 23574 1660
rect 23598 1658 23654 1660
rect 23678 1658 23734 1660
rect 23758 1658 23814 1660
rect 23518 1606 23564 1658
rect 23564 1606 23574 1658
rect 23598 1606 23628 1658
rect 23628 1606 23640 1658
rect 23640 1606 23654 1658
rect 23678 1606 23692 1658
rect 23692 1606 23704 1658
rect 23704 1606 23734 1658
rect 23758 1606 23768 1658
rect 23768 1606 23814 1658
rect 23518 1604 23574 1606
rect 23598 1604 23654 1606
rect 23678 1604 23734 1606
rect 23758 1604 23814 1606
rect 31223 1658 31279 1660
rect 31303 1658 31359 1660
rect 31383 1658 31439 1660
rect 31463 1658 31519 1660
rect 31223 1606 31269 1658
rect 31269 1606 31279 1658
rect 31303 1606 31333 1658
rect 31333 1606 31345 1658
rect 31345 1606 31359 1658
rect 31383 1606 31397 1658
rect 31397 1606 31409 1658
rect 31409 1606 31439 1658
rect 31463 1606 31473 1658
rect 31473 1606 31519 1658
rect 31223 1604 31279 1606
rect 31303 1604 31359 1606
rect 31383 1604 31439 1606
rect 31463 1604 31519 1606
rect 27371 1114 27427 1116
rect 27451 1114 27507 1116
rect 27531 1114 27587 1116
rect 27611 1114 27667 1116
rect 27371 1062 27417 1114
rect 27417 1062 27427 1114
rect 27451 1062 27481 1114
rect 27481 1062 27493 1114
rect 27493 1062 27507 1114
rect 27531 1062 27545 1114
rect 27545 1062 27557 1114
rect 27557 1062 27587 1114
rect 27611 1062 27621 1114
rect 27621 1062 27667 1114
rect 27371 1060 27427 1062
rect 27451 1060 27507 1062
rect 27531 1060 27587 1062
rect 27611 1060 27667 1062
rect 23518 570 23574 572
rect 23598 570 23654 572
rect 23678 570 23734 572
rect 23758 570 23814 572
rect 23518 518 23564 570
rect 23564 518 23574 570
rect 23598 518 23628 570
rect 23628 518 23640 570
rect 23640 518 23654 570
rect 23678 518 23692 570
rect 23692 518 23704 570
rect 23704 518 23734 570
rect 23758 518 23768 570
rect 23768 518 23814 570
rect 23518 516 23574 518
rect 23598 516 23654 518
rect 23678 516 23734 518
rect 23758 516 23814 518
rect 31223 570 31279 572
rect 31303 570 31359 572
rect 31383 570 31439 572
rect 31463 570 31519 572
rect 31223 518 31269 570
rect 31269 518 31279 570
rect 31303 518 31333 570
rect 31333 518 31345 570
rect 31345 518 31359 570
rect 31383 518 31397 570
rect 31397 518 31409 570
rect 31409 518 31439 570
rect 31463 518 31473 570
rect 31473 518 31519 570
rect 31223 516 31279 518
rect 31303 516 31359 518
rect 31383 516 31439 518
rect 31463 516 31519 518
<< metal3 >>
rect 8098 19072 8414 19073
rect 8098 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8414 19072
rect 8098 19007 8414 19008
rect 15803 19072 16119 19073
rect 15803 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16119 19072
rect 15803 19007 16119 19008
rect 23508 19072 23824 19073
rect 23508 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23824 19072
rect 23508 19007 23824 19008
rect 31213 19072 31529 19073
rect 31213 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31529 19072
rect 31213 19007 31529 19008
rect 4246 18528 4562 18529
rect 4246 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4562 18528
rect 4246 18463 4562 18464
rect 11951 18528 12267 18529
rect 11951 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12267 18528
rect 11951 18463 12267 18464
rect 19656 18528 19972 18529
rect 19656 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19972 18528
rect 19656 18463 19972 18464
rect 27361 18528 27677 18529
rect 27361 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27677 18528
rect 27361 18463 27677 18464
rect 8098 17984 8414 17985
rect 8098 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8414 17984
rect 8098 17919 8414 17920
rect 15803 17984 16119 17985
rect 15803 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16119 17984
rect 15803 17919 16119 17920
rect 23508 17984 23824 17985
rect 23508 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23824 17984
rect 23508 17919 23824 17920
rect 31213 17984 31529 17985
rect 31213 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31529 17984
rect 31213 17919 31529 17920
rect 4246 17440 4562 17441
rect 4246 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4562 17440
rect 4246 17375 4562 17376
rect 11951 17440 12267 17441
rect 11951 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12267 17440
rect 11951 17375 12267 17376
rect 19656 17440 19972 17441
rect 19656 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19972 17440
rect 19656 17375 19972 17376
rect 27361 17440 27677 17441
rect 27361 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27677 17440
rect 27361 17375 27677 17376
rect 8098 16896 8414 16897
rect 8098 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8414 16896
rect 8098 16831 8414 16832
rect 15803 16896 16119 16897
rect 15803 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16119 16896
rect 15803 16831 16119 16832
rect 23508 16896 23824 16897
rect 23508 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23824 16896
rect 23508 16831 23824 16832
rect 31213 16896 31529 16897
rect 31213 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31529 16896
rect 31213 16831 31529 16832
rect 4246 16352 4562 16353
rect 4246 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4562 16352
rect 4246 16287 4562 16288
rect 11951 16352 12267 16353
rect 11951 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12267 16352
rect 11951 16287 12267 16288
rect 19656 16352 19972 16353
rect 19656 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19972 16352
rect 19656 16287 19972 16288
rect 27361 16352 27677 16353
rect 27361 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27677 16352
rect 27361 16287 27677 16288
rect 8098 15808 8414 15809
rect 8098 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8414 15808
rect 8098 15743 8414 15744
rect 15803 15808 16119 15809
rect 15803 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16119 15808
rect 15803 15743 16119 15744
rect 23508 15808 23824 15809
rect 23508 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23824 15808
rect 23508 15743 23824 15744
rect 31213 15808 31529 15809
rect 31213 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31529 15808
rect 31213 15743 31529 15744
rect 4246 15264 4562 15265
rect 4246 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4562 15264
rect 4246 15199 4562 15200
rect 11951 15264 12267 15265
rect 11951 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12267 15264
rect 11951 15199 12267 15200
rect 19656 15264 19972 15265
rect 19656 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19972 15264
rect 19656 15199 19972 15200
rect 27361 15264 27677 15265
rect 27361 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27677 15264
rect 27361 15199 27677 15200
rect 8098 14720 8414 14721
rect 8098 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8414 14720
rect 8098 14655 8414 14656
rect 15803 14720 16119 14721
rect 15803 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16119 14720
rect 15803 14655 16119 14656
rect 23508 14720 23824 14721
rect 23508 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23824 14720
rect 23508 14655 23824 14656
rect 31213 14720 31529 14721
rect 31213 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31529 14720
rect 31213 14655 31529 14656
rect 4246 14176 4562 14177
rect 4246 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4562 14176
rect 4246 14111 4562 14112
rect 11951 14176 12267 14177
rect 11951 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12267 14176
rect 11951 14111 12267 14112
rect 19656 14176 19972 14177
rect 19656 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19972 14176
rect 19656 14111 19972 14112
rect 27361 14176 27677 14177
rect 27361 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27677 14176
rect 27361 14111 27677 14112
rect 8098 13632 8414 13633
rect 8098 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8414 13632
rect 8098 13567 8414 13568
rect 15803 13632 16119 13633
rect 15803 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16119 13632
rect 15803 13567 16119 13568
rect 23508 13632 23824 13633
rect 23508 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23824 13632
rect 23508 13567 23824 13568
rect 31213 13632 31529 13633
rect 31213 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31529 13632
rect 31213 13567 31529 13568
rect 4246 13088 4562 13089
rect 4246 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4562 13088
rect 4246 13023 4562 13024
rect 11951 13088 12267 13089
rect 11951 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12267 13088
rect 11951 13023 12267 13024
rect 19656 13088 19972 13089
rect 19656 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19972 13088
rect 19656 13023 19972 13024
rect 27361 13088 27677 13089
rect 27361 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27677 13088
rect 27361 13023 27677 13024
rect 8098 12544 8414 12545
rect 8098 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8414 12544
rect 8098 12479 8414 12480
rect 15803 12544 16119 12545
rect 15803 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16119 12544
rect 15803 12479 16119 12480
rect 23508 12544 23824 12545
rect 23508 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23824 12544
rect 23508 12479 23824 12480
rect 31213 12544 31529 12545
rect 31213 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31529 12544
rect 31213 12479 31529 12480
rect 4246 12000 4562 12001
rect 4246 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4562 12000
rect 4246 11935 4562 11936
rect 11951 12000 12267 12001
rect 11951 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12267 12000
rect 11951 11935 12267 11936
rect 19656 12000 19972 12001
rect 19656 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19972 12000
rect 19656 11935 19972 11936
rect 27361 12000 27677 12001
rect 27361 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27677 12000
rect 27361 11935 27677 11936
rect 8098 11456 8414 11457
rect 8098 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8414 11456
rect 8098 11391 8414 11392
rect 15803 11456 16119 11457
rect 15803 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16119 11456
rect 15803 11391 16119 11392
rect 23508 11456 23824 11457
rect 23508 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23824 11456
rect 23508 11391 23824 11392
rect 31213 11456 31529 11457
rect 31213 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31529 11456
rect 31213 11391 31529 11392
rect 4246 10912 4562 10913
rect 4246 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4562 10912
rect 4246 10847 4562 10848
rect 11951 10912 12267 10913
rect 11951 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12267 10912
rect 11951 10847 12267 10848
rect 19656 10912 19972 10913
rect 19656 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19972 10912
rect 19656 10847 19972 10848
rect 27361 10912 27677 10913
rect 27361 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27677 10912
rect 27361 10847 27677 10848
rect 8098 10368 8414 10369
rect 0 10298 400 10328
rect 8098 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8414 10368
rect 8098 10303 8414 10304
rect 15803 10368 16119 10369
rect 15803 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16119 10368
rect 15803 10303 16119 10304
rect 23508 10368 23824 10369
rect 23508 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23824 10368
rect 23508 10303 23824 10304
rect 31213 10368 31529 10369
rect 31213 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31529 10368
rect 31213 10303 31529 10304
rect 11881 10298 11947 10301
rect 0 10238 2790 10298
rect 0 10208 400 10238
rect 2730 10162 2790 10238
rect 8526 10296 11947 10298
rect 8526 10240 11886 10296
rect 11942 10240 11947 10296
rect 8526 10238 11947 10240
rect 8526 10162 8586 10238
rect 11881 10235 11947 10238
rect 31600 10296 32000 10328
rect 31600 10240 31666 10296
rect 31722 10240 32000 10296
rect 31600 10208 32000 10240
rect 2730 10102 8586 10162
rect 4246 9824 4562 9825
rect 4246 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4562 9824
rect 4246 9759 4562 9760
rect 11951 9824 12267 9825
rect 11951 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12267 9824
rect 11951 9759 12267 9760
rect 19656 9824 19972 9825
rect 19656 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19972 9824
rect 19656 9759 19972 9760
rect 27361 9824 27677 9825
rect 27361 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27677 9824
rect 27361 9759 27677 9760
rect 9581 9756 9647 9757
rect 15561 9756 15627 9757
rect 9581 9752 9628 9756
rect 9692 9754 9698 9756
rect 15510 9754 15516 9756
rect 9581 9696 9586 9752
rect 9581 9692 9628 9696
rect 9692 9694 9738 9754
rect 15470 9694 15516 9754
rect 15580 9752 15627 9756
rect 15622 9696 15627 9752
rect 9692 9692 9698 9694
rect 15510 9692 15516 9694
rect 15580 9692 15627 9696
rect 9581 9691 9647 9692
rect 15561 9691 15627 9692
rect 0 9618 400 9648
rect 10133 9618 10199 9621
rect 0 9616 10199 9618
rect 0 9560 10138 9616
rect 10194 9560 10199 9616
rect 0 9558 10199 9560
rect 0 9528 400 9558
rect 10133 9555 10199 9558
rect 28257 9618 28323 9621
rect 31600 9618 32000 9648
rect 28257 9616 32000 9618
rect 28257 9560 28262 9616
rect 28318 9560 32000 9616
rect 28257 9558 32000 9560
rect 28257 9555 28323 9558
rect 31600 9528 32000 9558
rect 8098 9280 8414 9281
rect 8098 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8414 9280
rect 8098 9215 8414 9216
rect 15803 9280 16119 9281
rect 15803 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16119 9280
rect 15803 9215 16119 9216
rect 23508 9280 23824 9281
rect 23508 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23824 9280
rect 23508 9215 23824 9216
rect 31213 9280 31529 9281
rect 31213 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31529 9280
rect 31213 9215 31529 9216
rect 8201 9074 8267 9077
rect 11789 9074 11855 9077
rect 8201 9072 11855 9074
rect 8201 9016 8206 9072
rect 8262 9016 11794 9072
rect 11850 9016 11855 9072
rect 8201 9014 11855 9016
rect 8201 9011 8267 9014
rect 11789 9011 11855 9014
rect 0 8938 400 8968
rect 11145 8938 11211 8941
rect 0 8936 11211 8938
rect 0 8880 11150 8936
rect 11206 8880 11211 8936
rect 0 8878 11211 8880
rect 0 8848 400 8878
rect 11145 8875 11211 8878
rect 28257 8938 28323 8941
rect 31600 8938 32000 8968
rect 28257 8936 32000 8938
rect 28257 8880 28262 8936
rect 28318 8880 32000 8936
rect 28257 8878 32000 8880
rect 28257 8875 28323 8878
rect 31600 8848 32000 8878
rect 4246 8736 4562 8737
rect 4246 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4562 8736
rect 4246 8671 4562 8672
rect 11951 8736 12267 8737
rect 11951 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12267 8736
rect 11951 8671 12267 8672
rect 19656 8736 19972 8737
rect 19656 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19972 8736
rect 19656 8671 19972 8672
rect 27361 8736 27677 8737
rect 27361 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27677 8736
rect 27361 8671 27677 8672
rect 9397 8530 9463 8533
rect 9397 8528 12450 8530
rect 9397 8472 9402 8528
rect 9458 8472 12450 8528
rect 9397 8470 12450 8472
rect 9397 8467 9463 8470
rect 11145 8394 11211 8397
rect 12157 8394 12223 8397
rect 11145 8392 12223 8394
rect 11145 8336 11150 8392
rect 11206 8336 12162 8392
rect 12218 8336 12223 8392
rect 11145 8334 12223 8336
rect 12390 8394 12450 8470
rect 12566 8394 12572 8396
rect 12390 8334 12572 8394
rect 11145 8331 11211 8334
rect 12157 8331 12223 8334
rect 12566 8332 12572 8334
rect 12636 8332 12642 8396
rect 0 8258 400 8288
rect 10961 8258 11027 8261
rect 13077 8258 13143 8261
rect 0 8198 2790 8258
rect 0 8168 400 8198
rect 2730 7986 2790 8198
rect 10961 8256 13143 8258
rect 10961 8200 10966 8256
rect 11022 8200 13082 8256
rect 13138 8200 13143 8256
rect 10961 8198 13143 8200
rect 10961 8195 11027 8198
rect 13077 8195 13143 8198
rect 8098 8192 8414 8193
rect 8098 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8414 8192
rect 8098 8127 8414 8128
rect 15803 8192 16119 8193
rect 15803 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16119 8192
rect 15803 8127 16119 8128
rect 23508 8192 23824 8193
rect 23508 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23824 8192
rect 23508 8127 23824 8128
rect 31213 8192 31529 8193
rect 31213 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31529 8192
rect 31213 8127 31529 8128
rect 11145 8122 11211 8125
rect 8526 8120 11211 8122
rect 8526 8064 11150 8120
rect 11206 8064 11211 8120
rect 8526 8062 11211 8064
rect 8526 7986 8586 8062
rect 11145 8059 11211 8062
rect 11973 8122 12039 8125
rect 14089 8122 14155 8125
rect 11973 8120 14155 8122
rect 11973 8064 11978 8120
rect 12034 8064 14094 8120
rect 14150 8064 14155 8120
rect 11973 8062 14155 8064
rect 11973 8059 12039 8062
rect 14089 8059 14155 8062
rect 2730 7926 8586 7986
rect 11605 7986 11671 7989
rect 12985 7986 13051 7989
rect 11605 7984 13051 7986
rect 11605 7928 11610 7984
rect 11666 7928 12990 7984
rect 13046 7928 13051 7984
rect 11605 7926 13051 7928
rect 11605 7923 11671 7926
rect 12985 7923 13051 7926
rect 12157 7850 12223 7853
rect 12893 7850 12959 7853
rect 12157 7848 12959 7850
rect 12157 7792 12162 7848
rect 12218 7792 12898 7848
rect 12954 7792 12959 7848
rect 12157 7790 12959 7792
rect 12157 7787 12223 7790
rect 12893 7787 12959 7790
rect 4246 7648 4562 7649
rect 4246 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4562 7648
rect 4246 7583 4562 7584
rect 11951 7648 12267 7649
rect 11951 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12267 7648
rect 11951 7583 12267 7584
rect 19656 7648 19972 7649
rect 19656 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19972 7648
rect 19656 7583 19972 7584
rect 27361 7648 27677 7649
rect 27361 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27677 7648
rect 27361 7583 27677 7584
rect 10133 7170 10199 7173
rect 10593 7170 10659 7173
rect 10133 7168 10659 7170
rect 10133 7112 10138 7168
rect 10194 7112 10598 7168
rect 10654 7112 10659 7168
rect 10133 7110 10659 7112
rect 10133 7107 10199 7110
rect 10593 7107 10659 7110
rect 8098 7104 8414 7105
rect 8098 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8414 7104
rect 8098 7039 8414 7040
rect 15803 7104 16119 7105
rect 15803 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16119 7104
rect 15803 7039 16119 7040
rect 23508 7104 23824 7105
rect 23508 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23824 7104
rect 23508 7039 23824 7040
rect 31213 7104 31529 7105
rect 31213 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31529 7104
rect 31213 7039 31529 7040
rect 10961 7034 11027 7037
rect 11697 7034 11763 7037
rect 10961 7032 11763 7034
rect 10961 6976 10966 7032
rect 11022 6976 11702 7032
rect 11758 6976 11763 7032
rect 10961 6974 11763 6976
rect 10961 6971 11027 6974
rect 11697 6971 11763 6974
rect 9622 6836 9628 6900
rect 9692 6898 9698 6900
rect 11881 6898 11947 6901
rect 9692 6896 11947 6898
rect 9692 6840 11886 6896
rect 11942 6840 11947 6896
rect 9692 6838 11947 6840
rect 9692 6836 9698 6838
rect 11881 6835 11947 6838
rect 12566 6836 12572 6900
rect 12636 6898 12642 6900
rect 12801 6898 12867 6901
rect 12636 6896 12867 6898
rect 12636 6840 12806 6896
rect 12862 6840 12867 6896
rect 12636 6838 12867 6840
rect 12636 6836 12642 6838
rect 12801 6835 12867 6838
rect 10041 6762 10107 6765
rect 12157 6762 12223 6765
rect 10041 6760 12223 6762
rect 10041 6704 10046 6760
rect 10102 6704 12162 6760
rect 12218 6704 12223 6760
rect 10041 6702 12223 6704
rect 10041 6699 10107 6702
rect 12157 6699 12223 6702
rect 9673 6626 9739 6629
rect 11513 6626 11579 6629
rect 11697 6626 11763 6629
rect 9673 6624 11763 6626
rect 9673 6568 9678 6624
rect 9734 6568 11518 6624
rect 11574 6568 11702 6624
rect 11758 6568 11763 6624
rect 9673 6566 11763 6568
rect 9673 6563 9739 6566
rect 11513 6563 11579 6566
rect 11697 6563 11763 6566
rect 4246 6560 4562 6561
rect 4246 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4562 6560
rect 4246 6495 4562 6496
rect 11951 6560 12267 6561
rect 11951 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12267 6560
rect 11951 6495 12267 6496
rect 19656 6560 19972 6561
rect 19656 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19972 6560
rect 19656 6495 19972 6496
rect 27361 6560 27677 6561
rect 27361 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27677 6560
rect 27361 6495 27677 6496
rect 10225 6490 10291 6493
rect 11697 6490 11763 6493
rect 10225 6488 11763 6490
rect 10225 6432 10230 6488
rect 10286 6432 11702 6488
rect 11758 6432 11763 6488
rect 10225 6430 11763 6432
rect 10225 6427 10291 6430
rect 11697 6427 11763 6430
rect 9857 6354 9923 6357
rect 10869 6354 10935 6357
rect 9857 6352 10935 6354
rect 9857 6296 9862 6352
rect 9918 6296 10874 6352
rect 10930 6296 10935 6352
rect 9857 6294 10935 6296
rect 9857 6291 9923 6294
rect 10869 6291 10935 6294
rect 8098 6016 8414 6017
rect 8098 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8414 6016
rect 8098 5951 8414 5952
rect 15803 6016 16119 6017
rect 15803 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16119 6016
rect 15803 5951 16119 5952
rect 23508 6016 23824 6017
rect 23508 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23824 6016
rect 23508 5951 23824 5952
rect 31213 6016 31529 6017
rect 31213 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31529 6016
rect 31213 5951 31529 5952
rect 4246 5472 4562 5473
rect 4246 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4562 5472
rect 4246 5407 4562 5408
rect 11951 5472 12267 5473
rect 11951 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12267 5472
rect 11951 5407 12267 5408
rect 19656 5472 19972 5473
rect 19656 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19972 5472
rect 19656 5407 19972 5408
rect 27361 5472 27677 5473
rect 27361 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27677 5472
rect 27361 5407 27677 5408
rect 8098 4928 8414 4929
rect 8098 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8414 4928
rect 8098 4863 8414 4864
rect 15803 4928 16119 4929
rect 15803 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16119 4928
rect 15803 4863 16119 4864
rect 23508 4928 23824 4929
rect 23508 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23824 4928
rect 23508 4863 23824 4864
rect 31213 4928 31529 4929
rect 31213 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31529 4928
rect 31213 4863 31529 4864
rect 4246 4384 4562 4385
rect 4246 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4562 4384
rect 4246 4319 4562 4320
rect 11951 4384 12267 4385
rect 11951 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12267 4384
rect 11951 4319 12267 4320
rect 19656 4384 19972 4385
rect 19656 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19972 4384
rect 19656 4319 19972 4320
rect 27361 4384 27677 4385
rect 27361 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27677 4384
rect 27361 4319 27677 4320
rect 15469 4044 15535 4045
rect 15469 4042 15516 4044
rect 15424 4040 15516 4042
rect 15424 3984 15474 4040
rect 15424 3982 15516 3984
rect 15469 3980 15516 3982
rect 15580 3980 15586 4044
rect 15469 3979 15535 3980
rect 8098 3840 8414 3841
rect 8098 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8414 3840
rect 8098 3775 8414 3776
rect 15803 3840 16119 3841
rect 15803 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16119 3840
rect 15803 3775 16119 3776
rect 23508 3840 23824 3841
rect 23508 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23824 3840
rect 23508 3775 23824 3776
rect 31213 3840 31529 3841
rect 31213 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31529 3840
rect 31213 3775 31529 3776
rect 4246 3296 4562 3297
rect 4246 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4562 3296
rect 4246 3231 4562 3232
rect 11951 3296 12267 3297
rect 11951 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12267 3296
rect 11951 3231 12267 3232
rect 19656 3296 19972 3297
rect 19656 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19972 3296
rect 19656 3231 19972 3232
rect 27361 3296 27677 3297
rect 27361 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27677 3296
rect 27361 3231 27677 3232
rect 8098 2752 8414 2753
rect 8098 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8414 2752
rect 8098 2687 8414 2688
rect 15803 2752 16119 2753
rect 15803 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16119 2752
rect 15803 2687 16119 2688
rect 23508 2752 23824 2753
rect 23508 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23824 2752
rect 23508 2687 23824 2688
rect 31213 2752 31529 2753
rect 31213 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31529 2752
rect 31213 2687 31529 2688
rect 4246 2208 4562 2209
rect 4246 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4562 2208
rect 4246 2143 4562 2144
rect 11951 2208 12267 2209
rect 11951 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12267 2208
rect 11951 2143 12267 2144
rect 19656 2208 19972 2209
rect 19656 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19972 2208
rect 19656 2143 19972 2144
rect 27361 2208 27677 2209
rect 27361 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27677 2208
rect 27361 2143 27677 2144
rect 8098 1664 8414 1665
rect 8098 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8414 1664
rect 8098 1599 8414 1600
rect 15803 1664 16119 1665
rect 15803 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16119 1664
rect 15803 1599 16119 1600
rect 23508 1664 23824 1665
rect 23508 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23824 1664
rect 23508 1599 23824 1600
rect 31213 1664 31529 1665
rect 31213 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31529 1664
rect 31213 1599 31529 1600
rect 4246 1120 4562 1121
rect 4246 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4562 1120
rect 4246 1055 4562 1056
rect 11951 1120 12267 1121
rect 11951 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12267 1120
rect 11951 1055 12267 1056
rect 19656 1120 19972 1121
rect 19656 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19972 1120
rect 19656 1055 19972 1056
rect 27361 1120 27677 1121
rect 27361 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27677 1120
rect 27361 1055 27677 1056
rect 8098 576 8414 577
rect 8098 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8414 576
rect 8098 511 8414 512
rect 15803 576 16119 577
rect 15803 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16119 576
rect 15803 511 16119 512
rect 23508 576 23824 577
rect 23508 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23824 576
rect 23508 511 23824 512
rect 31213 576 31529 577
rect 31213 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31529 576
rect 31213 511 31529 512
<< via3 >>
rect 8104 19068 8168 19072
rect 8104 19012 8108 19068
rect 8108 19012 8164 19068
rect 8164 19012 8168 19068
rect 8104 19008 8168 19012
rect 8184 19068 8248 19072
rect 8184 19012 8188 19068
rect 8188 19012 8244 19068
rect 8244 19012 8248 19068
rect 8184 19008 8248 19012
rect 8264 19068 8328 19072
rect 8264 19012 8268 19068
rect 8268 19012 8324 19068
rect 8324 19012 8328 19068
rect 8264 19008 8328 19012
rect 8344 19068 8408 19072
rect 8344 19012 8348 19068
rect 8348 19012 8404 19068
rect 8404 19012 8408 19068
rect 8344 19008 8408 19012
rect 15809 19068 15873 19072
rect 15809 19012 15813 19068
rect 15813 19012 15869 19068
rect 15869 19012 15873 19068
rect 15809 19008 15873 19012
rect 15889 19068 15953 19072
rect 15889 19012 15893 19068
rect 15893 19012 15949 19068
rect 15949 19012 15953 19068
rect 15889 19008 15953 19012
rect 15969 19068 16033 19072
rect 15969 19012 15973 19068
rect 15973 19012 16029 19068
rect 16029 19012 16033 19068
rect 15969 19008 16033 19012
rect 16049 19068 16113 19072
rect 16049 19012 16053 19068
rect 16053 19012 16109 19068
rect 16109 19012 16113 19068
rect 16049 19008 16113 19012
rect 23514 19068 23578 19072
rect 23514 19012 23518 19068
rect 23518 19012 23574 19068
rect 23574 19012 23578 19068
rect 23514 19008 23578 19012
rect 23594 19068 23658 19072
rect 23594 19012 23598 19068
rect 23598 19012 23654 19068
rect 23654 19012 23658 19068
rect 23594 19008 23658 19012
rect 23674 19068 23738 19072
rect 23674 19012 23678 19068
rect 23678 19012 23734 19068
rect 23734 19012 23738 19068
rect 23674 19008 23738 19012
rect 23754 19068 23818 19072
rect 23754 19012 23758 19068
rect 23758 19012 23814 19068
rect 23814 19012 23818 19068
rect 23754 19008 23818 19012
rect 31219 19068 31283 19072
rect 31219 19012 31223 19068
rect 31223 19012 31279 19068
rect 31279 19012 31283 19068
rect 31219 19008 31283 19012
rect 31299 19068 31363 19072
rect 31299 19012 31303 19068
rect 31303 19012 31359 19068
rect 31359 19012 31363 19068
rect 31299 19008 31363 19012
rect 31379 19068 31443 19072
rect 31379 19012 31383 19068
rect 31383 19012 31439 19068
rect 31439 19012 31443 19068
rect 31379 19008 31443 19012
rect 31459 19068 31523 19072
rect 31459 19012 31463 19068
rect 31463 19012 31519 19068
rect 31519 19012 31523 19068
rect 31459 19008 31523 19012
rect 4252 18524 4316 18528
rect 4252 18468 4256 18524
rect 4256 18468 4312 18524
rect 4312 18468 4316 18524
rect 4252 18464 4316 18468
rect 4332 18524 4396 18528
rect 4332 18468 4336 18524
rect 4336 18468 4392 18524
rect 4392 18468 4396 18524
rect 4332 18464 4396 18468
rect 4412 18524 4476 18528
rect 4412 18468 4416 18524
rect 4416 18468 4472 18524
rect 4472 18468 4476 18524
rect 4412 18464 4476 18468
rect 4492 18524 4556 18528
rect 4492 18468 4496 18524
rect 4496 18468 4552 18524
rect 4552 18468 4556 18524
rect 4492 18464 4556 18468
rect 11957 18524 12021 18528
rect 11957 18468 11961 18524
rect 11961 18468 12017 18524
rect 12017 18468 12021 18524
rect 11957 18464 12021 18468
rect 12037 18524 12101 18528
rect 12037 18468 12041 18524
rect 12041 18468 12097 18524
rect 12097 18468 12101 18524
rect 12037 18464 12101 18468
rect 12117 18524 12181 18528
rect 12117 18468 12121 18524
rect 12121 18468 12177 18524
rect 12177 18468 12181 18524
rect 12117 18464 12181 18468
rect 12197 18524 12261 18528
rect 12197 18468 12201 18524
rect 12201 18468 12257 18524
rect 12257 18468 12261 18524
rect 12197 18464 12261 18468
rect 19662 18524 19726 18528
rect 19662 18468 19666 18524
rect 19666 18468 19722 18524
rect 19722 18468 19726 18524
rect 19662 18464 19726 18468
rect 19742 18524 19806 18528
rect 19742 18468 19746 18524
rect 19746 18468 19802 18524
rect 19802 18468 19806 18524
rect 19742 18464 19806 18468
rect 19822 18524 19886 18528
rect 19822 18468 19826 18524
rect 19826 18468 19882 18524
rect 19882 18468 19886 18524
rect 19822 18464 19886 18468
rect 19902 18524 19966 18528
rect 19902 18468 19906 18524
rect 19906 18468 19962 18524
rect 19962 18468 19966 18524
rect 19902 18464 19966 18468
rect 27367 18524 27431 18528
rect 27367 18468 27371 18524
rect 27371 18468 27427 18524
rect 27427 18468 27431 18524
rect 27367 18464 27431 18468
rect 27447 18524 27511 18528
rect 27447 18468 27451 18524
rect 27451 18468 27507 18524
rect 27507 18468 27511 18524
rect 27447 18464 27511 18468
rect 27527 18524 27591 18528
rect 27527 18468 27531 18524
rect 27531 18468 27587 18524
rect 27587 18468 27591 18524
rect 27527 18464 27591 18468
rect 27607 18524 27671 18528
rect 27607 18468 27611 18524
rect 27611 18468 27667 18524
rect 27667 18468 27671 18524
rect 27607 18464 27671 18468
rect 8104 17980 8168 17984
rect 8104 17924 8108 17980
rect 8108 17924 8164 17980
rect 8164 17924 8168 17980
rect 8104 17920 8168 17924
rect 8184 17980 8248 17984
rect 8184 17924 8188 17980
rect 8188 17924 8244 17980
rect 8244 17924 8248 17980
rect 8184 17920 8248 17924
rect 8264 17980 8328 17984
rect 8264 17924 8268 17980
rect 8268 17924 8324 17980
rect 8324 17924 8328 17980
rect 8264 17920 8328 17924
rect 8344 17980 8408 17984
rect 8344 17924 8348 17980
rect 8348 17924 8404 17980
rect 8404 17924 8408 17980
rect 8344 17920 8408 17924
rect 15809 17980 15873 17984
rect 15809 17924 15813 17980
rect 15813 17924 15869 17980
rect 15869 17924 15873 17980
rect 15809 17920 15873 17924
rect 15889 17980 15953 17984
rect 15889 17924 15893 17980
rect 15893 17924 15949 17980
rect 15949 17924 15953 17980
rect 15889 17920 15953 17924
rect 15969 17980 16033 17984
rect 15969 17924 15973 17980
rect 15973 17924 16029 17980
rect 16029 17924 16033 17980
rect 15969 17920 16033 17924
rect 16049 17980 16113 17984
rect 16049 17924 16053 17980
rect 16053 17924 16109 17980
rect 16109 17924 16113 17980
rect 16049 17920 16113 17924
rect 23514 17980 23578 17984
rect 23514 17924 23518 17980
rect 23518 17924 23574 17980
rect 23574 17924 23578 17980
rect 23514 17920 23578 17924
rect 23594 17980 23658 17984
rect 23594 17924 23598 17980
rect 23598 17924 23654 17980
rect 23654 17924 23658 17980
rect 23594 17920 23658 17924
rect 23674 17980 23738 17984
rect 23674 17924 23678 17980
rect 23678 17924 23734 17980
rect 23734 17924 23738 17980
rect 23674 17920 23738 17924
rect 23754 17980 23818 17984
rect 23754 17924 23758 17980
rect 23758 17924 23814 17980
rect 23814 17924 23818 17980
rect 23754 17920 23818 17924
rect 31219 17980 31283 17984
rect 31219 17924 31223 17980
rect 31223 17924 31279 17980
rect 31279 17924 31283 17980
rect 31219 17920 31283 17924
rect 31299 17980 31363 17984
rect 31299 17924 31303 17980
rect 31303 17924 31359 17980
rect 31359 17924 31363 17980
rect 31299 17920 31363 17924
rect 31379 17980 31443 17984
rect 31379 17924 31383 17980
rect 31383 17924 31439 17980
rect 31439 17924 31443 17980
rect 31379 17920 31443 17924
rect 31459 17980 31523 17984
rect 31459 17924 31463 17980
rect 31463 17924 31519 17980
rect 31519 17924 31523 17980
rect 31459 17920 31523 17924
rect 4252 17436 4316 17440
rect 4252 17380 4256 17436
rect 4256 17380 4312 17436
rect 4312 17380 4316 17436
rect 4252 17376 4316 17380
rect 4332 17436 4396 17440
rect 4332 17380 4336 17436
rect 4336 17380 4392 17436
rect 4392 17380 4396 17436
rect 4332 17376 4396 17380
rect 4412 17436 4476 17440
rect 4412 17380 4416 17436
rect 4416 17380 4472 17436
rect 4472 17380 4476 17436
rect 4412 17376 4476 17380
rect 4492 17436 4556 17440
rect 4492 17380 4496 17436
rect 4496 17380 4552 17436
rect 4552 17380 4556 17436
rect 4492 17376 4556 17380
rect 11957 17436 12021 17440
rect 11957 17380 11961 17436
rect 11961 17380 12017 17436
rect 12017 17380 12021 17436
rect 11957 17376 12021 17380
rect 12037 17436 12101 17440
rect 12037 17380 12041 17436
rect 12041 17380 12097 17436
rect 12097 17380 12101 17436
rect 12037 17376 12101 17380
rect 12117 17436 12181 17440
rect 12117 17380 12121 17436
rect 12121 17380 12177 17436
rect 12177 17380 12181 17436
rect 12117 17376 12181 17380
rect 12197 17436 12261 17440
rect 12197 17380 12201 17436
rect 12201 17380 12257 17436
rect 12257 17380 12261 17436
rect 12197 17376 12261 17380
rect 19662 17436 19726 17440
rect 19662 17380 19666 17436
rect 19666 17380 19722 17436
rect 19722 17380 19726 17436
rect 19662 17376 19726 17380
rect 19742 17436 19806 17440
rect 19742 17380 19746 17436
rect 19746 17380 19802 17436
rect 19802 17380 19806 17436
rect 19742 17376 19806 17380
rect 19822 17436 19886 17440
rect 19822 17380 19826 17436
rect 19826 17380 19882 17436
rect 19882 17380 19886 17436
rect 19822 17376 19886 17380
rect 19902 17436 19966 17440
rect 19902 17380 19906 17436
rect 19906 17380 19962 17436
rect 19962 17380 19966 17436
rect 19902 17376 19966 17380
rect 27367 17436 27431 17440
rect 27367 17380 27371 17436
rect 27371 17380 27427 17436
rect 27427 17380 27431 17436
rect 27367 17376 27431 17380
rect 27447 17436 27511 17440
rect 27447 17380 27451 17436
rect 27451 17380 27507 17436
rect 27507 17380 27511 17436
rect 27447 17376 27511 17380
rect 27527 17436 27591 17440
rect 27527 17380 27531 17436
rect 27531 17380 27587 17436
rect 27587 17380 27591 17436
rect 27527 17376 27591 17380
rect 27607 17436 27671 17440
rect 27607 17380 27611 17436
rect 27611 17380 27667 17436
rect 27667 17380 27671 17436
rect 27607 17376 27671 17380
rect 8104 16892 8168 16896
rect 8104 16836 8108 16892
rect 8108 16836 8164 16892
rect 8164 16836 8168 16892
rect 8104 16832 8168 16836
rect 8184 16892 8248 16896
rect 8184 16836 8188 16892
rect 8188 16836 8244 16892
rect 8244 16836 8248 16892
rect 8184 16832 8248 16836
rect 8264 16892 8328 16896
rect 8264 16836 8268 16892
rect 8268 16836 8324 16892
rect 8324 16836 8328 16892
rect 8264 16832 8328 16836
rect 8344 16892 8408 16896
rect 8344 16836 8348 16892
rect 8348 16836 8404 16892
rect 8404 16836 8408 16892
rect 8344 16832 8408 16836
rect 15809 16892 15873 16896
rect 15809 16836 15813 16892
rect 15813 16836 15869 16892
rect 15869 16836 15873 16892
rect 15809 16832 15873 16836
rect 15889 16892 15953 16896
rect 15889 16836 15893 16892
rect 15893 16836 15949 16892
rect 15949 16836 15953 16892
rect 15889 16832 15953 16836
rect 15969 16892 16033 16896
rect 15969 16836 15973 16892
rect 15973 16836 16029 16892
rect 16029 16836 16033 16892
rect 15969 16832 16033 16836
rect 16049 16892 16113 16896
rect 16049 16836 16053 16892
rect 16053 16836 16109 16892
rect 16109 16836 16113 16892
rect 16049 16832 16113 16836
rect 23514 16892 23578 16896
rect 23514 16836 23518 16892
rect 23518 16836 23574 16892
rect 23574 16836 23578 16892
rect 23514 16832 23578 16836
rect 23594 16892 23658 16896
rect 23594 16836 23598 16892
rect 23598 16836 23654 16892
rect 23654 16836 23658 16892
rect 23594 16832 23658 16836
rect 23674 16892 23738 16896
rect 23674 16836 23678 16892
rect 23678 16836 23734 16892
rect 23734 16836 23738 16892
rect 23674 16832 23738 16836
rect 23754 16892 23818 16896
rect 23754 16836 23758 16892
rect 23758 16836 23814 16892
rect 23814 16836 23818 16892
rect 23754 16832 23818 16836
rect 31219 16892 31283 16896
rect 31219 16836 31223 16892
rect 31223 16836 31279 16892
rect 31279 16836 31283 16892
rect 31219 16832 31283 16836
rect 31299 16892 31363 16896
rect 31299 16836 31303 16892
rect 31303 16836 31359 16892
rect 31359 16836 31363 16892
rect 31299 16832 31363 16836
rect 31379 16892 31443 16896
rect 31379 16836 31383 16892
rect 31383 16836 31439 16892
rect 31439 16836 31443 16892
rect 31379 16832 31443 16836
rect 31459 16892 31523 16896
rect 31459 16836 31463 16892
rect 31463 16836 31519 16892
rect 31519 16836 31523 16892
rect 31459 16832 31523 16836
rect 4252 16348 4316 16352
rect 4252 16292 4256 16348
rect 4256 16292 4312 16348
rect 4312 16292 4316 16348
rect 4252 16288 4316 16292
rect 4332 16348 4396 16352
rect 4332 16292 4336 16348
rect 4336 16292 4392 16348
rect 4392 16292 4396 16348
rect 4332 16288 4396 16292
rect 4412 16348 4476 16352
rect 4412 16292 4416 16348
rect 4416 16292 4472 16348
rect 4472 16292 4476 16348
rect 4412 16288 4476 16292
rect 4492 16348 4556 16352
rect 4492 16292 4496 16348
rect 4496 16292 4552 16348
rect 4552 16292 4556 16348
rect 4492 16288 4556 16292
rect 11957 16348 12021 16352
rect 11957 16292 11961 16348
rect 11961 16292 12017 16348
rect 12017 16292 12021 16348
rect 11957 16288 12021 16292
rect 12037 16348 12101 16352
rect 12037 16292 12041 16348
rect 12041 16292 12097 16348
rect 12097 16292 12101 16348
rect 12037 16288 12101 16292
rect 12117 16348 12181 16352
rect 12117 16292 12121 16348
rect 12121 16292 12177 16348
rect 12177 16292 12181 16348
rect 12117 16288 12181 16292
rect 12197 16348 12261 16352
rect 12197 16292 12201 16348
rect 12201 16292 12257 16348
rect 12257 16292 12261 16348
rect 12197 16288 12261 16292
rect 19662 16348 19726 16352
rect 19662 16292 19666 16348
rect 19666 16292 19722 16348
rect 19722 16292 19726 16348
rect 19662 16288 19726 16292
rect 19742 16348 19806 16352
rect 19742 16292 19746 16348
rect 19746 16292 19802 16348
rect 19802 16292 19806 16348
rect 19742 16288 19806 16292
rect 19822 16348 19886 16352
rect 19822 16292 19826 16348
rect 19826 16292 19882 16348
rect 19882 16292 19886 16348
rect 19822 16288 19886 16292
rect 19902 16348 19966 16352
rect 19902 16292 19906 16348
rect 19906 16292 19962 16348
rect 19962 16292 19966 16348
rect 19902 16288 19966 16292
rect 27367 16348 27431 16352
rect 27367 16292 27371 16348
rect 27371 16292 27427 16348
rect 27427 16292 27431 16348
rect 27367 16288 27431 16292
rect 27447 16348 27511 16352
rect 27447 16292 27451 16348
rect 27451 16292 27507 16348
rect 27507 16292 27511 16348
rect 27447 16288 27511 16292
rect 27527 16348 27591 16352
rect 27527 16292 27531 16348
rect 27531 16292 27587 16348
rect 27587 16292 27591 16348
rect 27527 16288 27591 16292
rect 27607 16348 27671 16352
rect 27607 16292 27611 16348
rect 27611 16292 27667 16348
rect 27667 16292 27671 16348
rect 27607 16288 27671 16292
rect 8104 15804 8168 15808
rect 8104 15748 8108 15804
rect 8108 15748 8164 15804
rect 8164 15748 8168 15804
rect 8104 15744 8168 15748
rect 8184 15804 8248 15808
rect 8184 15748 8188 15804
rect 8188 15748 8244 15804
rect 8244 15748 8248 15804
rect 8184 15744 8248 15748
rect 8264 15804 8328 15808
rect 8264 15748 8268 15804
rect 8268 15748 8324 15804
rect 8324 15748 8328 15804
rect 8264 15744 8328 15748
rect 8344 15804 8408 15808
rect 8344 15748 8348 15804
rect 8348 15748 8404 15804
rect 8404 15748 8408 15804
rect 8344 15744 8408 15748
rect 15809 15804 15873 15808
rect 15809 15748 15813 15804
rect 15813 15748 15869 15804
rect 15869 15748 15873 15804
rect 15809 15744 15873 15748
rect 15889 15804 15953 15808
rect 15889 15748 15893 15804
rect 15893 15748 15949 15804
rect 15949 15748 15953 15804
rect 15889 15744 15953 15748
rect 15969 15804 16033 15808
rect 15969 15748 15973 15804
rect 15973 15748 16029 15804
rect 16029 15748 16033 15804
rect 15969 15744 16033 15748
rect 16049 15804 16113 15808
rect 16049 15748 16053 15804
rect 16053 15748 16109 15804
rect 16109 15748 16113 15804
rect 16049 15744 16113 15748
rect 23514 15804 23578 15808
rect 23514 15748 23518 15804
rect 23518 15748 23574 15804
rect 23574 15748 23578 15804
rect 23514 15744 23578 15748
rect 23594 15804 23658 15808
rect 23594 15748 23598 15804
rect 23598 15748 23654 15804
rect 23654 15748 23658 15804
rect 23594 15744 23658 15748
rect 23674 15804 23738 15808
rect 23674 15748 23678 15804
rect 23678 15748 23734 15804
rect 23734 15748 23738 15804
rect 23674 15744 23738 15748
rect 23754 15804 23818 15808
rect 23754 15748 23758 15804
rect 23758 15748 23814 15804
rect 23814 15748 23818 15804
rect 23754 15744 23818 15748
rect 31219 15804 31283 15808
rect 31219 15748 31223 15804
rect 31223 15748 31279 15804
rect 31279 15748 31283 15804
rect 31219 15744 31283 15748
rect 31299 15804 31363 15808
rect 31299 15748 31303 15804
rect 31303 15748 31359 15804
rect 31359 15748 31363 15804
rect 31299 15744 31363 15748
rect 31379 15804 31443 15808
rect 31379 15748 31383 15804
rect 31383 15748 31439 15804
rect 31439 15748 31443 15804
rect 31379 15744 31443 15748
rect 31459 15804 31523 15808
rect 31459 15748 31463 15804
rect 31463 15748 31519 15804
rect 31519 15748 31523 15804
rect 31459 15744 31523 15748
rect 4252 15260 4316 15264
rect 4252 15204 4256 15260
rect 4256 15204 4312 15260
rect 4312 15204 4316 15260
rect 4252 15200 4316 15204
rect 4332 15260 4396 15264
rect 4332 15204 4336 15260
rect 4336 15204 4392 15260
rect 4392 15204 4396 15260
rect 4332 15200 4396 15204
rect 4412 15260 4476 15264
rect 4412 15204 4416 15260
rect 4416 15204 4472 15260
rect 4472 15204 4476 15260
rect 4412 15200 4476 15204
rect 4492 15260 4556 15264
rect 4492 15204 4496 15260
rect 4496 15204 4552 15260
rect 4552 15204 4556 15260
rect 4492 15200 4556 15204
rect 11957 15260 12021 15264
rect 11957 15204 11961 15260
rect 11961 15204 12017 15260
rect 12017 15204 12021 15260
rect 11957 15200 12021 15204
rect 12037 15260 12101 15264
rect 12037 15204 12041 15260
rect 12041 15204 12097 15260
rect 12097 15204 12101 15260
rect 12037 15200 12101 15204
rect 12117 15260 12181 15264
rect 12117 15204 12121 15260
rect 12121 15204 12177 15260
rect 12177 15204 12181 15260
rect 12117 15200 12181 15204
rect 12197 15260 12261 15264
rect 12197 15204 12201 15260
rect 12201 15204 12257 15260
rect 12257 15204 12261 15260
rect 12197 15200 12261 15204
rect 19662 15260 19726 15264
rect 19662 15204 19666 15260
rect 19666 15204 19722 15260
rect 19722 15204 19726 15260
rect 19662 15200 19726 15204
rect 19742 15260 19806 15264
rect 19742 15204 19746 15260
rect 19746 15204 19802 15260
rect 19802 15204 19806 15260
rect 19742 15200 19806 15204
rect 19822 15260 19886 15264
rect 19822 15204 19826 15260
rect 19826 15204 19882 15260
rect 19882 15204 19886 15260
rect 19822 15200 19886 15204
rect 19902 15260 19966 15264
rect 19902 15204 19906 15260
rect 19906 15204 19962 15260
rect 19962 15204 19966 15260
rect 19902 15200 19966 15204
rect 27367 15260 27431 15264
rect 27367 15204 27371 15260
rect 27371 15204 27427 15260
rect 27427 15204 27431 15260
rect 27367 15200 27431 15204
rect 27447 15260 27511 15264
rect 27447 15204 27451 15260
rect 27451 15204 27507 15260
rect 27507 15204 27511 15260
rect 27447 15200 27511 15204
rect 27527 15260 27591 15264
rect 27527 15204 27531 15260
rect 27531 15204 27587 15260
rect 27587 15204 27591 15260
rect 27527 15200 27591 15204
rect 27607 15260 27671 15264
rect 27607 15204 27611 15260
rect 27611 15204 27667 15260
rect 27667 15204 27671 15260
rect 27607 15200 27671 15204
rect 8104 14716 8168 14720
rect 8104 14660 8108 14716
rect 8108 14660 8164 14716
rect 8164 14660 8168 14716
rect 8104 14656 8168 14660
rect 8184 14716 8248 14720
rect 8184 14660 8188 14716
rect 8188 14660 8244 14716
rect 8244 14660 8248 14716
rect 8184 14656 8248 14660
rect 8264 14716 8328 14720
rect 8264 14660 8268 14716
rect 8268 14660 8324 14716
rect 8324 14660 8328 14716
rect 8264 14656 8328 14660
rect 8344 14716 8408 14720
rect 8344 14660 8348 14716
rect 8348 14660 8404 14716
rect 8404 14660 8408 14716
rect 8344 14656 8408 14660
rect 15809 14716 15873 14720
rect 15809 14660 15813 14716
rect 15813 14660 15869 14716
rect 15869 14660 15873 14716
rect 15809 14656 15873 14660
rect 15889 14716 15953 14720
rect 15889 14660 15893 14716
rect 15893 14660 15949 14716
rect 15949 14660 15953 14716
rect 15889 14656 15953 14660
rect 15969 14716 16033 14720
rect 15969 14660 15973 14716
rect 15973 14660 16029 14716
rect 16029 14660 16033 14716
rect 15969 14656 16033 14660
rect 16049 14716 16113 14720
rect 16049 14660 16053 14716
rect 16053 14660 16109 14716
rect 16109 14660 16113 14716
rect 16049 14656 16113 14660
rect 23514 14716 23578 14720
rect 23514 14660 23518 14716
rect 23518 14660 23574 14716
rect 23574 14660 23578 14716
rect 23514 14656 23578 14660
rect 23594 14716 23658 14720
rect 23594 14660 23598 14716
rect 23598 14660 23654 14716
rect 23654 14660 23658 14716
rect 23594 14656 23658 14660
rect 23674 14716 23738 14720
rect 23674 14660 23678 14716
rect 23678 14660 23734 14716
rect 23734 14660 23738 14716
rect 23674 14656 23738 14660
rect 23754 14716 23818 14720
rect 23754 14660 23758 14716
rect 23758 14660 23814 14716
rect 23814 14660 23818 14716
rect 23754 14656 23818 14660
rect 31219 14716 31283 14720
rect 31219 14660 31223 14716
rect 31223 14660 31279 14716
rect 31279 14660 31283 14716
rect 31219 14656 31283 14660
rect 31299 14716 31363 14720
rect 31299 14660 31303 14716
rect 31303 14660 31359 14716
rect 31359 14660 31363 14716
rect 31299 14656 31363 14660
rect 31379 14716 31443 14720
rect 31379 14660 31383 14716
rect 31383 14660 31439 14716
rect 31439 14660 31443 14716
rect 31379 14656 31443 14660
rect 31459 14716 31523 14720
rect 31459 14660 31463 14716
rect 31463 14660 31519 14716
rect 31519 14660 31523 14716
rect 31459 14656 31523 14660
rect 4252 14172 4316 14176
rect 4252 14116 4256 14172
rect 4256 14116 4312 14172
rect 4312 14116 4316 14172
rect 4252 14112 4316 14116
rect 4332 14172 4396 14176
rect 4332 14116 4336 14172
rect 4336 14116 4392 14172
rect 4392 14116 4396 14172
rect 4332 14112 4396 14116
rect 4412 14172 4476 14176
rect 4412 14116 4416 14172
rect 4416 14116 4472 14172
rect 4472 14116 4476 14172
rect 4412 14112 4476 14116
rect 4492 14172 4556 14176
rect 4492 14116 4496 14172
rect 4496 14116 4552 14172
rect 4552 14116 4556 14172
rect 4492 14112 4556 14116
rect 11957 14172 12021 14176
rect 11957 14116 11961 14172
rect 11961 14116 12017 14172
rect 12017 14116 12021 14172
rect 11957 14112 12021 14116
rect 12037 14172 12101 14176
rect 12037 14116 12041 14172
rect 12041 14116 12097 14172
rect 12097 14116 12101 14172
rect 12037 14112 12101 14116
rect 12117 14172 12181 14176
rect 12117 14116 12121 14172
rect 12121 14116 12177 14172
rect 12177 14116 12181 14172
rect 12117 14112 12181 14116
rect 12197 14172 12261 14176
rect 12197 14116 12201 14172
rect 12201 14116 12257 14172
rect 12257 14116 12261 14172
rect 12197 14112 12261 14116
rect 19662 14172 19726 14176
rect 19662 14116 19666 14172
rect 19666 14116 19722 14172
rect 19722 14116 19726 14172
rect 19662 14112 19726 14116
rect 19742 14172 19806 14176
rect 19742 14116 19746 14172
rect 19746 14116 19802 14172
rect 19802 14116 19806 14172
rect 19742 14112 19806 14116
rect 19822 14172 19886 14176
rect 19822 14116 19826 14172
rect 19826 14116 19882 14172
rect 19882 14116 19886 14172
rect 19822 14112 19886 14116
rect 19902 14172 19966 14176
rect 19902 14116 19906 14172
rect 19906 14116 19962 14172
rect 19962 14116 19966 14172
rect 19902 14112 19966 14116
rect 27367 14172 27431 14176
rect 27367 14116 27371 14172
rect 27371 14116 27427 14172
rect 27427 14116 27431 14172
rect 27367 14112 27431 14116
rect 27447 14172 27511 14176
rect 27447 14116 27451 14172
rect 27451 14116 27507 14172
rect 27507 14116 27511 14172
rect 27447 14112 27511 14116
rect 27527 14172 27591 14176
rect 27527 14116 27531 14172
rect 27531 14116 27587 14172
rect 27587 14116 27591 14172
rect 27527 14112 27591 14116
rect 27607 14172 27671 14176
rect 27607 14116 27611 14172
rect 27611 14116 27667 14172
rect 27667 14116 27671 14172
rect 27607 14112 27671 14116
rect 8104 13628 8168 13632
rect 8104 13572 8108 13628
rect 8108 13572 8164 13628
rect 8164 13572 8168 13628
rect 8104 13568 8168 13572
rect 8184 13628 8248 13632
rect 8184 13572 8188 13628
rect 8188 13572 8244 13628
rect 8244 13572 8248 13628
rect 8184 13568 8248 13572
rect 8264 13628 8328 13632
rect 8264 13572 8268 13628
rect 8268 13572 8324 13628
rect 8324 13572 8328 13628
rect 8264 13568 8328 13572
rect 8344 13628 8408 13632
rect 8344 13572 8348 13628
rect 8348 13572 8404 13628
rect 8404 13572 8408 13628
rect 8344 13568 8408 13572
rect 15809 13628 15873 13632
rect 15809 13572 15813 13628
rect 15813 13572 15869 13628
rect 15869 13572 15873 13628
rect 15809 13568 15873 13572
rect 15889 13628 15953 13632
rect 15889 13572 15893 13628
rect 15893 13572 15949 13628
rect 15949 13572 15953 13628
rect 15889 13568 15953 13572
rect 15969 13628 16033 13632
rect 15969 13572 15973 13628
rect 15973 13572 16029 13628
rect 16029 13572 16033 13628
rect 15969 13568 16033 13572
rect 16049 13628 16113 13632
rect 16049 13572 16053 13628
rect 16053 13572 16109 13628
rect 16109 13572 16113 13628
rect 16049 13568 16113 13572
rect 23514 13628 23578 13632
rect 23514 13572 23518 13628
rect 23518 13572 23574 13628
rect 23574 13572 23578 13628
rect 23514 13568 23578 13572
rect 23594 13628 23658 13632
rect 23594 13572 23598 13628
rect 23598 13572 23654 13628
rect 23654 13572 23658 13628
rect 23594 13568 23658 13572
rect 23674 13628 23738 13632
rect 23674 13572 23678 13628
rect 23678 13572 23734 13628
rect 23734 13572 23738 13628
rect 23674 13568 23738 13572
rect 23754 13628 23818 13632
rect 23754 13572 23758 13628
rect 23758 13572 23814 13628
rect 23814 13572 23818 13628
rect 23754 13568 23818 13572
rect 31219 13628 31283 13632
rect 31219 13572 31223 13628
rect 31223 13572 31279 13628
rect 31279 13572 31283 13628
rect 31219 13568 31283 13572
rect 31299 13628 31363 13632
rect 31299 13572 31303 13628
rect 31303 13572 31359 13628
rect 31359 13572 31363 13628
rect 31299 13568 31363 13572
rect 31379 13628 31443 13632
rect 31379 13572 31383 13628
rect 31383 13572 31439 13628
rect 31439 13572 31443 13628
rect 31379 13568 31443 13572
rect 31459 13628 31523 13632
rect 31459 13572 31463 13628
rect 31463 13572 31519 13628
rect 31519 13572 31523 13628
rect 31459 13568 31523 13572
rect 4252 13084 4316 13088
rect 4252 13028 4256 13084
rect 4256 13028 4312 13084
rect 4312 13028 4316 13084
rect 4252 13024 4316 13028
rect 4332 13084 4396 13088
rect 4332 13028 4336 13084
rect 4336 13028 4392 13084
rect 4392 13028 4396 13084
rect 4332 13024 4396 13028
rect 4412 13084 4476 13088
rect 4412 13028 4416 13084
rect 4416 13028 4472 13084
rect 4472 13028 4476 13084
rect 4412 13024 4476 13028
rect 4492 13084 4556 13088
rect 4492 13028 4496 13084
rect 4496 13028 4552 13084
rect 4552 13028 4556 13084
rect 4492 13024 4556 13028
rect 11957 13084 12021 13088
rect 11957 13028 11961 13084
rect 11961 13028 12017 13084
rect 12017 13028 12021 13084
rect 11957 13024 12021 13028
rect 12037 13084 12101 13088
rect 12037 13028 12041 13084
rect 12041 13028 12097 13084
rect 12097 13028 12101 13084
rect 12037 13024 12101 13028
rect 12117 13084 12181 13088
rect 12117 13028 12121 13084
rect 12121 13028 12177 13084
rect 12177 13028 12181 13084
rect 12117 13024 12181 13028
rect 12197 13084 12261 13088
rect 12197 13028 12201 13084
rect 12201 13028 12257 13084
rect 12257 13028 12261 13084
rect 12197 13024 12261 13028
rect 19662 13084 19726 13088
rect 19662 13028 19666 13084
rect 19666 13028 19722 13084
rect 19722 13028 19726 13084
rect 19662 13024 19726 13028
rect 19742 13084 19806 13088
rect 19742 13028 19746 13084
rect 19746 13028 19802 13084
rect 19802 13028 19806 13084
rect 19742 13024 19806 13028
rect 19822 13084 19886 13088
rect 19822 13028 19826 13084
rect 19826 13028 19882 13084
rect 19882 13028 19886 13084
rect 19822 13024 19886 13028
rect 19902 13084 19966 13088
rect 19902 13028 19906 13084
rect 19906 13028 19962 13084
rect 19962 13028 19966 13084
rect 19902 13024 19966 13028
rect 27367 13084 27431 13088
rect 27367 13028 27371 13084
rect 27371 13028 27427 13084
rect 27427 13028 27431 13084
rect 27367 13024 27431 13028
rect 27447 13084 27511 13088
rect 27447 13028 27451 13084
rect 27451 13028 27507 13084
rect 27507 13028 27511 13084
rect 27447 13024 27511 13028
rect 27527 13084 27591 13088
rect 27527 13028 27531 13084
rect 27531 13028 27587 13084
rect 27587 13028 27591 13084
rect 27527 13024 27591 13028
rect 27607 13084 27671 13088
rect 27607 13028 27611 13084
rect 27611 13028 27667 13084
rect 27667 13028 27671 13084
rect 27607 13024 27671 13028
rect 8104 12540 8168 12544
rect 8104 12484 8108 12540
rect 8108 12484 8164 12540
rect 8164 12484 8168 12540
rect 8104 12480 8168 12484
rect 8184 12540 8248 12544
rect 8184 12484 8188 12540
rect 8188 12484 8244 12540
rect 8244 12484 8248 12540
rect 8184 12480 8248 12484
rect 8264 12540 8328 12544
rect 8264 12484 8268 12540
rect 8268 12484 8324 12540
rect 8324 12484 8328 12540
rect 8264 12480 8328 12484
rect 8344 12540 8408 12544
rect 8344 12484 8348 12540
rect 8348 12484 8404 12540
rect 8404 12484 8408 12540
rect 8344 12480 8408 12484
rect 15809 12540 15873 12544
rect 15809 12484 15813 12540
rect 15813 12484 15869 12540
rect 15869 12484 15873 12540
rect 15809 12480 15873 12484
rect 15889 12540 15953 12544
rect 15889 12484 15893 12540
rect 15893 12484 15949 12540
rect 15949 12484 15953 12540
rect 15889 12480 15953 12484
rect 15969 12540 16033 12544
rect 15969 12484 15973 12540
rect 15973 12484 16029 12540
rect 16029 12484 16033 12540
rect 15969 12480 16033 12484
rect 16049 12540 16113 12544
rect 16049 12484 16053 12540
rect 16053 12484 16109 12540
rect 16109 12484 16113 12540
rect 16049 12480 16113 12484
rect 23514 12540 23578 12544
rect 23514 12484 23518 12540
rect 23518 12484 23574 12540
rect 23574 12484 23578 12540
rect 23514 12480 23578 12484
rect 23594 12540 23658 12544
rect 23594 12484 23598 12540
rect 23598 12484 23654 12540
rect 23654 12484 23658 12540
rect 23594 12480 23658 12484
rect 23674 12540 23738 12544
rect 23674 12484 23678 12540
rect 23678 12484 23734 12540
rect 23734 12484 23738 12540
rect 23674 12480 23738 12484
rect 23754 12540 23818 12544
rect 23754 12484 23758 12540
rect 23758 12484 23814 12540
rect 23814 12484 23818 12540
rect 23754 12480 23818 12484
rect 31219 12540 31283 12544
rect 31219 12484 31223 12540
rect 31223 12484 31279 12540
rect 31279 12484 31283 12540
rect 31219 12480 31283 12484
rect 31299 12540 31363 12544
rect 31299 12484 31303 12540
rect 31303 12484 31359 12540
rect 31359 12484 31363 12540
rect 31299 12480 31363 12484
rect 31379 12540 31443 12544
rect 31379 12484 31383 12540
rect 31383 12484 31439 12540
rect 31439 12484 31443 12540
rect 31379 12480 31443 12484
rect 31459 12540 31523 12544
rect 31459 12484 31463 12540
rect 31463 12484 31519 12540
rect 31519 12484 31523 12540
rect 31459 12480 31523 12484
rect 4252 11996 4316 12000
rect 4252 11940 4256 11996
rect 4256 11940 4312 11996
rect 4312 11940 4316 11996
rect 4252 11936 4316 11940
rect 4332 11996 4396 12000
rect 4332 11940 4336 11996
rect 4336 11940 4392 11996
rect 4392 11940 4396 11996
rect 4332 11936 4396 11940
rect 4412 11996 4476 12000
rect 4412 11940 4416 11996
rect 4416 11940 4472 11996
rect 4472 11940 4476 11996
rect 4412 11936 4476 11940
rect 4492 11996 4556 12000
rect 4492 11940 4496 11996
rect 4496 11940 4552 11996
rect 4552 11940 4556 11996
rect 4492 11936 4556 11940
rect 11957 11996 12021 12000
rect 11957 11940 11961 11996
rect 11961 11940 12017 11996
rect 12017 11940 12021 11996
rect 11957 11936 12021 11940
rect 12037 11996 12101 12000
rect 12037 11940 12041 11996
rect 12041 11940 12097 11996
rect 12097 11940 12101 11996
rect 12037 11936 12101 11940
rect 12117 11996 12181 12000
rect 12117 11940 12121 11996
rect 12121 11940 12177 11996
rect 12177 11940 12181 11996
rect 12117 11936 12181 11940
rect 12197 11996 12261 12000
rect 12197 11940 12201 11996
rect 12201 11940 12257 11996
rect 12257 11940 12261 11996
rect 12197 11936 12261 11940
rect 19662 11996 19726 12000
rect 19662 11940 19666 11996
rect 19666 11940 19722 11996
rect 19722 11940 19726 11996
rect 19662 11936 19726 11940
rect 19742 11996 19806 12000
rect 19742 11940 19746 11996
rect 19746 11940 19802 11996
rect 19802 11940 19806 11996
rect 19742 11936 19806 11940
rect 19822 11996 19886 12000
rect 19822 11940 19826 11996
rect 19826 11940 19882 11996
rect 19882 11940 19886 11996
rect 19822 11936 19886 11940
rect 19902 11996 19966 12000
rect 19902 11940 19906 11996
rect 19906 11940 19962 11996
rect 19962 11940 19966 11996
rect 19902 11936 19966 11940
rect 27367 11996 27431 12000
rect 27367 11940 27371 11996
rect 27371 11940 27427 11996
rect 27427 11940 27431 11996
rect 27367 11936 27431 11940
rect 27447 11996 27511 12000
rect 27447 11940 27451 11996
rect 27451 11940 27507 11996
rect 27507 11940 27511 11996
rect 27447 11936 27511 11940
rect 27527 11996 27591 12000
rect 27527 11940 27531 11996
rect 27531 11940 27587 11996
rect 27587 11940 27591 11996
rect 27527 11936 27591 11940
rect 27607 11996 27671 12000
rect 27607 11940 27611 11996
rect 27611 11940 27667 11996
rect 27667 11940 27671 11996
rect 27607 11936 27671 11940
rect 8104 11452 8168 11456
rect 8104 11396 8108 11452
rect 8108 11396 8164 11452
rect 8164 11396 8168 11452
rect 8104 11392 8168 11396
rect 8184 11452 8248 11456
rect 8184 11396 8188 11452
rect 8188 11396 8244 11452
rect 8244 11396 8248 11452
rect 8184 11392 8248 11396
rect 8264 11452 8328 11456
rect 8264 11396 8268 11452
rect 8268 11396 8324 11452
rect 8324 11396 8328 11452
rect 8264 11392 8328 11396
rect 8344 11452 8408 11456
rect 8344 11396 8348 11452
rect 8348 11396 8404 11452
rect 8404 11396 8408 11452
rect 8344 11392 8408 11396
rect 15809 11452 15873 11456
rect 15809 11396 15813 11452
rect 15813 11396 15869 11452
rect 15869 11396 15873 11452
rect 15809 11392 15873 11396
rect 15889 11452 15953 11456
rect 15889 11396 15893 11452
rect 15893 11396 15949 11452
rect 15949 11396 15953 11452
rect 15889 11392 15953 11396
rect 15969 11452 16033 11456
rect 15969 11396 15973 11452
rect 15973 11396 16029 11452
rect 16029 11396 16033 11452
rect 15969 11392 16033 11396
rect 16049 11452 16113 11456
rect 16049 11396 16053 11452
rect 16053 11396 16109 11452
rect 16109 11396 16113 11452
rect 16049 11392 16113 11396
rect 23514 11452 23578 11456
rect 23514 11396 23518 11452
rect 23518 11396 23574 11452
rect 23574 11396 23578 11452
rect 23514 11392 23578 11396
rect 23594 11452 23658 11456
rect 23594 11396 23598 11452
rect 23598 11396 23654 11452
rect 23654 11396 23658 11452
rect 23594 11392 23658 11396
rect 23674 11452 23738 11456
rect 23674 11396 23678 11452
rect 23678 11396 23734 11452
rect 23734 11396 23738 11452
rect 23674 11392 23738 11396
rect 23754 11452 23818 11456
rect 23754 11396 23758 11452
rect 23758 11396 23814 11452
rect 23814 11396 23818 11452
rect 23754 11392 23818 11396
rect 31219 11452 31283 11456
rect 31219 11396 31223 11452
rect 31223 11396 31279 11452
rect 31279 11396 31283 11452
rect 31219 11392 31283 11396
rect 31299 11452 31363 11456
rect 31299 11396 31303 11452
rect 31303 11396 31359 11452
rect 31359 11396 31363 11452
rect 31299 11392 31363 11396
rect 31379 11452 31443 11456
rect 31379 11396 31383 11452
rect 31383 11396 31439 11452
rect 31439 11396 31443 11452
rect 31379 11392 31443 11396
rect 31459 11452 31523 11456
rect 31459 11396 31463 11452
rect 31463 11396 31519 11452
rect 31519 11396 31523 11452
rect 31459 11392 31523 11396
rect 4252 10908 4316 10912
rect 4252 10852 4256 10908
rect 4256 10852 4312 10908
rect 4312 10852 4316 10908
rect 4252 10848 4316 10852
rect 4332 10908 4396 10912
rect 4332 10852 4336 10908
rect 4336 10852 4392 10908
rect 4392 10852 4396 10908
rect 4332 10848 4396 10852
rect 4412 10908 4476 10912
rect 4412 10852 4416 10908
rect 4416 10852 4472 10908
rect 4472 10852 4476 10908
rect 4412 10848 4476 10852
rect 4492 10908 4556 10912
rect 4492 10852 4496 10908
rect 4496 10852 4552 10908
rect 4552 10852 4556 10908
rect 4492 10848 4556 10852
rect 11957 10908 12021 10912
rect 11957 10852 11961 10908
rect 11961 10852 12017 10908
rect 12017 10852 12021 10908
rect 11957 10848 12021 10852
rect 12037 10908 12101 10912
rect 12037 10852 12041 10908
rect 12041 10852 12097 10908
rect 12097 10852 12101 10908
rect 12037 10848 12101 10852
rect 12117 10908 12181 10912
rect 12117 10852 12121 10908
rect 12121 10852 12177 10908
rect 12177 10852 12181 10908
rect 12117 10848 12181 10852
rect 12197 10908 12261 10912
rect 12197 10852 12201 10908
rect 12201 10852 12257 10908
rect 12257 10852 12261 10908
rect 12197 10848 12261 10852
rect 19662 10908 19726 10912
rect 19662 10852 19666 10908
rect 19666 10852 19722 10908
rect 19722 10852 19726 10908
rect 19662 10848 19726 10852
rect 19742 10908 19806 10912
rect 19742 10852 19746 10908
rect 19746 10852 19802 10908
rect 19802 10852 19806 10908
rect 19742 10848 19806 10852
rect 19822 10908 19886 10912
rect 19822 10852 19826 10908
rect 19826 10852 19882 10908
rect 19882 10852 19886 10908
rect 19822 10848 19886 10852
rect 19902 10908 19966 10912
rect 19902 10852 19906 10908
rect 19906 10852 19962 10908
rect 19962 10852 19966 10908
rect 19902 10848 19966 10852
rect 27367 10908 27431 10912
rect 27367 10852 27371 10908
rect 27371 10852 27427 10908
rect 27427 10852 27431 10908
rect 27367 10848 27431 10852
rect 27447 10908 27511 10912
rect 27447 10852 27451 10908
rect 27451 10852 27507 10908
rect 27507 10852 27511 10908
rect 27447 10848 27511 10852
rect 27527 10908 27591 10912
rect 27527 10852 27531 10908
rect 27531 10852 27587 10908
rect 27587 10852 27591 10908
rect 27527 10848 27591 10852
rect 27607 10908 27671 10912
rect 27607 10852 27611 10908
rect 27611 10852 27667 10908
rect 27667 10852 27671 10908
rect 27607 10848 27671 10852
rect 8104 10364 8168 10368
rect 8104 10308 8108 10364
rect 8108 10308 8164 10364
rect 8164 10308 8168 10364
rect 8104 10304 8168 10308
rect 8184 10364 8248 10368
rect 8184 10308 8188 10364
rect 8188 10308 8244 10364
rect 8244 10308 8248 10364
rect 8184 10304 8248 10308
rect 8264 10364 8328 10368
rect 8264 10308 8268 10364
rect 8268 10308 8324 10364
rect 8324 10308 8328 10364
rect 8264 10304 8328 10308
rect 8344 10364 8408 10368
rect 8344 10308 8348 10364
rect 8348 10308 8404 10364
rect 8404 10308 8408 10364
rect 8344 10304 8408 10308
rect 15809 10364 15873 10368
rect 15809 10308 15813 10364
rect 15813 10308 15869 10364
rect 15869 10308 15873 10364
rect 15809 10304 15873 10308
rect 15889 10364 15953 10368
rect 15889 10308 15893 10364
rect 15893 10308 15949 10364
rect 15949 10308 15953 10364
rect 15889 10304 15953 10308
rect 15969 10364 16033 10368
rect 15969 10308 15973 10364
rect 15973 10308 16029 10364
rect 16029 10308 16033 10364
rect 15969 10304 16033 10308
rect 16049 10364 16113 10368
rect 16049 10308 16053 10364
rect 16053 10308 16109 10364
rect 16109 10308 16113 10364
rect 16049 10304 16113 10308
rect 23514 10364 23578 10368
rect 23514 10308 23518 10364
rect 23518 10308 23574 10364
rect 23574 10308 23578 10364
rect 23514 10304 23578 10308
rect 23594 10364 23658 10368
rect 23594 10308 23598 10364
rect 23598 10308 23654 10364
rect 23654 10308 23658 10364
rect 23594 10304 23658 10308
rect 23674 10364 23738 10368
rect 23674 10308 23678 10364
rect 23678 10308 23734 10364
rect 23734 10308 23738 10364
rect 23674 10304 23738 10308
rect 23754 10364 23818 10368
rect 23754 10308 23758 10364
rect 23758 10308 23814 10364
rect 23814 10308 23818 10364
rect 23754 10304 23818 10308
rect 31219 10364 31283 10368
rect 31219 10308 31223 10364
rect 31223 10308 31279 10364
rect 31279 10308 31283 10364
rect 31219 10304 31283 10308
rect 31299 10364 31363 10368
rect 31299 10308 31303 10364
rect 31303 10308 31359 10364
rect 31359 10308 31363 10364
rect 31299 10304 31363 10308
rect 31379 10364 31443 10368
rect 31379 10308 31383 10364
rect 31383 10308 31439 10364
rect 31439 10308 31443 10364
rect 31379 10304 31443 10308
rect 31459 10364 31523 10368
rect 31459 10308 31463 10364
rect 31463 10308 31519 10364
rect 31519 10308 31523 10364
rect 31459 10304 31523 10308
rect 4252 9820 4316 9824
rect 4252 9764 4256 9820
rect 4256 9764 4312 9820
rect 4312 9764 4316 9820
rect 4252 9760 4316 9764
rect 4332 9820 4396 9824
rect 4332 9764 4336 9820
rect 4336 9764 4392 9820
rect 4392 9764 4396 9820
rect 4332 9760 4396 9764
rect 4412 9820 4476 9824
rect 4412 9764 4416 9820
rect 4416 9764 4472 9820
rect 4472 9764 4476 9820
rect 4412 9760 4476 9764
rect 4492 9820 4556 9824
rect 4492 9764 4496 9820
rect 4496 9764 4552 9820
rect 4552 9764 4556 9820
rect 4492 9760 4556 9764
rect 11957 9820 12021 9824
rect 11957 9764 11961 9820
rect 11961 9764 12017 9820
rect 12017 9764 12021 9820
rect 11957 9760 12021 9764
rect 12037 9820 12101 9824
rect 12037 9764 12041 9820
rect 12041 9764 12097 9820
rect 12097 9764 12101 9820
rect 12037 9760 12101 9764
rect 12117 9820 12181 9824
rect 12117 9764 12121 9820
rect 12121 9764 12177 9820
rect 12177 9764 12181 9820
rect 12117 9760 12181 9764
rect 12197 9820 12261 9824
rect 12197 9764 12201 9820
rect 12201 9764 12257 9820
rect 12257 9764 12261 9820
rect 12197 9760 12261 9764
rect 19662 9820 19726 9824
rect 19662 9764 19666 9820
rect 19666 9764 19722 9820
rect 19722 9764 19726 9820
rect 19662 9760 19726 9764
rect 19742 9820 19806 9824
rect 19742 9764 19746 9820
rect 19746 9764 19802 9820
rect 19802 9764 19806 9820
rect 19742 9760 19806 9764
rect 19822 9820 19886 9824
rect 19822 9764 19826 9820
rect 19826 9764 19882 9820
rect 19882 9764 19886 9820
rect 19822 9760 19886 9764
rect 19902 9820 19966 9824
rect 19902 9764 19906 9820
rect 19906 9764 19962 9820
rect 19962 9764 19966 9820
rect 19902 9760 19966 9764
rect 27367 9820 27431 9824
rect 27367 9764 27371 9820
rect 27371 9764 27427 9820
rect 27427 9764 27431 9820
rect 27367 9760 27431 9764
rect 27447 9820 27511 9824
rect 27447 9764 27451 9820
rect 27451 9764 27507 9820
rect 27507 9764 27511 9820
rect 27447 9760 27511 9764
rect 27527 9820 27591 9824
rect 27527 9764 27531 9820
rect 27531 9764 27587 9820
rect 27587 9764 27591 9820
rect 27527 9760 27591 9764
rect 27607 9820 27671 9824
rect 27607 9764 27611 9820
rect 27611 9764 27667 9820
rect 27667 9764 27671 9820
rect 27607 9760 27671 9764
rect 9628 9752 9692 9756
rect 9628 9696 9642 9752
rect 9642 9696 9692 9752
rect 9628 9692 9692 9696
rect 15516 9752 15580 9756
rect 15516 9696 15566 9752
rect 15566 9696 15580 9752
rect 15516 9692 15580 9696
rect 8104 9276 8168 9280
rect 8104 9220 8108 9276
rect 8108 9220 8164 9276
rect 8164 9220 8168 9276
rect 8104 9216 8168 9220
rect 8184 9276 8248 9280
rect 8184 9220 8188 9276
rect 8188 9220 8244 9276
rect 8244 9220 8248 9276
rect 8184 9216 8248 9220
rect 8264 9276 8328 9280
rect 8264 9220 8268 9276
rect 8268 9220 8324 9276
rect 8324 9220 8328 9276
rect 8264 9216 8328 9220
rect 8344 9276 8408 9280
rect 8344 9220 8348 9276
rect 8348 9220 8404 9276
rect 8404 9220 8408 9276
rect 8344 9216 8408 9220
rect 15809 9276 15873 9280
rect 15809 9220 15813 9276
rect 15813 9220 15869 9276
rect 15869 9220 15873 9276
rect 15809 9216 15873 9220
rect 15889 9276 15953 9280
rect 15889 9220 15893 9276
rect 15893 9220 15949 9276
rect 15949 9220 15953 9276
rect 15889 9216 15953 9220
rect 15969 9276 16033 9280
rect 15969 9220 15973 9276
rect 15973 9220 16029 9276
rect 16029 9220 16033 9276
rect 15969 9216 16033 9220
rect 16049 9276 16113 9280
rect 16049 9220 16053 9276
rect 16053 9220 16109 9276
rect 16109 9220 16113 9276
rect 16049 9216 16113 9220
rect 23514 9276 23578 9280
rect 23514 9220 23518 9276
rect 23518 9220 23574 9276
rect 23574 9220 23578 9276
rect 23514 9216 23578 9220
rect 23594 9276 23658 9280
rect 23594 9220 23598 9276
rect 23598 9220 23654 9276
rect 23654 9220 23658 9276
rect 23594 9216 23658 9220
rect 23674 9276 23738 9280
rect 23674 9220 23678 9276
rect 23678 9220 23734 9276
rect 23734 9220 23738 9276
rect 23674 9216 23738 9220
rect 23754 9276 23818 9280
rect 23754 9220 23758 9276
rect 23758 9220 23814 9276
rect 23814 9220 23818 9276
rect 23754 9216 23818 9220
rect 31219 9276 31283 9280
rect 31219 9220 31223 9276
rect 31223 9220 31279 9276
rect 31279 9220 31283 9276
rect 31219 9216 31283 9220
rect 31299 9276 31363 9280
rect 31299 9220 31303 9276
rect 31303 9220 31359 9276
rect 31359 9220 31363 9276
rect 31299 9216 31363 9220
rect 31379 9276 31443 9280
rect 31379 9220 31383 9276
rect 31383 9220 31439 9276
rect 31439 9220 31443 9276
rect 31379 9216 31443 9220
rect 31459 9276 31523 9280
rect 31459 9220 31463 9276
rect 31463 9220 31519 9276
rect 31519 9220 31523 9276
rect 31459 9216 31523 9220
rect 4252 8732 4316 8736
rect 4252 8676 4256 8732
rect 4256 8676 4312 8732
rect 4312 8676 4316 8732
rect 4252 8672 4316 8676
rect 4332 8732 4396 8736
rect 4332 8676 4336 8732
rect 4336 8676 4392 8732
rect 4392 8676 4396 8732
rect 4332 8672 4396 8676
rect 4412 8732 4476 8736
rect 4412 8676 4416 8732
rect 4416 8676 4472 8732
rect 4472 8676 4476 8732
rect 4412 8672 4476 8676
rect 4492 8732 4556 8736
rect 4492 8676 4496 8732
rect 4496 8676 4552 8732
rect 4552 8676 4556 8732
rect 4492 8672 4556 8676
rect 11957 8732 12021 8736
rect 11957 8676 11961 8732
rect 11961 8676 12017 8732
rect 12017 8676 12021 8732
rect 11957 8672 12021 8676
rect 12037 8732 12101 8736
rect 12037 8676 12041 8732
rect 12041 8676 12097 8732
rect 12097 8676 12101 8732
rect 12037 8672 12101 8676
rect 12117 8732 12181 8736
rect 12117 8676 12121 8732
rect 12121 8676 12177 8732
rect 12177 8676 12181 8732
rect 12117 8672 12181 8676
rect 12197 8732 12261 8736
rect 12197 8676 12201 8732
rect 12201 8676 12257 8732
rect 12257 8676 12261 8732
rect 12197 8672 12261 8676
rect 19662 8732 19726 8736
rect 19662 8676 19666 8732
rect 19666 8676 19722 8732
rect 19722 8676 19726 8732
rect 19662 8672 19726 8676
rect 19742 8732 19806 8736
rect 19742 8676 19746 8732
rect 19746 8676 19802 8732
rect 19802 8676 19806 8732
rect 19742 8672 19806 8676
rect 19822 8732 19886 8736
rect 19822 8676 19826 8732
rect 19826 8676 19882 8732
rect 19882 8676 19886 8732
rect 19822 8672 19886 8676
rect 19902 8732 19966 8736
rect 19902 8676 19906 8732
rect 19906 8676 19962 8732
rect 19962 8676 19966 8732
rect 19902 8672 19966 8676
rect 27367 8732 27431 8736
rect 27367 8676 27371 8732
rect 27371 8676 27427 8732
rect 27427 8676 27431 8732
rect 27367 8672 27431 8676
rect 27447 8732 27511 8736
rect 27447 8676 27451 8732
rect 27451 8676 27507 8732
rect 27507 8676 27511 8732
rect 27447 8672 27511 8676
rect 27527 8732 27591 8736
rect 27527 8676 27531 8732
rect 27531 8676 27587 8732
rect 27587 8676 27591 8732
rect 27527 8672 27591 8676
rect 27607 8732 27671 8736
rect 27607 8676 27611 8732
rect 27611 8676 27667 8732
rect 27667 8676 27671 8732
rect 27607 8672 27671 8676
rect 12572 8332 12636 8396
rect 8104 8188 8168 8192
rect 8104 8132 8108 8188
rect 8108 8132 8164 8188
rect 8164 8132 8168 8188
rect 8104 8128 8168 8132
rect 8184 8188 8248 8192
rect 8184 8132 8188 8188
rect 8188 8132 8244 8188
rect 8244 8132 8248 8188
rect 8184 8128 8248 8132
rect 8264 8188 8328 8192
rect 8264 8132 8268 8188
rect 8268 8132 8324 8188
rect 8324 8132 8328 8188
rect 8264 8128 8328 8132
rect 8344 8188 8408 8192
rect 8344 8132 8348 8188
rect 8348 8132 8404 8188
rect 8404 8132 8408 8188
rect 8344 8128 8408 8132
rect 15809 8188 15873 8192
rect 15809 8132 15813 8188
rect 15813 8132 15869 8188
rect 15869 8132 15873 8188
rect 15809 8128 15873 8132
rect 15889 8188 15953 8192
rect 15889 8132 15893 8188
rect 15893 8132 15949 8188
rect 15949 8132 15953 8188
rect 15889 8128 15953 8132
rect 15969 8188 16033 8192
rect 15969 8132 15973 8188
rect 15973 8132 16029 8188
rect 16029 8132 16033 8188
rect 15969 8128 16033 8132
rect 16049 8188 16113 8192
rect 16049 8132 16053 8188
rect 16053 8132 16109 8188
rect 16109 8132 16113 8188
rect 16049 8128 16113 8132
rect 23514 8188 23578 8192
rect 23514 8132 23518 8188
rect 23518 8132 23574 8188
rect 23574 8132 23578 8188
rect 23514 8128 23578 8132
rect 23594 8188 23658 8192
rect 23594 8132 23598 8188
rect 23598 8132 23654 8188
rect 23654 8132 23658 8188
rect 23594 8128 23658 8132
rect 23674 8188 23738 8192
rect 23674 8132 23678 8188
rect 23678 8132 23734 8188
rect 23734 8132 23738 8188
rect 23674 8128 23738 8132
rect 23754 8188 23818 8192
rect 23754 8132 23758 8188
rect 23758 8132 23814 8188
rect 23814 8132 23818 8188
rect 23754 8128 23818 8132
rect 31219 8188 31283 8192
rect 31219 8132 31223 8188
rect 31223 8132 31279 8188
rect 31279 8132 31283 8188
rect 31219 8128 31283 8132
rect 31299 8188 31363 8192
rect 31299 8132 31303 8188
rect 31303 8132 31359 8188
rect 31359 8132 31363 8188
rect 31299 8128 31363 8132
rect 31379 8188 31443 8192
rect 31379 8132 31383 8188
rect 31383 8132 31439 8188
rect 31439 8132 31443 8188
rect 31379 8128 31443 8132
rect 31459 8188 31523 8192
rect 31459 8132 31463 8188
rect 31463 8132 31519 8188
rect 31519 8132 31523 8188
rect 31459 8128 31523 8132
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 4332 7644 4396 7648
rect 4332 7588 4336 7644
rect 4336 7588 4392 7644
rect 4392 7588 4396 7644
rect 4332 7584 4396 7588
rect 4412 7644 4476 7648
rect 4412 7588 4416 7644
rect 4416 7588 4472 7644
rect 4472 7588 4476 7644
rect 4412 7584 4476 7588
rect 4492 7644 4556 7648
rect 4492 7588 4496 7644
rect 4496 7588 4552 7644
rect 4552 7588 4556 7644
rect 4492 7584 4556 7588
rect 11957 7644 12021 7648
rect 11957 7588 11961 7644
rect 11961 7588 12017 7644
rect 12017 7588 12021 7644
rect 11957 7584 12021 7588
rect 12037 7644 12101 7648
rect 12037 7588 12041 7644
rect 12041 7588 12097 7644
rect 12097 7588 12101 7644
rect 12037 7584 12101 7588
rect 12117 7644 12181 7648
rect 12117 7588 12121 7644
rect 12121 7588 12177 7644
rect 12177 7588 12181 7644
rect 12117 7584 12181 7588
rect 12197 7644 12261 7648
rect 12197 7588 12201 7644
rect 12201 7588 12257 7644
rect 12257 7588 12261 7644
rect 12197 7584 12261 7588
rect 19662 7644 19726 7648
rect 19662 7588 19666 7644
rect 19666 7588 19722 7644
rect 19722 7588 19726 7644
rect 19662 7584 19726 7588
rect 19742 7644 19806 7648
rect 19742 7588 19746 7644
rect 19746 7588 19802 7644
rect 19802 7588 19806 7644
rect 19742 7584 19806 7588
rect 19822 7644 19886 7648
rect 19822 7588 19826 7644
rect 19826 7588 19882 7644
rect 19882 7588 19886 7644
rect 19822 7584 19886 7588
rect 19902 7644 19966 7648
rect 19902 7588 19906 7644
rect 19906 7588 19962 7644
rect 19962 7588 19966 7644
rect 19902 7584 19966 7588
rect 27367 7644 27431 7648
rect 27367 7588 27371 7644
rect 27371 7588 27427 7644
rect 27427 7588 27431 7644
rect 27367 7584 27431 7588
rect 27447 7644 27511 7648
rect 27447 7588 27451 7644
rect 27451 7588 27507 7644
rect 27507 7588 27511 7644
rect 27447 7584 27511 7588
rect 27527 7644 27591 7648
rect 27527 7588 27531 7644
rect 27531 7588 27587 7644
rect 27587 7588 27591 7644
rect 27527 7584 27591 7588
rect 27607 7644 27671 7648
rect 27607 7588 27611 7644
rect 27611 7588 27667 7644
rect 27667 7588 27671 7644
rect 27607 7584 27671 7588
rect 8104 7100 8168 7104
rect 8104 7044 8108 7100
rect 8108 7044 8164 7100
rect 8164 7044 8168 7100
rect 8104 7040 8168 7044
rect 8184 7100 8248 7104
rect 8184 7044 8188 7100
rect 8188 7044 8244 7100
rect 8244 7044 8248 7100
rect 8184 7040 8248 7044
rect 8264 7100 8328 7104
rect 8264 7044 8268 7100
rect 8268 7044 8324 7100
rect 8324 7044 8328 7100
rect 8264 7040 8328 7044
rect 8344 7100 8408 7104
rect 8344 7044 8348 7100
rect 8348 7044 8404 7100
rect 8404 7044 8408 7100
rect 8344 7040 8408 7044
rect 15809 7100 15873 7104
rect 15809 7044 15813 7100
rect 15813 7044 15869 7100
rect 15869 7044 15873 7100
rect 15809 7040 15873 7044
rect 15889 7100 15953 7104
rect 15889 7044 15893 7100
rect 15893 7044 15949 7100
rect 15949 7044 15953 7100
rect 15889 7040 15953 7044
rect 15969 7100 16033 7104
rect 15969 7044 15973 7100
rect 15973 7044 16029 7100
rect 16029 7044 16033 7100
rect 15969 7040 16033 7044
rect 16049 7100 16113 7104
rect 16049 7044 16053 7100
rect 16053 7044 16109 7100
rect 16109 7044 16113 7100
rect 16049 7040 16113 7044
rect 23514 7100 23578 7104
rect 23514 7044 23518 7100
rect 23518 7044 23574 7100
rect 23574 7044 23578 7100
rect 23514 7040 23578 7044
rect 23594 7100 23658 7104
rect 23594 7044 23598 7100
rect 23598 7044 23654 7100
rect 23654 7044 23658 7100
rect 23594 7040 23658 7044
rect 23674 7100 23738 7104
rect 23674 7044 23678 7100
rect 23678 7044 23734 7100
rect 23734 7044 23738 7100
rect 23674 7040 23738 7044
rect 23754 7100 23818 7104
rect 23754 7044 23758 7100
rect 23758 7044 23814 7100
rect 23814 7044 23818 7100
rect 23754 7040 23818 7044
rect 31219 7100 31283 7104
rect 31219 7044 31223 7100
rect 31223 7044 31279 7100
rect 31279 7044 31283 7100
rect 31219 7040 31283 7044
rect 31299 7100 31363 7104
rect 31299 7044 31303 7100
rect 31303 7044 31359 7100
rect 31359 7044 31363 7100
rect 31299 7040 31363 7044
rect 31379 7100 31443 7104
rect 31379 7044 31383 7100
rect 31383 7044 31439 7100
rect 31439 7044 31443 7100
rect 31379 7040 31443 7044
rect 31459 7100 31523 7104
rect 31459 7044 31463 7100
rect 31463 7044 31519 7100
rect 31519 7044 31523 7100
rect 31459 7040 31523 7044
rect 9628 6836 9692 6900
rect 12572 6836 12636 6900
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 4332 6556 4396 6560
rect 4332 6500 4336 6556
rect 4336 6500 4392 6556
rect 4392 6500 4396 6556
rect 4332 6496 4396 6500
rect 4412 6556 4476 6560
rect 4412 6500 4416 6556
rect 4416 6500 4472 6556
rect 4472 6500 4476 6556
rect 4412 6496 4476 6500
rect 4492 6556 4556 6560
rect 4492 6500 4496 6556
rect 4496 6500 4552 6556
rect 4552 6500 4556 6556
rect 4492 6496 4556 6500
rect 11957 6556 12021 6560
rect 11957 6500 11961 6556
rect 11961 6500 12017 6556
rect 12017 6500 12021 6556
rect 11957 6496 12021 6500
rect 12037 6556 12101 6560
rect 12037 6500 12041 6556
rect 12041 6500 12097 6556
rect 12097 6500 12101 6556
rect 12037 6496 12101 6500
rect 12117 6556 12181 6560
rect 12117 6500 12121 6556
rect 12121 6500 12177 6556
rect 12177 6500 12181 6556
rect 12117 6496 12181 6500
rect 12197 6556 12261 6560
rect 12197 6500 12201 6556
rect 12201 6500 12257 6556
rect 12257 6500 12261 6556
rect 12197 6496 12261 6500
rect 19662 6556 19726 6560
rect 19662 6500 19666 6556
rect 19666 6500 19722 6556
rect 19722 6500 19726 6556
rect 19662 6496 19726 6500
rect 19742 6556 19806 6560
rect 19742 6500 19746 6556
rect 19746 6500 19802 6556
rect 19802 6500 19806 6556
rect 19742 6496 19806 6500
rect 19822 6556 19886 6560
rect 19822 6500 19826 6556
rect 19826 6500 19882 6556
rect 19882 6500 19886 6556
rect 19822 6496 19886 6500
rect 19902 6556 19966 6560
rect 19902 6500 19906 6556
rect 19906 6500 19962 6556
rect 19962 6500 19966 6556
rect 19902 6496 19966 6500
rect 27367 6556 27431 6560
rect 27367 6500 27371 6556
rect 27371 6500 27427 6556
rect 27427 6500 27431 6556
rect 27367 6496 27431 6500
rect 27447 6556 27511 6560
rect 27447 6500 27451 6556
rect 27451 6500 27507 6556
rect 27507 6500 27511 6556
rect 27447 6496 27511 6500
rect 27527 6556 27591 6560
rect 27527 6500 27531 6556
rect 27531 6500 27587 6556
rect 27587 6500 27591 6556
rect 27527 6496 27591 6500
rect 27607 6556 27671 6560
rect 27607 6500 27611 6556
rect 27611 6500 27667 6556
rect 27667 6500 27671 6556
rect 27607 6496 27671 6500
rect 8104 6012 8168 6016
rect 8104 5956 8108 6012
rect 8108 5956 8164 6012
rect 8164 5956 8168 6012
rect 8104 5952 8168 5956
rect 8184 6012 8248 6016
rect 8184 5956 8188 6012
rect 8188 5956 8244 6012
rect 8244 5956 8248 6012
rect 8184 5952 8248 5956
rect 8264 6012 8328 6016
rect 8264 5956 8268 6012
rect 8268 5956 8324 6012
rect 8324 5956 8328 6012
rect 8264 5952 8328 5956
rect 8344 6012 8408 6016
rect 8344 5956 8348 6012
rect 8348 5956 8404 6012
rect 8404 5956 8408 6012
rect 8344 5952 8408 5956
rect 15809 6012 15873 6016
rect 15809 5956 15813 6012
rect 15813 5956 15869 6012
rect 15869 5956 15873 6012
rect 15809 5952 15873 5956
rect 15889 6012 15953 6016
rect 15889 5956 15893 6012
rect 15893 5956 15949 6012
rect 15949 5956 15953 6012
rect 15889 5952 15953 5956
rect 15969 6012 16033 6016
rect 15969 5956 15973 6012
rect 15973 5956 16029 6012
rect 16029 5956 16033 6012
rect 15969 5952 16033 5956
rect 16049 6012 16113 6016
rect 16049 5956 16053 6012
rect 16053 5956 16109 6012
rect 16109 5956 16113 6012
rect 16049 5952 16113 5956
rect 23514 6012 23578 6016
rect 23514 5956 23518 6012
rect 23518 5956 23574 6012
rect 23574 5956 23578 6012
rect 23514 5952 23578 5956
rect 23594 6012 23658 6016
rect 23594 5956 23598 6012
rect 23598 5956 23654 6012
rect 23654 5956 23658 6012
rect 23594 5952 23658 5956
rect 23674 6012 23738 6016
rect 23674 5956 23678 6012
rect 23678 5956 23734 6012
rect 23734 5956 23738 6012
rect 23674 5952 23738 5956
rect 23754 6012 23818 6016
rect 23754 5956 23758 6012
rect 23758 5956 23814 6012
rect 23814 5956 23818 6012
rect 23754 5952 23818 5956
rect 31219 6012 31283 6016
rect 31219 5956 31223 6012
rect 31223 5956 31279 6012
rect 31279 5956 31283 6012
rect 31219 5952 31283 5956
rect 31299 6012 31363 6016
rect 31299 5956 31303 6012
rect 31303 5956 31359 6012
rect 31359 5956 31363 6012
rect 31299 5952 31363 5956
rect 31379 6012 31443 6016
rect 31379 5956 31383 6012
rect 31383 5956 31439 6012
rect 31439 5956 31443 6012
rect 31379 5952 31443 5956
rect 31459 6012 31523 6016
rect 31459 5956 31463 6012
rect 31463 5956 31519 6012
rect 31519 5956 31523 6012
rect 31459 5952 31523 5956
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 4332 5468 4396 5472
rect 4332 5412 4336 5468
rect 4336 5412 4392 5468
rect 4392 5412 4396 5468
rect 4332 5408 4396 5412
rect 4412 5468 4476 5472
rect 4412 5412 4416 5468
rect 4416 5412 4472 5468
rect 4472 5412 4476 5468
rect 4412 5408 4476 5412
rect 4492 5468 4556 5472
rect 4492 5412 4496 5468
rect 4496 5412 4552 5468
rect 4552 5412 4556 5468
rect 4492 5408 4556 5412
rect 11957 5468 12021 5472
rect 11957 5412 11961 5468
rect 11961 5412 12017 5468
rect 12017 5412 12021 5468
rect 11957 5408 12021 5412
rect 12037 5468 12101 5472
rect 12037 5412 12041 5468
rect 12041 5412 12097 5468
rect 12097 5412 12101 5468
rect 12037 5408 12101 5412
rect 12117 5468 12181 5472
rect 12117 5412 12121 5468
rect 12121 5412 12177 5468
rect 12177 5412 12181 5468
rect 12117 5408 12181 5412
rect 12197 5468 12261 5472
rect 12197 5412 12201 5468
rect 12201 5412 12257 5468
rect 12257 5412 12261 5468
rect 12197 5408 12261 5412
rect 19662 5468 19726 5472
rect 19662 5412 19666 5468
rect 19666 5412 19722 5468
rect 19722 5412 19726 5468
rect 19662 5408 19726 5412
rect 19742 5468 19806 5472
rect 19742 5412 19746 5468
rect 19746 5412 19802 5468
rect 19802 5412 19806 5468
rect 19742 5408 19806 5412
rect 19822 5468 19886 5472
rect 19822 5412 19826 5468
rect 19826 5412 19882 5468
rect 19882 5412 19886 5468
rect 19822 5408 19886 5412
rect 19902 5468 19966 5472
rect 19902 5412 19906 5468
rect 19906 5412 19962 5468
rect 19962 5412 19966 5468
rect 19902 5408 19966 5412
rect 27367 5468 27431 5472
rect 27367 5412 27371 5468
rect 27371 5412 27427 5468
rect 27427 5412 27431 5468
rect 27367 5408 27431 5412
rect 27447 5468 27511 5472
rect 27447 5412 27451 5468
rect 27451 5412 27507 5468
rect 27507 5412 27511 5468
rect 27447 5408 27511 5412
rect 27527 5468 27591 5472
rect 27527 5412 27531 5468
rect 27531 5412 27587 5468
rect 27587 5412 27591 5468
rect 27527 5408 27591 5412
rect 27607 5468 27671 5472
rect 27607 5412 27611 5468
rect 27611 5412 27667 5468
rect 27667 5412 27671 5468
rect 27607 5408 27671 5412
rect 8104 4924 8168 4928
rect 8104 4868 8108 4924
rect 8108 4868 8164 4924
rect 8164 4868 8168 4924
rect 8104 4864 8168 4868
rect 8184 4924 8248 4928
rect 8184 4868 8188 4924
rect 8188 4868 8244 4924
rect 8244 4868 8248 4924
rect 8184 4864 8248 4868
rect 8264 4924 8328 4928
rect 8264 4868 8268 4924
rect 8268 4868 8324 4924
rect 8324 4868 8328 4924
rect 8264 4864 8328 4868
rect 8344 4924 8408 4928
rect 8344 4868 8348 4924
rect 8348 4868 8404 4924
rect 8404 4868 8408 4924
rect 8344 4864 8408 4868
rect 15809 4924 15873 4928
rect 15809 4868 15813 4924
rect 15813 4868 15869 4924
rect 15869 4868 15873 4924
rect 15809 4864 15873 4868
rect 15889 4924 15953 4928
rect 15889 4868 15893 4924
rect 15893 4868 15949 4924
rect 15949 4868 15953 4924
rect 15889 4864 15953 4868
rect 15969 4924 16033 4928
rect 15969 4868 15973 4924
rect 15973 4868 16029 4924
rect 16029 4868 16033 4924
rect 15969 4864 16033 4868
rect 16049 4924 16113 4928
rect 16049 4868 16053 4924
rect 16053 4868 16109 4924
rect 16109 4868 16113 4924
rect 16049 4864 16113 4868
rect 23514 4924 23578 4928
rect 23514 4868 23518 4924
rect 23518 4868 23574 4924
rect 23574 4868 23578 4924
rect 23514 4864 23578 4868
rect 23594 4924 23658 4928
rect 23594 4868 23598 4924
rect 23598 4868 23654 4924
rect 23654 4868 23658 4924
rect 23594 4864 23658 4868
rect 23674 4924 23738 4928
rect 23674 4868 23678 4924
rect 23678 4868 23734 4924
rect 23734 4868 23738 4924
rect 23674 4864 23738 4868
rect 23754 4924 23818 4928
rect 23754 4868 23758 4924
rect 23758 4868 23814 4924
rect 23814 4868 23818 4924
rect 23754 4864 23818 4868
rect 31219 4924 31283 4928
rect 31219 4868 31223 4924
rect 31223 4868 31279 4924
rect 31279 4868 31283 4924
rect 31219 4864 31283 4868
rect 31299 4924 31363 4928
rect 31299 4868 31303 4924
rect 31303 4868 31359 4924
rect 31359 4868 31363 4924
rect 31299 4864 31363 4868
rect 31379 4924 31443 4928
rect 31379 4868 31383 4924
rect 31383 4868 31439 4924
rect 31439 4868 31443 4924
rect 31379 4864 31443 4868
rect 31459 4924 31523 4928
rect 31459 4868 31463 4924
rect 31463 4868 31519 4924
rect 31519 4868 31523 4924
rect 31459 4864 31523 4868
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 4332 4380 4396 4384
rect 4332 4324 4336 4380
rect 4336 4324 4392 4380
rect 4392 4324 4396 4380
rect 4332 4320 4396 4324
rect 4412 4380 4476 4384
rect 4412 4324 4416 4380
rect 4416 4324 4472 4380
rect 4472 4324 4476 4380
rect 4412 4320 4476 4324
rect 4492 4380 4556 4384
rect 4492 4324 4496 4380
rect 4496 4324 4552 4380
rect 4552 4324 4556 4380
rect 4492 4320 4556 4324
rect 11957 4380 12021 4384
rect 11957 4324 11961 4380
rect 11961 4324 12017 4380
rect 12017 4324 12021 4380
rect 11957 4320 12021 4324
rect 12037 4380 12101 4384
rect 12037 4324 12041 4380
rect 12041 4324 12097 4380
rect 12097 4324 12101 4380
rect 12037 4320 12101 4324
rect 12117 4380 12181 4384
rect 12117 4324 12121 4380
rect 12121 4324 12177 4380
rect 12177 4324 12181 4380
rect 12117 4320 12181 4324
rect 12197 4380 12261 4384
rect 12197 4324 12201 4380
rect 12201 4324 12257 4380
rect 12257 4324 12261 4380
rect 12197 4320 12261 4324
rect 19662 4380 19726 4384
rect 19662 4324 19666 4380
rect 19666 4324 19722 4380
rect 19722 4324 19726 4380
rect 19662 4320 19726 4324
rect 19742 4380 19806 4384
rect 19742 4324 19746 4380
rect 19746 4324 19802 4380
rect 19802 4324 19806 4380
rect 19742 4320 19806 4324
rect 19822 4380 19886 4384
rect 19822 4324 19826 4380
rect 19826 4324 19882 4380
rect 19882 4324 19886 4380
rect 19822 4320 19886 4324
rect 19902 4380 19966 4384
rect 19902 4324 19906 4380
rect 19906 4324 19962 4380
rect 19962 4324 19966 4380
rect 19902 4320 19966 4324
rect 27367 4380 27431 4384
rect 27367 4324 27371 4380
rect 27371 4324 27427 4380
rect 27427 4324 27431 4380
rect 27367 4320 27431 4324
rect 27447 4380 27511 4384
rect 27447 4324 27451 4380
rect 27451 4324 27507 4380
rect 27507 4324 27511 4380
rect 27447 4320 27511 4324
rect 27527 4380 27591 4384
rect 27527 4324 27531 4380
rect 27531 4324 27587 4380
rect 27587 4324 27591 4380
rect 27527 4320 27591 4324
rect 27607 4380 27671 4384
rect 27607 4324 27611 4380
rect 27611 4324 27667 4380
rect 27667 4324 27671 4380
rect 27607 4320 27671 4324
rect 15516 4040 15580 4044
rect 15516 3984 15530 4040
rect 15530 3984 15580 4040
rect 15516 3980 15580 3984
rect 8104 3836 8168 3840
rect 8104 3780 8108 3836
rect 8108 3780 8164 3836
rect 8164 3780 8168 3836
rect 8104 3776 8168 3780
rect 8184 3836 8248 3840
rect 8184 3780 8188 3836
rect 8188 3780 8244 3836
rect 8244 3780 8248 3836
rect 8184 3776 8248 3780
rect 8264 3836 8328 3840
rect 8264 3780 8268 3836
rect 8268 3780 8324 3836
rect 8324 3780 8328 3836
rect 8264 3776 8328 3780
rect 8344 3836 8408 3840
rect 8344 3780 8348 3836
rect 8348 3780 8404 3836
rect 8404 3780 8408 3836
rect 8344 3776 8408 3780
rect 15809 3836 15873 3840
rect 15809 3780 15813 3836
rect 15813 3780 15869 3836
rect 15869 3780 15873 3836
rect 15809 3776 15873 3780
rect 15889 3836 15953 3840
rect 15889 3780 15893 3836
rect 15893 3780 15949 3836
rect 15949 3780 15953 3836
rect 15889 3776 15953 3780
rect 15969 3836 16033 3840
rect 15969 3780 15973 3836
rect 15973 3780 16029 3836
rect 16029 3780 16033 3836
rect 15969 3776 16033 3780
rect 16049 3836 16113 3840
rect 16049 3780 16053 3836
rect 16053 3780 16109 3836
rect 16109 3780 16113 3836
rect 16049 3776 16113 3780
rect 23514 3836 23578 3840
rect 23514 3780 23518 3836
rect 23518 3780 23574 3836
rect 23574 3780 23578 3836
rect 23514 3776 23578 3780
rect 23594 3836 23658 3840
rect 23594 3780 23598 3836
rect 23598 3780 23654 3836
rect 23654 3780 23658 3836
rect 23594 3776 23658 3780
rect 23674 3836 23738 3840
rect 23674 3780 23678 3836
rect 23678 3780 23734 3836
rect 23734 3780 23738 3836
rect 23674 3776 23738 3780
rect 23754 3836 23818 3840
rect 23754 3780 23758 3836
rect 23758 3780 23814 3836
rect 23814 3780 23818 3836
rect 23754 3776 23818 3780
rect 31219 3836 31283 3840
rect 31219 3780 31223 3836
rect 31223 3780 31279 3836
rect 31279 3780 31283 3836
rect 31219 3776 31283 3780
rect 31299 3836 31363 3840
rect 31299 3780 31303 3836
rect 31303 3780 31359 3836
rect 31359 3780 31363 3836
rect 31299 3776 31363 3780
rect 31379 3836 31443 3840
rect 31379 3780 31383 3836
rect 31383 3780 31439 3836
rect 31439 3780 31443 3836
rect 31379 3776 31443 3780
rect 31459 3836 31523 3840
rect 31459 3780 31463 3836
rect 31463 3780 31519 3836
rect 31519 3780 31523 3836
rect 31459 3776 31523 3780
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 4332 3292 4396 3296
rect 4332 3236 4336 3292
rect 4336 3236 4392 3292
rect 4392 3236 4396 3292
rect 4332 3232 4396 3236
rect 4412 3292 4476 3296
rect 4412 3236 4416 3292
rect 4416 3236 4472 3292
rect 4472 3236 4476 3292
rect 4412 3232 4476 3236
rect 4492 3292 4556 3296
rect 4492 3236 4496 3292
rect 4496 3236 4552 3292
rect 4552 3236 4556 3292
rect 4492 3232 4556 3236
rect 11957 3292 12021 3296
rect 11957 3236 11961 3292
rect 11961 3236 12017 3292
rect 12017 3236 12021 3292
rect 11957 3232 12021 3236
rect 12037 3292 12101 3296
rect 12037 3236 12041 3292
rect 12041 3236 12097 3292
rect 12097 3236 12101 3292
rect 12037 3232 12101 3236
rect 12117 3292 12181 3296
rect 12117 3236 12121 3292
rect 12121 3236 12177 3292
rect 12177 3236 12181 3292
rect 12117 3232 12181 3236
rect 12197 3292 12261 3296
rect 12197 3236 12201 3292
rect 12201 3236 12257 3292
rect 12257 3236 12261 3292
rect 12197 3232 12261 3236
rect 19662 3292 19726 3296
rect 19662 3236 19666 3292
rect 19666 3236 19722 3292
rect 19722 3236 19726 3292
rect 19662 3232 19726 3236
rect 19742 3292 19806 3296
rect 19742 3236 19746 3292
rect 19746 3236 19802 3292
rect 19802 3236 19806 3292
rect 19742 3232 19806 3236
rect 19822 3292 19886 3296
rect 19822 3236 19826 3292
rect 19826 3236 19882 3292
rect 19882 3236 19886 3292
rect 19822 3232 19886 3236
rect 19902 3292 19966 3296
rect 19902 3236 19906 3292
rect 19906 3236 19962 3292
rect 19962 3236 19966 3292
rect 19902 3232 19966 3236
rect 27367 3292 27431 3296
rect 27367 3236 27371 3292
rect 27371 3236 27427 3292
rect 27427 3236 27431 3292
rect 27367 3232 27431 3236
rect 27447 3292 27511 3296
rect 27447 3236 27451 3292
rect 27451 3236 27507 3292
rect 27507 3236 27511 3292
rect 27447 3232 27511 3236
rect 27527 3292 27591 3296
rect 27527 3236 27531 3292
rect 27531 3236 27587 3292
rect 27587 3236 27591 3292
rect 27527 3232 27591 3236
rect 27607 3292 27671 3296
rect 27607 3236 27611 3292
rect 27611 3236 27667 3292
rect 27667 3236 27671 3292
rect 27607 3232 27671 3236
rect 8104 2748 8168 2752
rect 8104 2692 8108 2748
rect 8108 2692 8164 2748
rect 8164 2692 8168 2748
rect 8104 2688 8168 2692
rect 8184 2748 8248 2752
rect 8184 2692 8188 2748
rect 8188 2692 8244 2748
rect 8244 2692 8248 2748
rect 8184 2688 8248 2692
rect 8264 2748 8328 2752
rect 8264 2692 8268 2748
rect 8268 2692 8324 2748
rect 8324 2692 8328 2748
rect 8264 2688 8328 2692
rect 8344 2748 8408 2752
rect 8344 2692 8348 2748
rect 8348 2692 8404 2748
rect 8404 2692 8408 2748
rect 8344 2688 8408 2692
rect 15809 2748 15873 2752
rect 15809 2692 15813 2748
rect 15813 2692 15869 2748
rect 15869 2692 15873 2748
rect 15809 2688 15873 2692
rect 15889 2748 15953 2752
rect 15889 2692 15893 2748
rect 15893 2692 15949 2748
rect 15949 2692 15953 2748
rect 15889 2688 15953 2692
rect 15969 2748 16033 2752
rect 15969 2692 15973 2748
rect 15973 2692 16029 2748
rect 16029 2692 16033 2748
rect 15969 2688 16033 2692
rect 16049 2748 16113 2752
rect 16049 2692 16053 2748
rect 16053 2692 16109 2748
rect 16109 2692 16113 2748
rect 16049 2688 16113 2692
rect 23514 2748 23578 2752
rect 23514 2692 23518 2748
rect 23518 2692 23574 2748
rect 23574 2692 23578 2748
rect 23514 2688 23578 2692
rect 23594 2748 23658 2752
rect 23594 2692 23598 2748
rect 23598 2692 23654 2748
rect 23654 2692 23658 2748
rect 23594 2688 23658 2692
rect 23674 2748 23738 2752
rect 23674 2692 23678 2748
rect 23678 2692 23734 2748
rect 23734 2692 23738 2748
rect 23674 2688 23738 2692
rect 23754 2748 23818 2752
rect 23754 2692 23758 2748
rect 23758 2692 23814 2748
rect 23814 2692 23818 2748
rect 23754 2688 23818 2692
rect 31219 2748 31283 2752
rect 31219 2692 31223 2748
rect 31223 2692 31279 2748
rect 31279 2692 31283 2748
rect 31219 2688 31283 2692
rect 31299 2748 31363 2752
rect 31299 2692 31303 2748
rect 31303 2692 31359 2748
rect 31359 2692 31363 2748
rect 31299 2688 31363 2692
rect 31379 2748 31443 2752
rect 31379 2692 31383 2748
rect 31383 2692 31439 2748
rect 31439 2692 31443 2748
rect 31379 2688 31443 2692
rect 31459 2748 31523 2752
rect 31459 2692 31463 2748
rect 31463 2692 31519 2748
rect 31519 2692 31523 2748
rect 31459 2688 31523 2692
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 4332 2204 4396 2208
rect 4332 2148 4336 2204
rect 4336 2148 4392 2204
rect 4392 2148 4396 2204
rect 4332 2144 4396 2148
rect 4412 2204 4476 2208
rect 4412 2148 4416 2204
rect 4416 2148 4472 2204
rect 4472 2148 4476 2204
rect 4412 2144 4476 2148
rect 4492 2204 4556 2208
rect 4492 2148 4496 2204
rect 4496 2148 4552 2204
rect 4552 2148 4556 2204
rect 4492 2144 4556 2148
rect 11957 2204 12021 2208
rect 11957 2148 11961 2204
rect 11961 2148 12017 2204
rect 12017 2148 12021 2204
rect 11957 2144 12021 2148
rect 12037 2204 12101 2208
rect 12037 2148 12041 2204
rect 12041 2148 12097 2204
rect 12097 2148 12101 2204
rect 12037 2144 12101 2148
rect 12117 2204 12181 2208
rect 12117 2148 12121 2204
rect 12121 2148 12177 2204
rect 12177 2148 12181 2204
rect 12117 2144 12181 2148
rect 12197 2204 12261 2208
rect 12197 2148 12201 2204
rect 12201 2148 12257 2204
rect 12257 2148 12261 2204
rect 12197 2144 12261 2148
rect 19662 2204 19726 2208
rect 19662 2148 19666 2204
rect 19666 2148 19722 2204
rect 19722 2148 19726 2204
rect 19662 2144 19726 2148
rect 19742 2204 19806 2208
rect 19742 2148 19746 2204
rect 19746 2148 19802 2204
rect 19802 2148 19806 2204
rect 19742 2144 19806 2148
rect 19822 2204 19886 2208
rect 19822 2148 19826 2204
rect 19826 2148 19882 2204
rect 19882 2148 19886 2204
rect 19822 2144 19886 2148
rect 19902 2204 19966 2208
rect 19902 2148 19906 2204
rect 19906 2148 19962 2204
rect 19962 2148 19966 2204
rect 19902 2144 19966 2148
rect 27367 2204 27431 2208
rect 27367 2148 27371 2204
rect 27371 2148 27427 2204
rect 27427 2148 27431 2204
rect 27367 2144 27431 2148
rect 27447 2204 27511 2208
rect 27447 2148 27451 2204
rect 27451 2148 27507 2204
rect 27507 2148 27511 2204
rect 27447 2144 27511 2148
rect 27527 2204 27591 2208
rect 27527 2148 27531 2204
rect 27531 2148 27587 2204
rect 27587 2148 27591 2204
rect 27527 2144 27591 2148
rect 27607 2204 27671 2208
rect 27607 2148 27611 2204
rect 27611 2148 27667 2204
rect 27667 2148 27671 2204
rect 27607 2144 27671 2148
rect 8104 1660 8168 1664
rect 8104 1604 8108 1660
rect 8108 1604 8164 1660
rect 8164 1604 8168 1660
rect 8104 1600 8168 1604
rect 8184 1660 8248 1664
rect 8184 1604 8188 1660
rect 8188 1604 8244 1660
rect 8244 1604 8248 1660
rect 8184 1600 8248 1604
rect 8264 1660 8328 1664
rect 8264 1604 8268 1660
rect 8268 1604 8324 1660
rect 8324 1604 8328 1660
rect 8264 1600 8328 1604
rect 8344 1660 8408 1664
rect 8344 1604 8348 1660
rect 8348 1604 8404 1660
rect 8404 1604 8408 1660
rect 8344 1600 8408 1604
rect 15809 1660 15873 1664
rect 15809 1604 15813 1660
rect 15813 1604 15869 1660
rect 15869 1604 15873 1660
rect 15809 1600 15873 1604
rect 15889 1660 15953 1664
rect 15889 1604 15893 1660
rect 15893 1604 15949 1660
rect 15949 1604 15953 1660
rect 15889 1600 15953 1604
rect 15969 1660 16033 1664
rect 15969 1604 15973 1660
rect 15973 1604 16029 1660
rect 16029 1604 16033 1660
rect 15969 1600 16033 1604
rect 16049 1660 16113 1664
rect 16049 1604 16053 1660
rect 16053 1604 16109 1660
rect 16109 1604 16113 1660
rect 16049 1600 16113 1604
rect 23514 1660 23578 1664
rect 23514 1604 23518 1660
rect 23518 1604 23574 1660
rect 23574 1604 23578 1660
rect 23514 1600 23578 1604
rect 23594 1660 23658 1664
rect 23594 1604 23598 1660
rect 23598 1604 23654 1660
rect 23654 1604 23658 1660
rect 23594 1600 23658 1604
rect 23674 1660 23738 1664
rect 23674 1604 23678 1660
rect 23678 1604 23734 1660
rect 23734 1604 23738 1660
rect 23674 1600 23738 1604
rect 23754 1660 23818 1664
rect 23754 1604 23758 1660
rect 23758 1604 23814 1660
rect 23814 1604 23818 1660
rect 23754 1600 23818 1604
rect 31219 1660 31283 1664
rect 31219 1604 31223 1660
rect 31223 1604 31279 1660
rect 31279 1604 31283 1660
rect 31219 1600 31283 1604
rect 31299 1660 31363 1664
rect 31299 1604 31303 1660
rect 31303 1604 31359 1660
rect 31359 1604 31363 1660
rect 31299 1600 31363 1604
rect 31379 1660 31443 1664
rect 31379 1604 31383 1660
rect 31383 1604 31439 1660
rect 31439 1604 31443 1660
rect 31379 1600 31443 1604
rect 31459 1660 31523 1664
rect 31459 1604 31463 1660
rect 31463 1604 31519 1660
rect 31519 1604 31523 1660
rect 31459 1600 31523 1604
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 4332 1116 4396 1120
rect 4332 1060 4336 1116
rect 4336 1060 4392 1116
rect 4392 1060 4396 1116
rect 4332 1056 4396 1060
rect 4412 1116 4476 1120
rect 4412 1060 4416 1116
rect 4416 1060 4472 1116
rect 4472 1060 4476 1116
rect 4412 1056 4476 1060
rect 4492 1116 4556 1120
rect 4492 1060 4496 1116
rect 4496 1060 4552 1116
rect 4552 1060 4556 1116
rect 4492 1056 4556 1060
rect 11957 1116 12021 1120
rect 11957 1060 11961 1116
rect 11961 1060 12017 1116
rect 12017 1060 12021 1116
rect 11957 1056 12021 1060
rect 12037 1116 12101 1120
rect 12037 1060 12041 1116
rect 12041 1060 12097 1116
rect 12097 1060 12101 1116
rect 12037 1056 12101 1060
rect 12117 1116 12181 1120
rect 12117 1060 12121 1116
rect 12121 1060 12177 1116
rect 12177 1060 12181 1116
rect 12117 1056 12181 1060
rect 12197 1116 12261 1120
rect 12197 1060 12201 1116
rect 12201 1060 12257 1116
rect 12257 1060 12261 1116
rect 12197 1056 12261 1060
rect 19662 1116 19726 1120
rect 19662 1060 19666 1116
rect 19666 1060 19722 1116
rect 19722 1060 19726 1116
rect 19662 1056 19726 1060
rect 19742 1116 19806 1120
rect 19742 1060 19746 1116
rect 19746 1060 19802 1116
rect 19802 1060 19806 1116
rect 19742 1056 19806 1060
rect 19822 1116 19886 1120
rect 19822 1060 19826 1116
rect 19826 1060 19882 1116
rect 19882 1060 19886 1116
rect 19822 1056 19886 1060
rect 19902 1116 19966 1120
rect 19902 1060 19906 1116
rect 19906 1060 19962 1116
rect 19962 1060 19966 1116
rect 19902 1056 19966 1060
rect 27367 1116 27431 1120
rect 27367 1060 27371 1116
rect 27371 1060 27427 1116
rect 27427 1060 27431 1116
rect 27367 1056 27431 1060
rect 27447 1116 27511 1120
rect 27447 1060 27451 1116
rect 27451 1060 27507 1116
rect 27507 1060 27511 1116
rect 27447 1056 27511 1060
rect 27527 1116 27591 1120
rect 27527 1060 27531 1116
rect 27531 1060 27587 1116
rect 27587 1060 27591 1116
rect 27527 1056 27591 1060
rect 27607 1116 27671 1120
rect 27607 1060 27611 1116
rect 27611 1060 27667 1116
rect 27667 1060 27671 1116
rect 27607 1056 27671 1060
rect 8104 572 8168 576
rect 8104 516 8108 572
rect 8108 516 8164 572
rect 8164 516 8168 572
rect 8104 512 8168 516
rect 8184 572 8248 576
rect 8184 516 8188 572
rect 8188 516 8244 572
rect 8244 516 8248 572
rect 8184 512 8248 516
rect 8264 572 8328 576
rect 8264 516 8268 572
rect 8268 516 8324 572
rect 8324 516 8328 572
rect 8264 512 8328 516
rect 8344 572 8408 576
rect 8344 516 8348 572
rect 8348 516 8404 572
rect 8404 516 8408 572
rect 8344 512 8408 516
rect 15809 572 15873 576
rect 15809 516 15813 572
rect 15813 516 15869 572
rect 15869 516 15873 572
rect 15809 512 15873 516
rect 15889 572 15953 576
rect 15889 516 15893 572
rect 15893 516 15949 572
rect 15949 516 15953 572
rect 15889 512 15953 516
rect 15969 572 16033 576
rect 15969 516 15973 572
rect 15973 516 16029 572
rect 16029 516 16033 572
rect 15969 512 16033 516
rect 16049 572 16113 576
rect 16049 516 16053 572
rect 16053 516 16109 572
rect 16109 516 16113 572
rect 16049 512 16113 516
rect 23514 572 23578 576
rect 23514 516 23518 572
rect 23518 516 23574 572
rect 23574 516 23578 572
rect 23514 512 23578 516
rect 23594 572 23658 576
rect 23594 516 23598 572
rect 23598 516 23654 572
rect 23654 516 23658 572
rect 23594 512 23658 516
rect 23674 572 23738 576
rect 23674 516 23678 572
rect 23678 516 23734 572
rect 23734 516 23738 572
rect 23674 512 23738 516
rect 23754 572 23818 576
rect 23754 516 23758 572
rect 23758 516 23814 572
rect 23814 516 23818 572
rect 23754 512 23818 516
rect 31219 572 31283 576
rect 31219 516 31223 572
rect 31223 516 31279 572
rect 31279 516 31283 572
rect 31219 512 31283 516
rect 31299 572 31363 576
rect 31299 516 31303 572
rect 31303 516 31359 572
rect 31359 516 31363 572
rect 31299 512 31363 516
rect 31379 572 31443 576
rect 31379 516 31383 572
rect 31383 516 31439 572
rect 31439 516 31443 572
rect 31379 512 31443 516
rect 31459 572 31523 576
rect 31459 516 31463 572
rect 31463 516 31519 572
rect 31519 516 31523 572
rect 31459 512 31523 516
<< metal4 >>
rect 4244 18528 4564 19088
rect 4244 18464 4252 18528
rect 4316 18464 4332 18528
rect 4396 18464 4412 18528
rect 4476 18464 4492 18528
rect 4556 18464 4564 18528
rect 4244 17440 4564 18464
rect 4244 17376 4252 17440
rect 4316 17376 4332 17440
rect 4396 17376 4412 17440
rect 4476 17376 4492 17440
rect 4556 17376 4564 17440
rect 4244 16352 4564 17376
rect 4244 16288 4252 16352
rect 4316 16288 4332 16352
rect 4396 16288 4412 16352
rect 4476 16288 4492 16352
rect 4556 16288 4564 16352
rect 4244 15264 4564 16288
rect 4244 15200 4252 15264
rect 4316 15200 4332 15264
rect 4396 15200 4412 15264
rect 4476 15200 4492 15264
rect 4556 15200 4564 15264
rect 4244 14176 4564 15200
rect 4244 14112 4252 14176
rect 4316 14112 4332 14176
rect 4396 14112 4412 14176
rect 4476 14112 4492 14176
rect 4556 14112 4564 14176
rect 4244 13088 4564 14112
rect 4244 13024 4252 13088
rect 4316 13024 4332 13088
rect 4396 13024 4412 13088
rect 4476 13024 4492 13088
rect 4556 13024 4564 13088
rect 4244 12000 4564 13024
rect 4244 11936 4252 12000
rect 4316 11936 4332 12000
rect 4396 11936 4412 12000
rect 4476 11936 4492 12000
rect 4556 11936 4564 12000
rect 4244 10912 4564 11936
rect 4244 10848 4252 10912
rect 4316 10848 4332 10912
rect 4396 10848 4412 10912
rect 4476 10848 4492 10912
rect 4556 10848 4564 10912
rect 4244 9824 4564 10848
rect 4244 9760 4252 9824
rect 4316 9760 4332 9824
rect 4396 9760 4412 9824
rect 4476 9760 4492 9824
rect 4556 9760 4564 9824
rect 4244 8736 4564 9760
rect 4244 8672 4252 8736
rect 4316 8672 4332 8736
rect 4396 8672 4412 8736
rect 4476 8672 4492 8736
rect 4556 8672 4564 8736
rect 4244 7648 4564 8672
rect 4244 7584 4252 7648
rect 4316 7584 4332 7648
rect 4396 7584 4412 7648
rect 4476 7584 4492 7648
rect 4556 7584 4564 7648
rect 4244 6560 4564 7584
rect 4244 6496 4252 6560
rect 4316 6496 4332 6560
rect 4396 6496 4412 6560
rect 4476 6496 4492 6560
rect 4556 6496 4564 6560
rect 4244 5472 4564 6496
rect 4244 5408 4252 5472
rect 4316 5408 4332 5472
rect 4396 5408 4412 5472
rect 4476 5408 4492 5472
rect 4556 5408 4564 5472
rect 4244 4384 4564 5408
rect 4244 4320 4252 4384
rect 4316 4320 4332 4384
rect 4396 4320 4412 4384
rect 4476 4320 4492 4384
rect 4556 4320 4564 4384
rect 4244 3296 4564 4320
rect 4244 3232 4252 3296
rect 4316 3232 4332 3296
rect 4396 3232 4412 3296
rect 4476 3232 4492 3296
rect 4556 3232 4564 3296
rect 4244 2208 4564 3232
rect 4244 2144 4252 2208
rect 4316 2144 4332 2208
rect 4396 2144 4412 2208
rect 4476 2144 4492 2208
rect 4556 2144 4564 2208
rect 4244 1120 4564 2144
rect 4244 1056 4252 1120
rect 4316 1056 4332 1120
rect 4396 1056 4412 1120
rect 4476 1056 4492 1120
rect 4556 1056 4564 1120
rect 4244 496 4564 1056
rect 8096 19072 8416 19088
rect 8096 19008 8104 19072
rect 8168 19008 8184 19072
rect 8248 19008 8264 19072
rect 8328 19008 8344 19072
rect 8408 19008 8416 19072
rect 8096 17984 8416 19008
rect 8096 17920 8104 17984
rect 8168 17920 8184 17984
rect 8248 17920 8264 17984
rect 8328 17920 8344 17984
rect 8408 17920 8416 17984
rect 8096 16896 8416 17920
rect 8096 16832 8104 16896
rect 8168 16832 8184 16896
rect 8248 16832 8264 16896
rect 8328 16832 8344 16896
rect 8408 16832 8416 16896
rect 8096 15808 8416 16832
rect 8096 15744 8104 15808
rect 8168 15744 8184 15808
rect 8248 15744 8264 15808
rect 8328 15744 8344 15808
rect 8408 15744 8416 15808
rect 8096 14720 8416 15744
rect 8096 14656 8104 14720
rect 8168 14656 8184 14720
rect 8248 14656 8264 14720
rect 8328 14656 8344 14720
rect 8408 14656 8416 14720
rect 8096 13632 8416 14656
rect 8096 13568 8104 13632
rect 8168 13568 8184 13632
rect 8248 13568 8264 13632
rect 8328 13568 8344 13632
rect 8408 13568 8416 13632
rect 8096 12544 8416 13568
rect 8096 12480 8104 12544
rect 8168 12480 8184 12544
rect 8248 12480 8264 12544
rect 8328 12480 8344 12544
rect 8408 12480 8416 12544
rect 8096 11456 8416 12480
rect 8096 11392 8104 11456
rect 8168 11392 8184 11456
rect 8248 11392 8264 11456
rect 8328 11392 8344 11456
rect 8408 11392 8416 11456
rect 8096 10368 8416 11392
rect 8096 10304 8104 10368
rect 8168 10304 8184 10368
rect 8248 10304 8264 10368
rect 8328 10304 8344 10368
rect 8408 10304 8416 10368
rect 8096 9280 8416 10304
rect 11949 18528 12269 19088
rect 11949 18464 11957 18528
rect 12021 18464 12037 18528
rect 12101 18464 12117 18528
rect 12181 18464 12197 18528
rect 12261 18464 12269 18528
rect 11949 17440 12269 18464
rect 11949 17376 11957 17440
rect 12021 17376 12037 17440
rect 12101 17376 12117 17440
rect 12181 17376 12197 17440
rect 12261 17376 12269 17440
rect 11949 16352 12269 17376
rect 11949 16288 11957 16352
rect 12021 16288 12037 16352
rect 12101 16288 12117 16352
rect 12181 16288 12197 16352
rect 12261 16288 12269 16352
rect 11949 15264 12269 16288
rect 11949 15200 11957 15264
rect 12021 15200 12037 15264
rect 12101 15200 12117 15264
rect 12181 15200 12197 15264
rect 12261 15200 12269 15264
rect 11949 14176 12269 15200
rect 11949 14112 11957 14176
rect 12021 14112 12037 14176
rect 12101 14112 12117 14176
rect 12181 14112 12197 14176
rect 12261 14112 12269 14176
rect 11949 13088 12269 14112
rect 11949 13024 11957 13088
rect 12021 13024 12037 13088
rect 12101 13024 12117 13088
rect 12181 13024 12197 13088
rect 12261 13024 12269 13088
rect 11949 12000 12269 13024
rect 11949 11936 11957 12000
rect 12021 11936 12037 12000
rect 12101 11936 12117 12000
rect 12181 11936 12197 12000
rect 12261 11936 12269 12000
rect 11949 10912 12269 11936
rect 11949 10848 11957 10912
rect 12021 10848 12037 10912
rect 12101 10848 12117 10912
rect 12181 10848 12197 10912
rect 12261 10848 12269 10912
rect 11949 9824 12269 10848
rect 11949 9760 11957 9824
rect 12021 9760 12037 9824
rect 12101 9760 12117 9824
rect 12181 9760 12197 9824
rect 12261 9760 12269 9824
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 8096 9216 8104 9280
rect 8168 9216 8184 9280
rect 8248 9216 8264 9280
rect 8328 9216 8344 9280
rect 8408 9216 8416 9280
rect 8096 8192 8416 9216
rect 8096 8128 8104 8192
rect 8168 8128 8184 8192
rect 8248 8128 8264 8192
rect 8328 8128 8344 8192
rect 8408 8128 8416 8192
rect 8096 7104 8416 8128
rect 8096 7040 8104 7104
rect 8168 7040 8184 7104
rect 8248 7040 8264 7104
rect 8328 7040 8344 7104
rect 8408 7040 8416 7104
rect 8096 6016 8416 7040
rect 9630 6901 9690 9691
rect 11949 8736 12269 9760
rect 15801 19072 16121 19088
rect 15801 19008 15809 19072
rect 15873 19008 15889 19072
rect 15953 19008 15969 19072
rect 16033 19008 16049 19072
rect 16113 19008 16121 19072
rect 15801 17984 16121 19008
rect 15801 17920 15809 17984
rect 15873 17920 15889 17984
rect 15953 17920 15969 17984
rect 16033 17920 16049 17984
rect 16113 17920 16121 17984
rect 15801 16896 16121 17920
rect 15801 16832 15809 16896
rect 15873 16832 15889 16896
rect 15953 16832 15969 16896
rect 16033 16832 16049 16896
rect 16113 16832 16121 16896
rect 15801 15808 16121 16832
rect 15801 15744 15809 15808
rect 15873 15744 15889 15808
rect 15953 15744 15969 15808
rect 16033 15744 16049 15808
rect 16113 15744 16121 15808
rect 15801 14720 16121 15744
rect 15801 14656 15809 14720
rect 15873 14656 15889 14720
rect 15953 14656 15969 14720
rect 16033 14656 16049 14720
rect 16113 14656 16121 14720
rect 15801 13632 16121 14656
rect 15801 13568 15809 13632
rect 15873 13568 15889 13632
rect 15953 13568 15969 13632
rect 16033 13568 16049 13632
rect 16113 13568 16121 13632
rect 15801 12544 16121 13568
rect 15801 12480 15809 12544
rect 15873 12480 15889 12544
rect 15953 12480 15969 12544
rect 16033 12480 16049 12544
rect 16113 12480 16121 12544
rect 15801 11456 16121 12480
rect 15801 11392 15809 11456
rect 15873 11392 15889 11456
rect 15953 11392 15969 11456
rect 16033 11392 16049 11456
rect 16113 11392 16121 11456
rect 15801 10368 16121 11392
rect 15801 10304 15809 10368
rect 15873 10304 15889 10368
rect 15953 10304 15969 10368
rect 16033 10304 16049 10368
rect 16113 10304 16121 10368
rect 15515 9756 15581 9757
rect 15515 9692 15516 9756
rect 15580 9692 15581 9756
rect 15515 9691 15581 9692
rect 11949 8672 11957 8736
rect 12021 8672 12037 8736
rect 12101 8672 12117 8736
rect 12181 8672 12197 8736
rect 12261 8672 12269 8736
rect 11949 7648 12269 8672
rect 12571 8396 12637 8397
rect 12571 8332 12572 8396
rect 12636 8332 12637 8396
rect 12571 8331 12637 8332
rect 11949 7584 11957 7648
rect 12021 7584 12037 7648
rect 12101 7584 12117 7648
rect 12181 7584 12197 7648
rect 12261 7584 12269 7648
rect 9627 6900 9693 6901
rect 9627 6836 9628 6900
rect 9692 6836 9693 6900
rect 9627 6835 9693 6836
rect 8096 5952 8104 6016
rect 8168 5952 8184 6016
rect 8248 5952 8264 6016
rect 8328 5952 8344 6016
rect 8408 5952 8416 6016
rect 8096 4928 8416 5952
rect 8096 4864 8104 4928
rect 8168 4864 8184 4928
rect 8248 4864 8264 4928
rect 8328 4864 8344 4928
rect 8408 4864 8416 4928
rect 8096 3840 8416 4864
rect 8096 3776 8104 3840
rect 8168 3776 8184 3840
rect 8248 3776 8264 3840
rect 8328 3776 8344 3840
rect 8408 3776 8416 3840
rect 8096 2752 8416 3776
rect 8096 2688 8104 2752
rect 8168 2688 8184 2752
rect 8248 2688 8264 2752
rect 8328 2688 8344 2752
rect 8408 2688 8416 2752
rect 8096 1664 8416 2688
rect 8096 1600 8104 1664
rect 8168 1600 8184 1664
rect 8248 1600 8264 1664
rect 8328 1600 8344 1664
rect 8408 1600 8416 1664
rect 8096 576 8416 1600
rect 8096 512 8104 576
rect 8168 512 8184 576
rect 8248 512 8264 576
rect 8328 512 8344 576
rect 8408 512 8416 576
rect 8096 496 8416 512
rect 11949 6560 12269 7584
rect 12574 6901 12634 8331
rect 12571 6900 12637 6901
rect 12571 6836 12572 6900
rect 12636 6836 12637 6900
rect 12571 6835 12637 6836
rect 11949 6496 11957 6560
rect 12021 6496 12037 6560
rect 12101 6496 12117 6560
rect 12181 6496 12197 6560
rect 12261 6496 12269 6560
rect 11949 5472 12269 6496
rect 11949 5408 11957 5472
rect 12021 5408 12037 5472
rect 12101 5408 12117 5472
rect 12181 5408 12197 5472
rect 12261 5408 12269 5472
rect 11949 4384 12269 5408
rect 11949 4320 11957 4384
rect 12021 4320 12037 4384
rect 12101 4320 12117 4384
rect 12181 4320 12197 4384
rect 12261 4320 12269 4384
rect 11949 3296 12269 4320
rect 15518 4045 15578 9691
rect 15801 9280 16121 10304
rect 15801 9216 15809 9280
rect 15873 9216 15889 9280
rect 15953 9216 15969 9280
rect 16033 9216 16049 9280
rect 16113 9216 16121 9280
rect 15801 8192 16121 9216
rect 15801 8128 15809 8192
rect 15873 8128 15889 8192
rect 15953 8128 15969 8192
rect 16033 8128 16049 8192
rect 16113 8128 16121 8192
rect 15801 7104 16121 8128
rect 15801 7040 15809 7104
rect 15873 7040 15889 7104
rect 15953 7040 15969 7104
rect 16033 7040 16049 7104
rect 16113 7040 16121 7104
rect 15801 6016 16121 7040
rect 15801 5952 15809 6016
rect 15873 5952 15889 6016
rect 15953 5952 15969 6016
rect 16033 5952 16049 6016
rect 16113 5952 16121 6016
rect 15801 4928 16121 5952
rect 15801 4864 15809 4928
rect 15873 4864 15889 4928
rect 15953 4864 15969 4928
rect 16033 4864 16049 4928
rect 16113 4864 16121 4928
rect 15515 4044 15581 4045
rect 15515 3980 15516 4044
rect 15580 3980 15581 4044
rect 15515 3979 15581 3980
rect 11949 3232 11957 3296
rect 12021 3232 12037 3296
rect 12101 3232 12117 3296
rect 12181 3232 12197 3296
rect 12261 3232 12269 3296
rect 11949 2208 12269 3232
rect 11949 2144 11957 2208
rect 12021 2144 12037 2208
rect 12101 2144 12117 2208
rect 12181 2144 12197 2208
rect 12261 2144 12269 2208
rect 11949 1120 12269 2144
rect 11949 1056 11957 1120
rect 12021 1056 12037 1120
rect 12101 1056 12117 1120
rect 12181 1056 12197 1120
rect 12261 1056 12269 1120
rect 11949 496 12269 1056
rect 15801 3840 16121 4864
rect 15801 3776 15809 3840
rect 15873 3776 15889 3840
rect 15953 3776 15969 3840
rect 16033 3776 16049 3840
rect 16113 3776 16121 3840
rect 15801 2752 16121 3776
rect 15801 2688 15809 2752
rect 15873 2688 15889 2752
rect 15953 2688 15969 2752
rect 16033 2688 16049 2752
rect 16113 2688 16121 2752
rect 15801 1664 16121 2688
rect 15801 1600 15809 1664
rect 15873 1600 15889 1664
rect 15953 1600 15969 1664
rect 16033 1600 16049 1664
rect 16113 1600 16121 1664
rect 15801 576 16121 1600
rect 15801 512 15809 576
rect 15873 512 15889 576
rect 15953 512 15969 576
rect 16033 512 16049 576
rect 16113 512 16121 576
rect 15801 496 16121 512
rect 19654 18528 19974 19088
rect 19654 18464 19662 18528
rect 19726 18464 19742 18528
rect 19806 18464 19822 18528
rect 19886 18464 19902 18528
rect 19966 18464 19974 18528
rect 19654 17440 19974 18464
rect 19654 17376 19662 17440
rect 19726 17376 19742 17440
rect 19806 17376 19822 17440
rect 19886 17376 19902 17440
rect 19966 17376 19974 17440
rect 19654 16352 19974 17376
rect 19654 16288 19662 16352
rect 19726 16288 19742 16352
rect 19806 16288 19822 16352
rect 19886 16288 19902 16352
rect 19966 16288 19974 16352
rect 19654 15264 19974 16288
rect 19654 15200 19662 15264
rect 19726 15200 19742 15264
rect 19806 15200 19822 15264
rect 19886 15200 19902 15264
rect 19966 15200 19974 15264
rect 19654 14176 19974 15200
rect 19654 14112 19662 14176
rect 19726 14112 19742 14176
rect 19806 14112 19822 14176
rect 19886 14112 19902 14176
rect 19966 14112 19974 14176
rect 19654 13088 19974 14112
rect 19654 13024 19662 13088
rect 19726 13024 19742 13088
rect 19806 13024 19822 13088
rect 19886 13024 19902 13088
rect 19966 13024 19974 13088
rect 19654 12000 19974 13024
rect 19654 11936 19662 12000
rect 19726 11936 19742 12000
rect 19806 11936 19822 12000
rect 19886 11936 19902 12000
rect 19966 11936 19974 12000
rect 19654 10912 19974 11936
rect 19654 10848 19662 10912
rect 19726 10848 19742 10912
rect 19806 10848 19822 10912
rect 19886 10848 19902 10912
rect 19966 10848 19974 10912
rect 19654 9824 19974 10848
rect 19654 9760 19662 9824
rect 19726 9760 19742 9824
rect 19806 9760 19822 9824
rect 19886 9760 19902 9824
rect 19966 9760 19974 9824
rect 19654 8736 19974 9760
rect 19654 8672 19662 8736
rect 19726 8672 19742 8736
rect 19806 8672 19822 8736
rect 19886 8672 19902 8736
rect 19966 8672 19974 8736
rect 19654 7648 19974 8672
rect 19654 7584 19662 7648
rect 19726 7584 19742 7648
rect 19806 7584 19822 7648
rect 19886 7584 19902 7648
rect 19966 7584 19974 7648
rect 19654 6560 19974 7584
rect 19654 6496 19662 6560
rect 19726 6496 19742 6560
rect 19806 6496 19822 6560
rect 19886 6496 19902 6560
rect 19966 6496 19974 6560
rect 19654 5472 19974 6496
rect 19654 5408 19662 5472
rect 19726 5408 19742 5472
rect 19806 5408 19822 5472
rect 19886 5408 19902 5472
rect 19966 5408 19974 5472
rect 19654 4384 19974 5408
rect 19654 4320 19662 4384
rect 19726 4320 19742 4384
rect 19806 4320 19822 4384
rect 19886 4320 19902 4384
rect 19966 4320 19974 4384
rect 19654 3296 19974 4320
rect 19654 3232 19662 3296
rect 19726 3232 19742 3296
rect 19806 3232 19822 3296
rect 19886 3232 19902 3296
rect 19966 3232 19974 3296
rect 19654 2208 19974 3232
rect 19654 2144 19662 2208
rect 19726 2144 19742 2208
rect 19806 2144 19822 2208
rect 19886 2144 19902 2208
rect 19966 2144 19974 2208
rect 19654 1120 19974 2144
rect 19654 1056 19662 1120
rect 19726 1056 19742 1120
rect 19806 1056 19822 1120
rect 19886 1056 19902 1120
rect 19966 1056 19974 1120
rect 19654 496 19974 1056
rect 23506 19072 23826 19088
rect 23506 19008 23514 19072
rect 23578 19008 23594 19072
rect 23658 19008 23674 19072
rect 23738 19008 23754 19072
rect 23818 19008 23826 19072
rect 23506 17984 23826 19008
rect 23506 17920 23514 17984
rect 23578 17920 23594 17984
rect 23658 17920 23674 17984
rect 23738 17920 23754 17984
rect 23818 17920 23826 17984
rect 23506 16896 23826 17920
rect 23506 16832 23514 16896
rect 23578 16832 23594 16896
rect 23658 16832 23674 16896
rect 23738 16832 23754 16896
rect 23818 16832 23826 16896
rect 23506 15808 23826 16832
rect 23506 15744 23514 15808
rect 23578 15744 23594 15808
rect 23658 15744 23674 15808
rect 23738 15744 23754 15808
rect 23818 15744 23826 15808
rect 23506 14720 23826 15744
rect 23506 14656 23514 14720
rect 23578 14656 23594 14720
rect 23658 14656 23674 14720
rect 23738 14656 23754 14720
rect 23818 14656 23826 14720
rect 23506 13632 23826 14656
rect 23506 13568 23514 13632
rect 23578 13568 23594 13632
rect 23658 13568 23674 13632
rect 23738 13568 23754 13632
rect 23818 13568 23826 13632
rect 23506 12544 23826 13568
rect 23506 12480 23514 12544
rect 23578 12480 23594 12544
rect 23658 12480 23674 12544
rect 23738 12480 23754 12544
rect 23818 12480 23826 12544
rect 23506 11456 23826 12480
rect 23506 11392 23514 11456
rect 23578 11392 23594 11456
rect 23658 11392 23674 11456
rect 23738 11392 23754 11456
rect 23818 11392 23826 11456
rect 23506 10368 23826 11392
rect 23506 10304 23514 10368
rect 23578 10304 23594 10368
rect 23658 10304 23674 10368
rect 23738 10304 23754 10368
rect 23818 10304 23826 10368
rect 23506 9280 23826 10304
rect 23506 9216 23514 9280
rect 23578 9216 23594 9280
rect 23658 9216 23674 9280
rect 23738 9216 23754 9280
rect 23818 9216 23826 9280
rect 23506 8192 23826 9216
rect 23506 8128 23514 8192
rect 23578 8128 23594 8192
rect 23658 8128 23674 8192
rect 23738 8128 23754 8192
rect 23818 8128 23826 8192
rect 23506 7104 23826 8128
rect 23506 7040 23514 7104
rect 23578 7040 23594 7104
rect 23658 7040 23674 7104
rect 23738 7040 23754 7104
rect 23818 7040 23826 7104
rect 23506 6016 23826 7040
rect 23506 5952 23514 6016
rect 23578 5952 23594 6016
rect 23658 5952 23674 6016
rect 23738 5952 23754 6016
rect 23818 5952 23826 6016
rect 23506 4928 23826 5952
rect 23506 4864 23514 4928
rect 23578 4864 23594 4928
rect 23658 4864 23674 4928
rect 23738 4864 23754 4928
rect 23818 4864 23826 4928
rect 23506 3840 23826 4864
rect 23506 3776 23514 3840
rect 23578 3776 23594 3840
rect 23658 3776 23674 3840
rect 23738 3776 23754 3840
rect 23818 3776 23826 3840
rect 23506 2752 23826 3776
rect 23506 2688 23514 2752
rect 23578 2688 23594 2752
rect 23658 2688 23674 2752
rect 23738 2688 23754 2752
rect 23818 2688 23826 2752
rect 23506 1664 23826 2688
rect 23506 1600 23514 1664
rect 23578 1600 23594 1664
rect 23658 1600 23674 1664
rect 23738 1600 23754 1664
rect 23818 1600 23826 1664
rect 23506 576 23826 1600
rect 23506 512 23514 576
rect 23578 512 23594 576
rect 23658 512 23674 576
rect 23738 512 23754 576
rect 23818 512 23826 576
rect 23506 496 23826 512
rect 27359 18528 27679 19088
rect 27359 18464 27367 18528
rect 27431 18464 27447 18528
rect 27511 18464 27527 18528
rect 27591 18464 27607 18528
rect 27671 18464 27679 18528
rect 27359 17440 27679 18464
rect 27359 17376 27367 17440
rect 27431 17376 27447 17440
rect 27511 17376 27527 17440
rect 27591 17376 27607 17440
rect 27671 17376 27679 17440
rect 27359 16352 27679 17376
rect 27359 16288 27367 16352
rect 27431 16288 27447 16352
rect 27511 16288 27527 16352
rect 27591 16288 27607 16352
rect 27671 16288 27679 16352
rect 27359 15264 27679 16288
rect 27359 15200 27367 15264
rect 27431 15200 27447 15264
rect 27511 15200 27527 15264
rect 27591 15200 27607 15264
rect 27671 15200 27679 15264
rect 27359 14176 27679 15200
rect 27359 14112 27367 14176
rect 27431 14112 27447 14176
rect 27511 14112 27527 14176
rect 27591 14112 27607 14176
rect 27671 14112 27679 14176
rect 27359 13088 27679 14112
rect 27359 13024 27367 13088
rect 27431 13024 27447 13088
rect 27511 13024 27527 13088
rect 27591 13024 27607 13088
rect 27671 13024 27679 13088
rect 27359 12000 27679 13024
rect 27359 11936 27367 12000
rect 27431 11936 27447 12000
rect 27511 11936 27527 12000
rect 27591 11936 27607 12000
rect 27671 11936 27679 12000
rect 27359 10912 27679 11936
rect 27359 10848 27367 10912
rect 27431 10848 27447 10912
rect 27511 10848 27527 10912
rect 27591 10848 27607 10912
rect 27671 10848 27679 10912
rect 27359 9824 27679 10848
rect 27359 9760 27367 9824
rect 27431 9760 27447 9824
rect 27511 9760 27527 9824
rect 27591 9760 27607 9824
rect 27671 9760 27679 9824
rect 27359 8736 27679 9760
rect 27359 8672 27367 8736
rect 27431 8672 27447 8736
rect 27511 8672 27527 8736
rect 27591 8672 27607 8736
rect 27671 8672 27679 8736
rect 27359 7648 27679 8672
rect 27359 7584 27367 7648
rect 27431 7584 27447 7648
rect 27511 7584 27527 7648
rect 27591 7584 27607 7648
rect 27671 7584 27679 7648
rect 27359 6560 27679 7584
rect 27359 6496 27367 6560
rect 27431 6496 27447 6560
rect 27511 6496 27527 6560
rect 27591 6496 27607 6560
rect 27671 6496 27679 6560
rect 27359 5472 27679 6496
rect 27359 5408 27367 5472
rect 27431 5408 27447 5472
rect 27511 5408 27527 5472
rect 27591 5408 27607 5472
rect 27671 5408 27679 5472
rect 27359 4384 27679 5408
rect 27359 4320 27367 4384
rect 27431 4320 27447 4384
rect 27511 4320 27527 4384
rect 27591 4320 27607 4384
rect 27671 4320 27679 4384
rect 27359 3296 27679 4320
rect 27359 3232 27367 3296
rect 27431 3232 27447 3296
rect 27511 3232 27527 3296
rect 27591 3232 27607 3296
rect 27671 3232 27679 3296
rect 27359 2208 27679 3232
rect 27359 2144 27367 2208
rect 27431 2144 27447 2208
rect 27511 2144 27527 2208
rect 27591 2144 27607 2208
rect 27671 2144 27679 2208
rect 27359 1120 27679 2144
rect 27359 1056 27367 1120
rect 27431 1056 27447 1120
rect 27511 1056 27527 1120
rect 27591 1056 27607 1120
rect 27671 1056 27679 1120
rect 27359 496 27679 1056
rect 31211 19072 31531 19088
rect 31211 19008 31219 19072
rect 31283 19008 31299 19072
rect 31363 19008 31379 19072
rect 31443 19008 31459 19072
rect 31523 19008 31531 19072
rect 31211 17984 31531 19008
rect 31211 17920 31219 17984
rect 31283 17920 31299 17984
rect 31363 17920 31379 17984
rect 31443 17920 31459 17984
rect 31523 17920 31531 17984
rect 31211 16896 31531 17920
rect 31211 16832 31219 16896
rect 31283 16832 31299 16896
rect 31363 16832 31379 16896
rect 31443 16832 31459 16896
rect 31523 16832 31531 16896
rect 31211 15808 31531 16832
rect 31211 15744 31219 15808
rect 31283 15744 31299 15808
rect 31363 15744 31379 15808
rect 31443 15744 31459 15808
rect 31523 15744 31531 15808
rect 31211 14720 31531 15744
rect 31211 14656 31219 14720
rect 31283 14656 31299 14720
rect 31363 14656 31379 14720
rect 31443 14656 31459 14720
rect 31523 14656 31531 14720
rect 31211 13632 31531 14656
rect 31211 13568 31219 13632
rect 31283 13568 31299 13632
rect 31363 13568 31379 13632
rect 31443 13568 31459 13632
rect 31523 13568 31531 13632
rect 31211 12544 31531 13568
rect 31211 12480 31219 12544
rect 31283 12480 31299 12544
rect 31363 12480 31379 12544
rect 31443 12480 31459 12544
rect 31523 12480 31531 12544
rect 31211 11456 31531 12480
rect 31211 11392 31219 11456
rect 31283 11392 31299 11456
rect 31363 11392 31379 11456
rect 31443 11392 31459 11456
rect 31523 11392 31531 11456
rect 31211 10368 31531 11392
rect 31211 10304 31219 10368
rect 31283 10304 31299 10368
rect 31363 10304 31379 10368
rect 31443 10304 31459 10368
rect 31523 10304 31531 10368
rect 31211 9280 31531 10304
rect 31211 9216 31219 9280
rect 31283 9216 31299 9280
rect 31363 9216 31379 9280
rect 31443 9216 31459 9280
rect 31523 9216 31531 9280
rect 31211 8192 31531 9216
rect 31211 8128 31219 8192
rect 31283 8128 31299 8192
rect 31363 8128 31379 8192
rect 31443 8128 31459 8192
rect 31523 8128 31531 8192
rect 31211 7104 31531 8128
rect 31211 7040 31219 7104
rect 31283 7040 31299 7104
rect 31363 7040 31379 7104
rect 31443 7040 31459 7104
rect 31523 7040 31531 7104
rect 31211 6016 31531 7040
rect 31211 5952 31219 6016
rect 31283 5952 31299 6016
rect 31363 5952 31379 6016
rect 31443 5952 31459 6016
rect 31523 5952 31531 6016
rect 31211 4928 31531 5952
rect 31211 4864 31219 4928
rect 31283 4864 31299 4928
rect 31363 4864 31379 4928
rect 31443 4864 31459 4928
rect 31523 4864 31531 4928
rect 31211 3840 31531 4864
rect 31211 3776 31219 3840
rect 31283 3776 31299 3840
rect 31363 3776 31379 3840
rect 31443 3776 31459 3840
rect 31523 3776 31531 3840
rect 31211 2752 31531 3776
rect 31211 2688 31219 2752
rect 31283 2688 31299 2752
rect 31363 2688 31379 2752
rect 31443 2688 31459 2752
rect 31523 2688 31531 2752
rect 31211 1664 31531 2688
rect 31211 1600 31219 1664
rect 31283 1600 31299 1664
rect 31363 1600 31379 1664
rect 31443 1600 31459 1664
rect 31523 1600 31531 1664
rect 31211 576 31531 1600
rect 31211 512 31219 576
rect 31283 512 31299 576
rect 31363 512 31379 576
rect 31443 512 31459 576
rect 31523 512 31531 576
rect 31211 496 31531 512
use sky130_fd_sc_hd__inv_2  _10__3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12512 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__4
timestamp 1701704242
transform -1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__5
timestamp 1701704242
transform 1 0 14076 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__6
timestamp 1701704242
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__7
timestamp 1701704242
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__8
timestamp 1701704242
transform 1 0 17388 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__9
timestamp 1701704242
transform 1 0 17020 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__10
timestamp 1701704242
transform -1 0 16744 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__11
timestamp 1701704242
transform -1 0 16284 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__12
timestamp 1701704242
transform -1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__13
timestamp 1701704242
transform -1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__14
timestamp 1701704242
transform -1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__15
timestamp 1701704242
transform 1 0 10304 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__16
timestamp 1701704242
transform -1 0 12420 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _10__17
timestamp 1701704242
transform -1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12328 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _12_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13156 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _13_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13340 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _14_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13708 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _15_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 14536 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1701704242
transform 1 0 14628 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _17_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15640 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _18_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 15180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _19_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17020 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _20_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 16468 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _21_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 17572 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1701704242
transform -1 0 16560 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _23_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 14076 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _24_
timestamp 1701704242
transform 1 0 14536 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _25_
timestamp 1701704242
transform 1 0 16560 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _26_
timestamp 1701704242
transform 1 0 11500 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _27_
timestamp 1701704242
transform 1 0 13892 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _28_
timestamp 1701704242
transform 1 0 16560 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _29_
timestamp 1701704242
transform 1 0 18308 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _30_
timestamp 1701704242
transform 1 0 18216 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _31_
timestamp 1701704242
transform 1 0 18676 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _32_
timestamp 1701704242
transform 1 0 18308 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _33_
timestamp 1701704242
transform 1 0 16836 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _34_
timestamp 1701704242
transform 1 0 15364 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _35_
timestamp 1701704242
transform 1 0 13524 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _36_
timestamp 1701704242
transform 1 0 10948 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _37_
timestamp 1701704242
transform 1 0 9108 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _38_
timestamp 1701704242
transform 1 0 9016 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _39_
timestamp 1701704242
transform 1 0 13524 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _40_
timestamp 1701704242
transform 1 0 9108 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _41_
timestamp 1701704242
transform 1 0 10212 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _42_
timestamp 1701704242
transform 1 0 16836 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _43_
timestamp 1701704242
transform 1 0 18400 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _44_
timestamp 1701704242
transform 1 0 18676 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _45_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 18676 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _46_
timestamp 1701704242
transform 1 0 19872 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _47_
timestamp 1701704242
transform -1 0 19964 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _48_
timestamp 1701704242
transform 1 0 12788 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _49_
timestamp 1701704242
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _50_
timestamp 1701704242
transform 1 0 18676 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _51_
timestamp 1701704242
transform 1 0 19780 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _52_
timestamp 1701704242
transform 1 0 19688 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _53_
timestamp 1701704242
transform 1 0 20240 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _54_
timestamp 1701704242
transform 1 0 19780 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _55_
timestamp 1701704242
transform 1 0 18676 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _56_
timestamp 1701704242
transform 1 0 16836 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _57_
timestamp 1701704242
transform -1 0 14904 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _58_
timestamp 1701704242
transform 1 0 12420 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _59_
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _60_
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _61_
timestamp 1701704242
transform 1 0 14996 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _62_
timestamp 1701704242
transform 1 0 10580 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _63_
timestamp 1701704242
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _64_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 15916 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_stop pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13892 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net3
timestamp 1701704242
transform 1 0 14076 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_i_stop
timestamp 1701704242
transform -1 0 13340 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net3
timestamp 1701704242
transform -1 0 13708 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_i_stop
timestamp 1701704242
transform 1 0 16560 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net3
timestamp 1701704242
transform 1 0 16376 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__nor2_1  dly_stg1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg2
timestamp 1701704242
transform -1 0 12880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  dly_stg5 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10856 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg6_187
timestamp 1701704242
transform 1 0 12972 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_70
timestamp 1701704242
transform 1 0 12052 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_71
timestamp 1701704242
transform -1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg9_72
timestamp 1701704242
transform 1 0 12328 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_108
timestamp 1701704242
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_109
timestamp 1701704242
transform 1 0 11776 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_110
timestamp 1701704242
transform -1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_111
timestamp 1701704242
transform -1 0 12052 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_112
timestamp 1701704242
transform 1 0 17572 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_113
timestamp 1701704242
transform 1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_114
timestamp 1701704242
transform 1 0 13800 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg10_115
timestamp 1701704242
transform -1 0 13708 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_154
timestamp 1701704242
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_155
timestamp 1701704242
transform -1 0 13156 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg11_156
timestamp 1701704242
transform 1 0 13616 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_73
timestamp 1701704242
transform 1 0 13800 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_74
timestamp 1701704242
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_75
timestamp 1701704242
transform -1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  dly_stg12_76
timestamp 1701704242
transform -1 0 14444 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  dly_strt_inv_chain_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1701704242
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1701704242
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1701704242
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1701704242
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1701704242
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1701704242
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1701704242
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1701704242
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1701704242
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1701704242
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1701704242
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1701704242
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1701704242
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1701704242
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1701704242
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1701704242
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1701704242
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1701704242
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1701704242
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1701704242
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1701704242
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1701704242
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_321 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_329
timestamp 1701704242
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1701704242
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1701704242
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1701704242
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1701704242
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1701704242
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1701704242
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1701704242
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1701704242
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1701704242
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1701704242
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1701704242
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1701704242
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1701704242
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1701704242
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1701704242
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1701704242
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1701704242
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1701704242
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1701704242
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1701704242
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1701704242
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 1701704242
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1701704242
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1701704242
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1701704242
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1701704242
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1701704242
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1701704242
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1701704242
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1701704242
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1701704242
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1701704242
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1701704242
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1701704242
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1701704242
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1701704242
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1701704242
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1701704242
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1701704242
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1701704242
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1701704242
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1701704242
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1701704242
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1701704242
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1701704242
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1701704242
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1701704242
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1701704242
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1701704242
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1701704242
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1701704242
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1701704242
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1701704242
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1701704242
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1701704242
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1701704242
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1701704242
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1701704242
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1701704242
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1701704242
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1701704242
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1701704242
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1701704242
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1701704242
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1701704242
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1701704242
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1701704242
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 1701704242
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1701704242
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1701704242
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1701704242
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1701704242
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1701704242
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1701704242
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1701704242
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1701704242
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1701704242
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1701704242
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1701704242
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1701704242
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1701704242
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1701704242
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1701704242
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1701704242
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1701704242
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1701704242
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1701704242
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1701704242
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1701704242
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1701704242
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1701704242
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_321
timestamp 1701704242
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_329
timestamp 1701704242
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1701704242
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1701704242
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1701704242
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1701704242
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1701704242
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1701704242
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1701704242
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1701704242
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1701704242
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1701704242
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1701704242
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1701704242
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1701704242
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1701704242
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1701704242
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1701704242
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1701704242
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1701704242
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1701704242
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1701704242
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1701704242
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1701704242
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1701704242
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1701704242
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 1701704242
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1701704242
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1701704242
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1701704242
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1701704242
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1701704242
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1701704242
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1701704242
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1701704242
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1701704242
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1701704242
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1701704242
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1701704242
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1701704242
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1701704242
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1701704242
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1701704242
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1701704242
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1701704242
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1701704242
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1701704242
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1701704242
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1701704242
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1701704242
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1701704242
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1701704242
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_321
timestamp 1701704242
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_329
timestamp 1701704242
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1701704242
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1701704242
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1701704242
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1701704242
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1701704242
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1701704242
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1701704242
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1701704242
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1701704242
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1701704242
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1701704242
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1701704242
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1701704242
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1701704242
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1701704242
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1701704242
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1701704242
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1701704242
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1701704242
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1701704242
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1701704242
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1701704242
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1701704242
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1701704242
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1701704242
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_329
timestamp 1701704242
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1701704242
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1701704242
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1701704242
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1701704242
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1701704242
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1701704242
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1701704242
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1701704242
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1701704242
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1701704242
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1701704242
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1701704242
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1701704242
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1701704242
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1701704242
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1701704242
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1701704242
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1701704242
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1701704242
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1701704242
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1701704242
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1701704242
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1701704242
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1701704242
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1701704242
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1701704242
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_321
timestamp 1701704242
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_329
timestamp 1701704242
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1701704242
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1701704242
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1701704242
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1701704242
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1701704242
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1701704242
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_119
timestamp 1701704242
transform 1 0 11500 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_125
timestamp 1701704242
transform 1 0 12052 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_129 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_137
timestamp 1701704242
transform 1 0 13156 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_143
timestamp 1701704242
transform 1 0 13708 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_147
timestamp 1701704242
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1701704242
transform 1 0 15180 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1701704242
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1701704242
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1701704242
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1701704242
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1701704242
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1701704242
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1701704242
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1701704242
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1701704242
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1701704242
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1701704242
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1701704242
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1701704242
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1701704242
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1701704242
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1701704242
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1701704242
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_329
timestamp 1701704242
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1701704242
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1701704242
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1701704242
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1701704242
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1701704242
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1701704242
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_109
timestamp 1701704242
transform 1 0 10580 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1701704242
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_150
timestamp 1701704242
transform 1 0 14352 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_154
timestamp 1701704242
transform 1 0 14720 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_161
timestamp 1701704242
transform 1 0 15364 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_171
timestamp 1701704242
transform 1 0 16284 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_183
timestamp 1701704242
transform 1 0 17388 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1701704242
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1701704242
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1701704242
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1701704242
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1701704242
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1701704242
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1701704242
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1701704242
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1701704242
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1701704242
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1701704242
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1701704242
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1701704242
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1701704242
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_321
timestamp 1701704242
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 1701704242
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1701704242
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1701704242
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1701704242
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1701704242
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1701704242
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1701704242
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_93
timestamp 1701704242
transform 1 0 9108 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_101
timestamp 1701704242
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_128
timestamp 1701704242
transform 1 0 12328 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_156
timestamp 1701704242
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_160
timestamp 1701704242
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_175
timestamp 1701704242
transform 1 0 16652 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_197
timestamp 1701704242
transform 1 0 18676 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_209
timestamp 1701704242
transform 1 0 19780 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp 1701704242
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1701704242
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1701704242
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1701704242
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1701704242
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1701704242
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1701704242
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1701704242
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1701704242
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1701704242
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1701704242
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_329
timestamp 1701704242
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1701704242
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1701704242
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1701704242
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1701704242
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1701704242
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1701704242
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1701704242
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1701704242
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_97
timestamp 1701704242
transform 1 0 9476 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_135
timestamp 1701704242
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_157
timestamp 1701704242
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1701704242
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_212
timestamp 1701704242
transform 1 0 20056 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_224
timestamp 1701704242
transform 1 0 21160 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_236
timestamp 1701704242
transform 1 0 22264 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_248
timestamp 1701704242
transform 1 0 23368 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1701704242
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1701704242
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1701704242
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1701704242
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1701704242
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1701704242
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1701704242
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_321
timestamp 1701704242
transform 1 0 30084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_329
timestamp 1701704242
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1701704242
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1701704242
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1701704242
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1701704242
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1701704242
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1701704242
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_81
timestamp 1701704242
transform 1 0 8004 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1701704242
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_172
timestamp 1701704242
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_218
timestamp 1701704242
transform 1 0 20608 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1701704242
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1701704242
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1701704242
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1701704242
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1701704242
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1701704242
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1701704242
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1701704242
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1701704242
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1701704242
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_329
timestamp 1701704242
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1701704242
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1701704242
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1701704242
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1701704242
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_77
timestamp 1701704242
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1701704242
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_222
timestamp 1701704242
transform 1 0 20976 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_234
timestamp 1701704242
transform 1 0 22080 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_246
timestamp 1701704242
transform 1 0 23184 0 1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1701704242
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1701704242
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1701704242
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1701704242
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1701704242
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1701704242
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1701704242
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_321
timestamp 1701704242
transform 1 0 30084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_329
timestamp 1701704242
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1701704242
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1701704242
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1701704242
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_69
timestamp 1701704242
transform 1 0 6900 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_108
timestamp 1701704242
transform 1 0 10488 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_119
timestamp 1701704242
transform 1 0 11500 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_143
timestamp 1701704242
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1701704242
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_231
timestamp 1701704242
transform 1 0 21804 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_243
timestamp 1701704242
transform 1 0 22908 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_255
timestamp 1701704242
transform 1 0 24012 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_267
timestamp 1701704242
transform 1 0 25116 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1701704242
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1701704242
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1701704242
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1701704242
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1701704242
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_329
timestamp 1701704242
transform 1 0 30820 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1701704242
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1701704242
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1701704242
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1701704242
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1701704242
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_77
timestamp 1701704242
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1701704242
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_115
timestamp 1701704242
transform 1 0 11132 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1701704242
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_167
timestamp 1701704242
transform 1 0 15916 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1701704242
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1701704242
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1701704242
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1701704242
transform 1 0 23092 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1701704242
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1701704242
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1701704242
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1701704242
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1701704242
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1701704242
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1701704242
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1701704242
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1701704242
transform 1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_329
timestamp 1701704242
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1701704242
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1701704242
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1701704242
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1701704242
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1701704242
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1701704242
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_81
timestamp 1701704242
transform 1 0 8004 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_87
timestamp 1701704242
transform 1 0 8556 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_140
timestamp 1701704242
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1701704242
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1701704242
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_218
timestamp 1701704242
transform 1 0 20608 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1701704242
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1701704242
transform 1 0 22356 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1701704242
transform 1 0 23460 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1701704242
transform 1 0 24564 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1701704242
transform 1 0 25668 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1701704242
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1701704242
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1701704242
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1701704242
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1701704242
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_329
timestamp 1701704242
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1701704242
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1701704242
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1701704242
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1701704242
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1701704242
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1701704242
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1701704242
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1701704242
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_93
timestamp 1701704242
transform 1 0 9108 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_127
timestamp 1701704242
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1701704242
transform 1 0 13524 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_157
timestamp 1701704242
transform 1 0 14996 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_164
timestamp 1701704242
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_171
timestamp 1701704242
transform 1 0 16284 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_212
timestamp 1701704242
transform 1 0 20056 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_224
timestamp 1701704242
transform 1 0 21160 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_236
timestamp 1701704242
transform 1 0 22264 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 1701704242
transform 1 0 23368 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1701704242
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1701704242
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1701704242
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1701704242
transform 1 0 27140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1701704242
transform 1 0 28244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1701704242
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1701704242
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_321
timestamp 1701704242
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_329
timestamp 1701704242
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1701704242
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1701704242
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1701704242
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1701704242
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1701704242
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1701704242
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1701704242
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_105
timestamp 1701704242
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_123
timestamp 1701704242
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_150
timestamp 1701704242
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_175
timestamp 1701704242
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_193
timestamp 1701704242
transform 1 0 18308 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_216
timestamp 1701704242
transform 1 0 20424 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1701704242
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1701704242
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1701704242
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1701704242
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1701704242
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1701704242
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1701704242
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1701704242
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1701704242
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1701704242
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_329
timestamp 1701704242
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1701704242
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1701704242
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1701704242
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1701704242
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1701704242
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1701704242
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1701704242
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1701704242
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1701704242
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1701704242
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1701704242
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_109
timestamp 1701704242
transform 1 0 10580 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1701704242
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1701704242
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_152
timestamp 1701704242
transform 1 0 14536 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_156
timestamp 1701704242
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_163
timestamp 1701704242
transform 1 0 15548 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_179
timestamp 1701704242
transform 1 0 17020 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_188
timestamp 1701704242
transform 1 0 17848 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_213
timestamp 1701704242
transform 1 0 20148 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_225
timestamp 1701704242
transform 1 0 21252 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_237
timestamp 1701704242
transform 1 0 22356 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1701704242
transform 1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1701704242
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1701704242
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1701704242
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1701704242
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1701704242
transform 1 0 28244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1701704242
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1701704242
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_321
timestamp 1701704242
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_329
timestamp 1701704242
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1701704242
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1701704242
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1701704242
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1701704242
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1701704242
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1701704242
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1701704242
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1701704242
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1701704242
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1701704242
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1701704242
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1701704242
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1701704242
transform 1 0 10948 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_121
timestamp 1701704242
transform 1 0 11684 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_131
timestamp 1701704242
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_138
timestamp 1701704242
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_143
timestamp 1701704242
transform 1 0 13708 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_163
timestamp 1701704242
transform 1 0 15548 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1701704242
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1701704242
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_190
timestamp 1701704242
transform 1 0 18032 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_202
timestamp 1701704242
transform 1 0 19136 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_211
timestamp 1701704242
transform 1 0 19964 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1701704242
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1701704242
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1701704242
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1701704242
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1701704242
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1701704242
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1701704242
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1701704242
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1701704242
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1701704242
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1701704242
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_329
timestamp 1701704242
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1701704242
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1701704242
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1701704242
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1701704242
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1701704242
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1701704242
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1701704242
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1701704242
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1701704242
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1701704242
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1701704242
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1701704242
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1701704242
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1701704242
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1701704242
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1701704242
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1701704242
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1701704242
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1701704242
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1701704242
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1701704242
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1701704242
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1701704242
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1701704242
transform 1 0 20884 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1701704242
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1701704242
transform 1 0 23092 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1701704242
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1701704242
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1701704242
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1701704242
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1701704242
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1701704242
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1701704242
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1701704242
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_321
timestamp 1701704242
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_329
timestamp 1701704242
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1701704242
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1701704242
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1701704242
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1701704242
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1701704242
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1701704242
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1701704242
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1701704242
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1701704242
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1701704242
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1701704242
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1701704242
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1701704242
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1701704242
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1701704242
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1701704242
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1701704242
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1701704242
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1701704242
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1701704242
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1701704242
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1701704242
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1701704242
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1701704242
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1701704242
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1701704242
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1701704242
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1701704242
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1701704242
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1701704242
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1701704242
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1701704242
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1701704242
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1701704242
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_329
timestamp 1701704242
transform 1 0 30820 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1701704242
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1701704242
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1701704242
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1701704242
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1701704242
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1701704242
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1701704242
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1701704242
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1701704242
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1701704242
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1701704242
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1701704242
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1701704242
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1701704242
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1701704242
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1701704242
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1701704242
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1701704242
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1701704242
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1701704242
transform 1 0 17940 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1701704242
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1701704242
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1701704242
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1701704242
transform 1 0 20884 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1701704242
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1701704242
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1701704242
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1701704242
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1701704242
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1701704242
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1701704242
transform 1 0 27140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1701704242
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1701704242
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1701704242
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_321
timestamp 1701704242
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_329
timestamp 1701704242
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1701704242
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1701704242
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1701704242
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1701704242
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1701704242
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1701704242
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1701704242
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1701704242
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1701704242
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1701704242
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1701704242
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1701704242
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1701704242
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1701704242
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1701704242
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1701704242
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1701704242
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1701704242
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1701704242
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1701704242
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1701704242
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1701704242
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1701704242
transform 1 0 20516 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1701704242
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1701704242
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1701704242
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1701704242
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1701704242
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1701704242
transform 1 0 25668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1701704242
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1701704242
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1701704242
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1701704242
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1701704242
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_329
timestamp 1701704242
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1701704242
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1701704242
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1701704242
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1701704242
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1701704242
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1701704242
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1701704242
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1701704242
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1701704242
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1701704242
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1701704242
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1701704242
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1701704242
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1701704242
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1701704242
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1701704242
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1701704242
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1701704242
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1701704242
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1701704242
transform 1 0 17940 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1701704242
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1701704242
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1701704242
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1701704242
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1701704242
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1701704242
transform 1 0 23092 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1701704242
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1701704242
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1701704242
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1701704242
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1701704242
transform 1 0 27140 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1701704242
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1701704242
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1701704242
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1701704242
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_329
timestamp 1701704242
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1701704242
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1701704242
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1701704242
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1701704242
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1701704242
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1701704242
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1701704242
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1701704242
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1701704242
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1701704242
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1701704242
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1701704242
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1701704242
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1701704242
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1701704242
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1701704242
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1701704242
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1701704242
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1701704242
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1701704242
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1701704242
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1701704242
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1701704242
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1701704242
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1701704242
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1701704242
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1701704242
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1701704242
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1701704242
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1701704242
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1701704242
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1701704242
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1701704242
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1701704242
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_329
timestamp 1701704242
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1701704242
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1701704242
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1701704242
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1701704242
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1701704242
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1701704242
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1701704242
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1701704242
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1701704242
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1701704242
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1701704242
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1701704242
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1701704242
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1701704242
transform 1 0 12788 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1701704242
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1701704242
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1701704242
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1701704242
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1701704242
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1701704242
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1701704242
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1701704242
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1701704242
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1701704242
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1701704242
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1701704242
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1701704242
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1701704242
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1701704242
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1701704242
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1701704242
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1701704242
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1701704242
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1701704242
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_321
timestamp 1701704242
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_329
timestamp 1701704242
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1701704242
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1701704242
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1701704242
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1701704242
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1701704242
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1701704242
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1701704242
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1701704242
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1701704242
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1701704242
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1701704242
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1701704242
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1701704242
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1701704242
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1701704242
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1701704242
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1701704242
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1701704242
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1701704242
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1701704242
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1701704242
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1701704242
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1701704242
transform 1 0 20516 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1701704242
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1701704242
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1701704242
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1701704242
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1701704242
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1701704242
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1701704242
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1701704242
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1701704242
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1701704242
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1701704242
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_329
timestamp 1701704242
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1701704242
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1701704242
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1701704242
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1701704242
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1701704242
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1701704242
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1701704242
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1701704242
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1701704242
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1701704242
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1701704242
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1701704242
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1701704242
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1701704242
transform 1 0 12788 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1701704242
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1701704242
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1701704242
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1701704242
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1701704242
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1701704242
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1701704242
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1701704242
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1701704242
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1701704242
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1701704242
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1701704242
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1701704242
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1701704242
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1701704242
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1701704242
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1701704242
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1701704242
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1701704242
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1701704242
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_321
timestamp 1701704242
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_329
timestamp 1701704242
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1701704242
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1701704242
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1701704242
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1701704242
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1701704242
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1701704242
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1701704242
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1701704242
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1701704242
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1701704242
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1701704242
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1701704242
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1701704242
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1701704242
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1701704242
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1701704242
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1701704242
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1701704242
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1701704242
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1701704242
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1701704242
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1701704242
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1701704242
transform 1 0 20516 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1701704242
transform 1 0 21068 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1701704242
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1701704242
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1701704242
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1701704242
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1701704242
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1701704242
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1701704242
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1701704242
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1701704242
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1701704242
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_329
timestamp 1701704242
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1701704242
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1701704242
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1701704242
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1701704242
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1701704242
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1701704242
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1701704242
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1701704242
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1701704242
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1701704242
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1701704242
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1701704242
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1701704242
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1701704242
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1701704242
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1701704242
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1701704242
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1701704242
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1701704242
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1701704242
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1701704242
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1701704242
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1701704242
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1701704242
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1701704242
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1701704242
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1701704242
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1701704242
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1701704242
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1701704242
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1701704242
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1701704242
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1701704242
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1701704242
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1701704242
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_329
timestamp 1701704242
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1701704242
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1701704242
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 1701704242
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1701704242
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1701704242
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1701704242
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1701704242
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1701704242
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1701704242
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1701704242
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1701704242
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1701704242
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1701704242
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1701704242
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_137
timestamp 1701704242
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_141
timestamp 1701704242
transform 1 0 13524 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_145
timestamp 1701704242
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_157
timestamp 1701704242
transform 1 0 14996 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1701704242
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1701704242
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1701704242
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_193
timestamp 1701704242
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_197
timestamp 1701704242
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_209
timestamp 1701704242
transform 1 0 19780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1701704242
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1701704242
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1701704242
transform 1 0 22356 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_249
timestamp 1701704242
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_253
timestamp 1701704242
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_265
timestamp 1701704242
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1701704242
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1701704242
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1701704242
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_305
timestamp 1701704242
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_309
timestamp 1701704242
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_321
timestamp 1701704242
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_329
timestamp 1701704242
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[1\].dly_stg3
timestamp 1701704242
transform 1 0 15732 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_18
timestamp 1701704242
transform -1 0 16284 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_19
timestamp 1701704242
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_20
timestamp 1701704242
transform -1 0 16192 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[1\].dly_stg4_21
timestamp 1701704242
transform 1 0 17204 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[2\].dly_stg3
timestamp 1701704242
transform 1 0 15640 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_22
timestamp 1701704242
transform 1 0 19780 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_23
timestamp 1701704242
transform -1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_24
timestamp 1701704242
transform -1 0 17848 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[2\].dly_stg4_25
timestamp 1701704242
transform 1 0 19504 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[3\].dly_stg3
timestamp 1701704242
transform -1 0 19504 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_26
timestamp 1701704242
transform -1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_27
timestamp 1701704242
transform 1 0 18124 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_28
timestamp 1701704242
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[3\].dly_stg4_29
timestamp 1701704242
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[4\].dly_stg3
timestamp 1701704242
transform -1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_30
timestamp 1701704242
transform -1 0 15640 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_31
timestamp 1701704242
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_32
timestamp 1701704242
transform 1 0 18216 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[4\].dly_stg4_33
timestamp 1701704242
transform 1 0 19780 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[5\].dly_stg3
timestamp 1701704242
transform -1 0 20424 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_34
timestamp 1701704242
transform -1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_35
timestamp 1701704242
transform -1 0 18676 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_36
timestamp 1701704242
transform 1 0 15456 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[5\].dly_stg4_37
timestamp 1701704242
transform 1 0 20332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[6\].dly_stg3
timestamp 1701704242
transform 1 0 13432 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_38
timestamp 1701704242
transform -1 0 13800 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_39
timestamp 1701704242
transform -1 0 15088 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_40
timestamp 1701704242
transform -1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[6\].dly_stg4_41
timestamp 1701704242
transform 1 0 20700 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[7\].dly_stg3
timestamp 1701704242
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_42
timestamp 1701704242
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_43
timestamp 1701704242
transform -1 0 13432 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_44
timestamp 1701704242
transform 1 0 12880 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[7\].dly_stg4_45
timestamp 1701704242
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[8\].dly_stg3
timestamp 1701704242
transform -1 0 12604 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_46
timestamp 1701704242
transform -1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_47
timestamp 1701704242
transform 1 0 13156 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_48
timestamp 1701704242
transform -1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[8\].dly_stg4_49
timestamp 1701704242
transform -1 0 14076 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[9\].dly_stg3
timestamp 1701704242
transform -1 0 13156 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_50
timestamp 1701704242
transform 1 0 13248 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_51
timestamp 1701704242
transform 1 0 11500 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_52
timestamp 1701704242
transform 1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[9\].dly_stg4_53
timestamp 1701704242
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[10\].dly_stg3
timestamp 1701704242
transform 1 0 9844 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_54
timestamp 1701704242
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_55
timestamp 1701704242
transform 1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_56
timestamp 1701704242
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[10\].dly_stg4_57
timestamp 1701704242
transform -1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[11\].dly_stg3
timestamp 1701704242
transform -1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_58
timestamp 1701704242
transform -1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_59
timestamp 1701704242
transform 1 0 12696 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_60
timestamp 1701704242
transform 1 0 12236 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[11\].dly_stg4_61
timestamp 1701704242
transform -1 0 8280 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[12\].dly_stg3
timestamp 1701704242
transform 1 0 8464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_62
timestamp 1701704242
transform -1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_63
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_64
timestamp 1701704242
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[12\].dly_stg4_65
timestamp 1701704242
transform -1 0 11776 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[13\].dly_stg3
timestamp 1701704242
transform 1 0 8188 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_66
timestamp 1701704242
transform 1 0 12052 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_67
timestamp 1701704242
transform 1 0 10672 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_68
timestamp 1701704242
transform 1 0 11776 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[13\].dly_stg4_69
timestamp 1701704242
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  g_dly_chain\[14\].dly_stg3
timestamp 1701704242
transform 1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain\[14\].dly_stg4_186
timestamp 1701704242
transform 1 0 11224 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_116
timestamp 1701704242
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_117
timestamp 1701704242
transform -1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_118
timestamp 1701704242
transform -1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_119
timestamp 1701704242
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_120
timestamp 1701704242
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg7_121
timestamp 1701704242
transform -1 0 16928 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[0\].dly_stg8_157
timestamp 1701704242
transform 1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_77
timestamp 1701704242
transform 1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_78
timestamp 1701704242
transform -1 0 18308 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_79
timestamp 1701704242
transform -1 0 16652 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_80
timestamp 1701704242
transform 1 0 19504 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_81
timestamp 1701704242
transform 1 0 17848 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg7_82
timestamp 1701704242
transform -1 0 16468 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[1\].dly_stg8_122
timestamp 1701704242
transform 1 0 16284 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_158
timestamp 1701704242
transform 1 0 19780 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_159
timestamp 1701704242
transform 1 0 16560 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_160
timestamp 1701704242
transform 1 0 17756 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_161
timestamp 1701704242
transform 1 0 20792 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_162
timestamp 1701704242
transform -1 0 20608 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg7_163
timestamp 1701704242
transform 1 0 17296 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[2\].dly_stg8_83
timestamp 1701704242
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_123
timestamp 1701704242
transform 1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_124
timestamp 1701704242
transform 1 0 17940 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_125
timestamp 1701704242
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_126
timestamp 1701704242
transform -1 0 17020 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_127
timestamp 1701704242
transform 1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg7_128
timestamp 1701704242
transform 1 0 16744 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[3\].dly_stg8_164
timestamp 1701704242
transform -1 0 20332 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_84
timestamp 1701704242
transform 1 0 19504 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_85
timestamp 1701704242
transform 1 0 15088 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_86
timestamp 1701704242
transform 1 0 21252 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_87
timestamp 1701704242
transform -1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_88
timestamp 1701704242
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg7_89
timestamp 1701704242
transform 1 0 17572 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[4\].dly_stg8_129
timestamp 1701704242
transform 1 0 21528 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_165
timestamp 1701704242
transform 1 0 20424 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_166
timestamp 1701704242
transform -1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_167
timestamp 1701704242
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_168
timestamp 1701704242
transform -1 0 14720 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_169
timestamp 1701704242
transform -1 0 16652 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg7_170
timestamp 1701704242
transform -1 0 14260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[5\].dly_stg8_90
timestamp 1701704242
transform -1 0 16376 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_130
timestamp 1701704242
transform 1 0 15732 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_131
timestamp 1701704242
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_132
timestamp 1701704242
transform -1 0 14536 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_133
timestamp 1701704242
transform -1 0 11224 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_134
timestamp 1701704242
transform -1 0 14076 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg7_135
timestamp 1701704242
transform 1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[6\].dly_stg8_171
timestamp 1701704242
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_91
timestamp 1701704242
transform 1 0 14076 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_92
timestamp 1701704242
transform -1 0 13340 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_93
timestamp 1701704242
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_94
timestamp 1701704242
transform -1 0 10948 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_95
timestamp 1701704242
transform -1 0 14076 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg7_96
timestamp 1701704242
transform -1 0 12880 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[7\].dly_stg8_136
timestamp 1701704242
transform -1 0 13432 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_172
timestamp 1701704242
transform -1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_173
timestamp 1701704242
transform 1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_174
timestamp 1701704242
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_175
timestamp 1701704242
transform 1 0 11224 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_176
timestamp 1701704242
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg7_177
timestamp 1701704242
transform 1 0 9292 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[8\].dly_stg8_97
timestamp 1701704242
transform -1 0 12328 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_137
timestamp 1701704242
transform -1 0 8832 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_138
timestamp 1701704242
transform -1 0 7912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_139
timestamp 1701704242
transform 1 0 7912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_140
timestamp 1701704242
transform 1 0 11776 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_141
timestamp 1701704242
transform 1 0 12420 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg7_142
timestamp 1701704242
transform -1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[9\].dly_stg8_178
timestamp 1701704242
transform 1 0 12788 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_98
timestamp 1701704242
transform -1 0 8924 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_99
timestamp 1701704242
transform 1 0 10580 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_100
timestamp 1701704242
transform 1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_101
timestamp 1701704242
transform -1 0 11960 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_102
timestamp 1701704242
transform 1 0 11960 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg7_103
timestamp 1701704242
transform 1 0 9568 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[10\].dly_stg8_143
timestamp 1701704242
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_179
timestamp 1701704242
transform 1 0 11592 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_180
timestamp 1701704242
transform 1 0 8832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_181
timestamp 1701704242
transform -1 0 8740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_182
timestamp 1701704242
transform 1 0 11500 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_183
timestamp 1701704242
transform -1 0 8832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg7_184
timestamp 1701704242
transform 1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[11\].dly_stg8_104
timestamp 1701704242
transform -1 0 9016 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_144
timestamp 1701704242
transform -1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_145
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_146
timestamp 1701704242
transform 1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_147
timestamp 1701704242
transform 1 0 9476 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_148
timestamp 1701704242
transform -1 0 10120 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg7_149
timestamp 1701704242
transform -1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[12\].dly_stg8_185
timestamp 1701704242
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_105
timestamp 1701704242
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg7_106
timestamp 1701704242
transform -1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  g_dly_chain_interleave\[13\].dly_stg7_107 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11224 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_150
timestamp 1701704242
transform 1 0 9936 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_151
timestamp 1701704242
transform 1 0 12328 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_152
timestamp 1701704242
transform 1 0 12052 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  g_dly_chain_interleave\[13\].dly_stg8_153
timestamp 1701704242
transform -1 0 9936 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[0\].dly_stp_1
timestamp 1701704242
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_stp\[1\].dly_stp_2
timestamp 1701704242
transform -1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[1\].inv_chain
timestamp 1701704242
transform -1 0 13248 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  g_dly_strt\[2\].inv_chain
timestamp 1701704242
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1701704242
transform -1 0 13892 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1701704242
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1701704242
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1701704242
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1701704242
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1701704242
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1701704242
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1701704242
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1701704242
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1701704242
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1701704242
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1701704242
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1701704242
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1701704242
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1701704242
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1701704242
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1701704242
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1701704242
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1701704242
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1701704242
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1701704242
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1701704242
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1701704242
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1701704242
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1701704242
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1701704242
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1701704242
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1701704242
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1701704242
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1701704242
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1701704242
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1701704242
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1701704242
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1701704242
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1701704242
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1701704242
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1701704242
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 1701704242
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 1701704242
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 1701704242
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 1701704242
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 1701704242
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 1701704242
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 1701704242
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 1701704242
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 1701704242
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 1701704242
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 1701704242
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 1701704242
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 1701704242
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 1701704242
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 1701704242
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 1701704242
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 1701704242
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 1701704242
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 1701704242
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 1701704242
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 1701704242
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 1701704242
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1701704242
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 1701704242
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1701704242
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1701704242
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1701704242
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1701704242
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1701704242
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1701704242
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1701704242
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1701704242
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 1701704242
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 1701704242
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 1701704242
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 1701704242
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 1701704242
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 1701704242
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 1701704242
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 1701704242
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 1701704242
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 1701704242
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 1701704242
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 1701704242
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 1701704242
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 1701704242
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 1701704242
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1701704242
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 1701704242
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 1701704242
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1701704242
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 1701704242
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1701704242
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1701704242
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1701704242
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1701704242
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1701704242
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1701704242
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1701704242
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1701704242
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1701704242
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1701704242
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1701704242
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1701704242
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1701704242
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1701704242
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1701704242
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1701704242
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1701704242
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1701704242
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1701704242
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1701704242
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1701704242
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1701704242
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1701704242
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1701704242
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1701704242
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1701704242
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1701704242
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1701704242
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1701704242
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1701704242
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1701704242
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1701704242
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1701704242
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1701704242
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1701704242
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1701704242
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1701704242
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1701704242
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1701704242
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 1701704242
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 1701704242
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1701704242
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1701704242
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 1701704242
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 1701704242
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 1701704242
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1701704242
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1701704242
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 1701704242
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 1701704242
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 1701704242
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 1701704242
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 1701704242
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 1701704242
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 1701704242
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 1701704242
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 1701704242
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 1701704242
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 1701704242
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 1701704242
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 1701704242
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 1701704242
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 1701704242
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 1701704242
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 1701704242
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 1701704242
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 1701704242
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 1701704242
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 1701704242
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 1701704242
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 1701704242
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 1701704242
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 1701704242
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 1701704242
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 1701704242
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 1701704242
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 1701704242
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 1701704242
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 1701704242
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 1701704242
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 1701704242
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 1701704242
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 1701704242
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 1701704242
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 1701704242
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 1701704242
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 1701704242
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 1701704242
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 1701704242
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 1701704242
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 1701704242
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 1701704242
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 1701704242
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 1701704242
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 1701704242
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1701704242
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 8096 496 8416 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15801 496 16121 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23506 496 23826 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 31211 496 31531 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4244 496 4564 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11949 496 12269 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19654 496 19974 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 27359 496 27679 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 13542 19600 13598 20000 0 FreeSans 224 90 0 0 i_start
port 2 nsew signal input
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 i_stop
port 3 nsew signal input
flabel metal2 s 18694 19600 18750 20000 0 FreeSans 224 90 0 0 o_result_ctr[0]
port 4 nsew signal tristate
flabel metal2 s 19982 19600 20038 20000 0 FreeSans 224 90 0 0 o_result_ctr[1]
port 5 nsew signal tristate
flabel metal2 s 19338 19600 19394 20000 0 FreeSans 224 90 0 0 o_result_ctr[2]
port 6 nsew signal tristate
flabel metal2 s 12898 19600 12954 20000 0 FreeSans 224 90 0 0 o_result_ring[0]
port 7 nsew signal tristate
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 o_result_ring[10]
port 8 nsew signal tristate
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 o_result_ring[11]
port 9 nsew signal tristate
flabel metal3 s 0 8848 400 8968 0 FreeSans 480 0 0 0 o_result_ring[12]
port 10 nsew signal tristate
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 o_result_ring[13]
port 11 nsew signal tristate
flabel metal3 s 0 9528 400 9648 0 FreeSans 480 0 0 0 o_result_ring[14]
port 12 nsew signal tristate
flabel metal3 s 0 10208 400 10328 0 FreeSans 480 0 0 0 o_result_ring[15]
port 13 nsew signal tristate
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 o_result_ring[1]
port 14 nsew signal tristate
flabel metal2 s 18050 19600 18106 20000 0 FreeSans 224 90 0 0 o_result_ring[2]
port 15 nsew signal tristate
flabel metal3 s 31600 10208 32000 10328 0 FreeSans 480 0 0 0 o_result_ring[3]
port 16 nsew signal tristate
flabel metal3 s 31600 9528 32000 9648 0 FreeSans 480 0 0 0 o_result_ring[4]
port 17 nsew signal tristate
flabel metal3 s 31600 8848 32000 8968 0 FreeSans 480 0 0 0 o_result_ring[5]
port 18 nsew signal tristate
flabel metal2 s 19982 0 20038 400 0 FreeSans 224 90 0 0 o_result_ring[6]
port 19 nsew signal tristate
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 o_result_ring[7]
port 20 nsew signal tristate
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 o_result_ring[8]
port 21 nsew signal tristate
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 o_result_ring[9]
port 22 nsew signal tristate
rlabel via1 16041 19040 16041 19040 0 VGND
rlabel metal1 15962 18496 15962 18496 0 VPWR
rlabel metal2 14674 12070 14674 12070 0 _00_
rlabel metal1 14945 11254 14945 11254 0 _01_
rlabel metal1 16682 12342 16682 12342 0 _02_
rlabel viali 13386 10097 13386 10097 0 _03_
rlabel metal2 13754 11492 13754 11492 0 _04_
rlabel metal1 14858 11696 14858 11696 0 _05_
rlabel metal1 15318 10778 15318 10778 0 _06_
rlabel metal1 17158 11866 17158 11866 0 _07_
rlabel metal1 17004 11594 17004 11594 0 _08_
rlabel metal1 16744 11798 16744 11798 0 _09_
rlabel metal1 14260 9146 14260 9146 0 clknet_0_i_stop
rlabel metal2 15410 9214 15410 9214 0 clknet_0_net3
rlabel metal2 12466 9996 12466 9996 0 clknet_1_0__leaf_i_stop
rlabel metal1 11178 11220 11178 11220 0 clknet_1_0__leaf_net3
rlabel metal2 18446 11424 18446 11424 0 clknet_1_1__leaf_i_stop
rlabel metal1 16238 10608 16238 10608 0 clknet_1_1__leaf_net3
rlabel metal1 13708 18802 13708 18802 0 i_start
rlabel metal2 13938 6256 13938 6256 0 i_stop
rlabel metal1 13616 11186 13616 11186 0 net1
rlabel metal2 17158 9044 17158 9044 0 net10
rlabel metal1 12282 6188 12282 6188 0 net100
rlabel metal1 12650 6834 12650 6834 0 net101
rlabel metal1 11776 6426 11776 6426 0 net102
rlabel metal2 12098 5848 12098 5848 0 net103
rlabel metal1 10810 6426 10810 6426 0 net104
rlabel metal1 11316 6630 11316 6630 0 net105
rlabel metal1 11224 10098 11224 10098 0 net106
rlabel metal1 9798 10234 9798 10234 0 net107
rlabel metal1 14766 10642 14766 10642 0 net108
rlabel metal1 16882 10506 16882 10506 0 net109
rlabel metal1 15870 7956 15870 7956 0 net11
rlabel metal1 13386 10642 13386 10642 0 net111
rlabel via1 11817 11662 11817 11662 0 net112
rlabel metal1 17618 11594 17618 11594 0 net113
rlabel metal1 15088 10642 15088 10642 0 net114
rlabel metal1 14030 11798 14030 11798 0 net115
rlabel metal1 13386 11288 13386 11288 0 net116
rlabel metal1 17250 10540 17250 10540 0 net117
rlabel metal1 16192 8398 16192 8398 0 net118
rlabel metal1 13800 10778 13800 10778 0 net119
rlabel metal1 16054 10574 16054 10574 0 net12
rlabel metal1 16238 9520 16238 9520 0 net120
rlabel metal1 16284 9146 16284 9146 0 net121
rlabel metal1 16330 10506 16330 10506 0 net122
rlabel metal2 16422 9792 16422 9792 0 net123
rlabel metal1 19826 7276 19826 7276 0 net124
rlabel metal1 18170 7310 18170 7310 0 net125
rlabel metal1 20654 9588 20654 9588 0 net126
rlabel metal1 15594 7888 15594 7888 0 net127
rlabel metal1 18400 6834 18400 6834 0 net128
rlabel metal1 17020 6630 17020 6630 0 net129
rlabel metal1 10074 8602 10074 8602 0 net13
rlabel metal1 19504 6698 19504 6698 0 net130
rlabel metal1 15962 6222 15962 6222 0 net131
rlabel viali 12922 7912 12922 7912 0 net132
rlabel metal2 14398 8160 14398 8160 0 net133
rlabel metal1 13570 6188 13570 6188 0 net134
rlabel metal1 13984 6970 13984 6970 0 net135
rlabel metal1 15042 6086 15042 6086 0 net136
rlabel metal2 13294 7616 13294 7616 0 net137
rlabel metal1 8602 8058 8602 8058 0 net138
rlabel metal1 9890 6834 9890 6834 0 net139
rlabel metal1 8418 9044 8418 9044 0 net14
rlabel metal2 9522 8500 9522 8500 0 net140
rlabel metal2 12558 6188 12558 6188 0 net141
rlabel metal1 13018 6800 13018 6800 0 net142
rlabel metal1 11362 6426 11362 6426 0 net143
rlabel metal1 12972 6630 12972 6630 0 net144
rlabel metal2 9062 10404 9062 10404 0 net145
rlabel metal1 11822 7956 11822 7956 0 net146
rlabel metal1 10672 8398 10672 8398 0 net147
rlabel metal1 12052 6834 12052 6834 0 net148
rlabel metal1 12098 10064 12098 10064 0 net149
rlabel metal2 8694 7548 8694 7548 0 net15
rlabel metal1 8878 9146 8878 9146 0 net150
rlabel metal1 10810 10166 10810 10166 0 net152
rlabel metal1 13110 10064 13110 10064 0 net153
rlabel metal1 10150 10506 10150 10506 0 net154
rlabel metal1 13938 10540 13938 10540 0 net155
rlabel metal1 12926 10098 12926 10098 0 net156
rlabel metal1 13524 10234 13524 10234 0 net157
rlabel metal1 14122 10778 14122 10778 0 net158
rlabel metal1 20286 10098 20286 10098 0 net159
rlabel metal1 10672 6222 10672 6222 0 net16
rlabel metal1 17710 7344 17710 7344 0 net160
rlabel metal1 18216 8398 18216 8398 0 net161
rlabel metal1 20562 6698 20562 6698 0 net162
rlabel metal1 20378 9486 20378 9486 0 net163
rlabel metal1 18216 8602 18216 8602 0 net164
rlabel metal1 20470 9350 20470 9350 0 net165
rlabel metal1 20654 8398 20654 8398 0 net166
rlabel metal1 14674 6834 14674 6834 0 net167
rlabel metal1 15042 7956 15042 7956 0 net168
rlabel metal2 14582 6562 14582 6562 0 net169
rlabel metal1 11684 5882 11684 5882 0 net17
rlabel metal1 16514 6868 16514 6868 0 net170
rlabel metal1 13892 8058 13892 8058 0 net171
rlabel metal2 14674 8432 14674 8432 0 net172
rlabel metal2 9798 6766 9798 6766 0 net173
rlabel metal1 11178 6256 11178 6256 0 net174
rlabel metal1 11408 7922 11408 7922 0 net175
rlabel metal2 13110 8823 13110 8823 0 net176
rlabel metal4 12604 7616 12604 7616 0 net177
rlabel metal2 9430 7004 9430 7004 0 net178
rlabel metal1 12834 5882 12834 5882 0 net179
rlabel metal1 10626 10166 10626 10166 0 net18
rlabel metal1 11776 8398 11776 8398 0 net180
rlabel metal2 8970 10642 8970 10642 0 net181
rlabel metal2 8786 7344 8786 7344 0 net182
rlabel metal1 11546 9486 11546 9486 0 net183
rlabel metal1 8924 9622 8924 9622 0 net184
rlabel metal1 8602 6800 8602 6800 0 net185
rlabel via2 12190 6715 12190 6715 0 net186
rlabel metal2 11362 10336 11362 10336 0 net187
rlabel metal1 13018 10200 13018 10200 0 net188
rlabel metal1 17342 8364 17342 8364 0 net19
rlabel via1 13731 9486 13731 9486 0 net2
rlabel metal1 15686 7990 15686 7990 0 net21
rlabel metal1 17107 10098 17107 10098 0 net22
rlabel metal1 18354 10540 18354 10540 0 net23
rlabel metal2 17710 8942 17710 8942 0 net25
rlabel metal1 19131 10166 19131 10166 0 net26
rlabel metal1 19550 7344 19550 7344 0 net27
rlabel metal2 17250 7004 17250 7004 0 net29
rlabel metal1 14260 9486 14260 9486 0 net3
rlabel metal1 18993 9078 18993 9078 0 net30
rlabel metal1 15916 7718 15916 7718 0 net31
rlabel metal1 18860 7514 18860 7514 0 net33
rlabel metal1 19688 7446 19688 7446 0 net34
rlabel metal2 12650 8602 12650 8602 0 net35
rlabel metal1 15548 6698 15548 6698 0 net37
rlabel metal1 19085 7922 19085 7922 0 net38
rlabel metal1 12098 8330 12098 8330 0 net39
rlabel metal1 12926 5780 12926 5780 0 net4
rlabel metal1 15318 6188 15318 6188 0 net41
rlabel metal1 17705 7922 17705 7922 0 net42
rlabel metal1 9338 8330 9338 8330 0 net43
rlabel metal1 12558 7888 12558 7888 0 net45
rlabel metal1 15916 6426 15916 6426 0 net46
rlabel metal1 8786 7990 8786 7990 0 net47
rlabel metal2 13110 6987 13110 6987 0 net49
rlabel metal1 12374 7956 12374 7956 0 net5
rlabel metal1 13892 5882 13892 5882 0 net50
rlabel metal1 10488 8398 10488 8398 0 net52
rlabel metal2 11270 6630 11270 6630 0 net53
rlabel metal2 11362 6528 11362 6528 0 net54
rlabel metal1 8970 9486 8970 9486 0 net56
rlabel metal1 11086 6188 11086 6188 0 net57
rlabel metal1 9138 7990 9138 7990 0 net58
rlabel metal1 10166 8398 10166 8398 0 net59
rlabel metal2 15134 6426 15134 6426 0 net6
rlabel metal1 12282 6086 12282 6086 0 net61
rlabel via1 9333 9010 9333 9010 0 net62
rlabel metal1 10258 10064 10258 10064 0 net63
rlabel via2 8234 9027 8234 9027 0 net65
rlabel metal1 13652 8398 13652 8398 0 net66
rlabel metal1 10626 8262 10626 8262 0 net68
rlabel metal1 12374 10506 12374 10506 0 net69
rlabel metal1 15548 6970 15548 6970 0 net7
rlabel via1 9425 9486 9425 9486 0 net70
rlabel metal2 12190 11492 12190 11492 0 net71
rlabel metal2 10718 10608 10718 10608 0 net72
rlabel metal1 14398 10540 14398 10540 0 net73
rlabel metal1 16514 8398 16514 8398 0 net74
rlabel metal1 15778 10642 15778 10642 0 net75
rlabel metal2 12742 10336 12742 10336 0 net76
rlabel metal1 14255 10166 14255 10166 0 net77
rlabel metal1 19458 10574 19458 10574 0 net78
rlabel metal2 17802 9180 17802 9180 0 net79
rlabel metal2 17434 7582 17434 7582 0 net8
rlabel metal2 16514 9962 16514 9962 0 net80
rlabel metal1 19734 9486 19734 9486 0 net81
rlabel metal1 18032 8534 18032 8534 0 net82
rlabel metal1 16100 8058 16100 8058 0 net83
rlabel metal1 18216 8534 18216 8534 0 net84
rlabel metal1 20010 7514 20010 7514 0 net85
rlabel metal1 15456 6834 15456 6834 0 net86
rlabel metal1 19412 6834 19412 6834 0 net87
rlabel metal2 13846 8296 13846 8296 0 net88
rlabel metal1 16284 6970 16284 6970 0 net89
rlabel metal1 17066 6868 17066 6868 0 net9
rlabel metal1 17986 6630 17986 6630 0 net90
rlabel metal1 15594 7786 15594 7786 0 net91
rlabel metal1 14122 5746 14122 5746 0 net92
rlabel metal1 12972 6426 12972 6426 0 net93
rlabel metal2 12834 7922 12834 7922 0 net94
rlabel metal2 10810 7854 10810 7854 0 net95
rlabel metal1 13662 6426 13662 6426 0 net96
rlabel metal1 12604 7718 12604 7718 0 net97
rlabel metal1 13156 6970 13156 6970 0 net98
rlabel metal2 8234 9690 8234 9690 0 net99
rlabel metal2 18722 18099 18722 18099 0 o_result_ctr[0]
rlabel metal2 20056 11322 20056 11322 0 o_result_ctr[1]
rlabel metal2 19366 18099 19366 18099 0 o_result_ctr[2]
rlabel metal2 12926 18099 12926 18099 0 o_result_ring[0]
rlabel metal2 12282 619 12282 619 0 o_result_ring[10]
rlabel metal3 1533 8228 1533 8228 0 o_result_ring[11]
rlabel metal2 11178 8857 11178 8857 0 o_result_ring[12]
rlabel metal1 14766 4114 14766 4114 0 o_result_ring[13]
rlabel via2 10166 9605 10166 9605 0 o_result_ring[14]
rlabel metal3 1533 10268 1533 10268 0 o_result_ring[15]
rlabel via3 15525 4012 15525 4012 0 o_result_ring[1]
rlabel metal2 18078 18099 18078 18099 0 o_result_ring[2]
rlabel metal2 31694 10217 31694 10217 0 o_result_ring[3]
rlabel metal2 28290 9367 28290 9367 0 o_result_ring[4]
rlabel via2 28290 8891 28290 8891 0 o_result_ring[5]
rlabel metal2 20010 4036 20010 4036 0 o_result_ring[6]
rlabel metal2 18722 1557 18722 1557 0 o_result_ring[7]
rlabel metal2 16790 415 16790 415 0 o_result_ring[8]
rlabel metal2 14858 415 14858 415 0 o_result_ring[9]
rlabel metal1 18722 10574 18722 10574 0 r_dly_store_ctr\[0\]
rlabel metal1 20010 11288 20010 11288 0 r_dly_store_ctr\[1\]
rlabel metal2 20102 12070 20102 12070 0 r_dly_store_ctr\[2\]
rlabel metal1 12926 11254 12926 11254 0 r_dly_store_ring\[0\]
rlabel metal1 12374 7208 12374 7208 0 r_dly_store_ring\[10\]
rlabel metal1 11086 8024 11086 8024 0 r_dly_store_ring\[11\]
rlabel metal1 10948 9010 10948 9010 0 r_dly_store_ring\[12\]
rlabel metal1 15042 8330 15042 8330 0 r_dly_store_ring\[13\]
rlabel metal1 10626 9418 10626 9418 0 r_dly_store_ring\[14\]
rlabel metal1 11730 10506 11730 10506 0 r_dly_store_ring\[15\]
rlabel metal1 15502 10200 15502 10200 0 r_dly_store_ring\[1\]
rlabel metal1 18400 9418 18400 9418 0 r_dly_store_ring\[2\]
rlabel metal1 19918 10200 19918 10200 0 r_dly_store_ring\[3\]
rlabel metal1 19826 9112 19826 9112 0 r_dly_store_ring\[4\]
rlabel metal1 20240 8602 20240 8602 0 r_dly_store_ring\[5\]
rlabel metal1 19826 7990 19826 7990 0 r_dly_store_ring\[6\]
rlabel metal1 18814 7344 18814 7344 0 r_dly_store_ring\[7\]
rlabel metal1 16974 7208 16974 7208 0 r_dly_store_ring\[8\]
rlabel metal1 14858 6902 14858 6902 0 r_dly_store_ring\[9\]
rlabel metal1 14950 11526 14950 11526 0 r_ring_ctr\[0\]
rlabel metal2 16514 11492 16514 11492 0 r_ring_ctr\[1\]
rlabel metal1 18400 12070 18400 12070 0 r_ring_ctr\[2\]
rlabel metal1 12581 10234 12581 10234 0 w_dly_strt\[1\]
rlabel metal1 12282 12240 12282 12240 0 w_dly_strt\[2\]
rlabel metal1 12374 11254 12374 11254 0 w_dly_strt\[3\]
rlabel metal1 14122 12308 14122 12308 0 w_ring_ctr_clk
rlabel metal2 13202 10404 13202 10404 0 w_strt_pulse
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
