* PEX produced on Fri Mar 29 11:25:02 PM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tdc_ring.ext - technology: sky130A

.subckt tdc_ring dbg_reset dbg_ring_ctr[0] dbg_ring_ctr[1] dbg_ring_ctr[2] dbg_ring_sig[10]
+ dbg_ring_sig[11] dbg_ring_sig[12] dbg_ring_sig[13] dbg_ring_sig[14] dbg_ring_sig[15]
+ dbg_ring_sig[2] dbg_ring_sig[5] dbg_ring_sig[7] dbg_ring_sig[9] i_start o_result_ctr[1]
+ o_result_ctr[2] o_result_ring[10] o_result_ring[12] o_result_ring[14] o_result_ring[15]
+ o_result_ring[2] o_result_ring[5] o_result_ring[7] o_result_ring[4] o_result_ring[9]
+ o_result_ring[1] dbg_ring_sig[4] dbg_ring_sig[1] dbg_ring_sig[6] o_result_ring[6]
+ o_result_ring[11] o_result_ring[3] o_result_ring[8] o_result_ring[0] o_result_ctr[0]
+ dbg_ring_sig[3] dbg_ring_sig[8] dbg_ring_sig[0] i_stop o_result_ring[13] VGND VPWR
X0 a_16861_11989# a_16643_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1 VGND a_15071_11146# _01_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5 a_16459_10383# a_16109_10383# a_16364_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X9 VPWR a_13323_10058# w_ring_buf[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X10 net6 a_15667_7671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X13 VGND r_dly_store_ring[8] a_16127_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X14 w_ring_buf[1] a_16495_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X16 r_dly_store_ring[6] a_10443_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 r_dly_store_ring[3] a_19827_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 a_16677_10625# a_16459_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X24 a_13441_12021# a_13275_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VPWR a_18151_9839# o_result_ring[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 a_19793_8207# w_ring_buf[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_14223_12015# a_13441_12021# a_14139_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X33 a_18027_8181# w_ring_buf[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X34 VPWR a_14563_9295# dbg_ring_sig[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X37 a_17208_12393# a_16293_12021# a_16861_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X38 o_result_ring[8] a_16127_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X44 VPWR w_ring_norsz[8] a_14103_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X46 VPWR a_19991_9295# o_result_ring[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X47 VGND net1 w_ring_int_norsz[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X48 VGND a_10699_7119# o_result_ring[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X49 dbg_ring_ctr[2] a_18763_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X57 a_19973_11837# a_19439_11471# a_19878_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X59 a_19142_10749# a_18703_10383# a_19057_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X61 a_12500_11445# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X65 a_12173_8751# w_ring_int_norsz[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X66 r_dly_store_ring[14] a_10443_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X67 w_ring_norsz[1] w_ring_int_norsz[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VGND a_20303_8573# a_20471_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X72 VGND a_14583_7387# a_14541_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X78 VPWR a_10563_8372# w_ring_buf[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X79 w_ring_norsz[1] net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X84 a_11901_8751# w_ring_norsz[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X89 w_ring_buf[3] a_18703_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X91 VGND a_18763_11445# dbg_ring_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X94 VGND a_20175_10383# o_result_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X96 r_dly_store_ctr[1] a_20471_11739# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X101 a_9765_8751# w_ring_buf[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X104 a_12500_11445# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X107 o_result_ring[1] a_18151_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X112 r_dly_store_ring[1] a_17711_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X118 VPWR i_start a_12355_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X119 a_11759_8372# w_ring_norsz[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X121 VGND net7 a_11343_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X124 VGND a_10975_9839# o_result_ring[6] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X132 VGND a_20911_11471# o_result_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X138 a_12797_10933# a_12631_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
R0 VGND net15 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X140 a_14415_7485# a_13551_7119# a_14158_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X141 a_17635_7663# a_16937_7669# a_17378_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X142 VGND a_10443_7637# a_10401_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X143 a_17562_12381# _05_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X144 a_11141_10933# a_10975_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X145 VGND a_12355_591# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X147 net2 a_9814_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X149 a_12725_9545# w_ring_int_norsz[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X150 VPWR w_ring_norsz[4] a_14001_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X160 VPWR w_ring_int_norsz[5] a_13717_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X164 VPWR a_10018_9813# a_9945_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X165 VGND a_9747_7093# dbg_ring_sig[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X166 r_dly_store_ctr[2] a_19735_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X169 VGND a_10275_9839# a_10443_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X172 VPWR net5 _04_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X173 r_dly_store_ring[9] a_20379_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X177 a_20387_8573# a_19605_8207# a_20303_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X179 dbg_ring_sig[8] a_14563_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X181 a_16459_10383# a_15943_10383# a_16364_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
R1 net14 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X185 VGND w_ring_norsz[11] w_ring_int_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X186 o_result_ctr[0] a_20175_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X187 VPWR w_ring_norsz[9] a_17405_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X189 a_17627_9839# a_16845_9845# a_17543_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X190 w_ring_norsz[15] net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X194 VGND net7 a_13275_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X195 a_16293_9545# w_ring_norsz[1] a_16209_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 VGND _07_ a_18057_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X200 o_result_ring[4] a_14839_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X202 VGND r_ring_ctr[0] a_18141_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X203 o_result_ring[8] a_16127_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X208 VPWR a_10018_8725# a_9945_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X210 _05_ net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X211 a_9556_8181# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X216 w_ring_norsz[2] net4 a_15937_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X219 VPWR w_ring_norsz[12] a_14747_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X220 a_20429_11471# a_19439_11471# a_20303_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X225 VGND a_14747_12015# o_result_ring[0] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X226 VPWR a_18887_7119# dbg_ring_sig[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X228 VPWR a_14583_7387# a_14499_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X229 a_18869_10383# a_18703_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X233 VGND w_ring_norsz[9] a_18887_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X234 VPWR a_17383_12319# a_17370_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X244 VGND w_ring_buf[1] a_16771_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X247 a_19912_10217# a_19513_9845# a_19786_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R2 g_ring3[12].stg01_11.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X261 VPWR a_18027_8181# dbg_ring_sig[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X262 a_14369_8457# net1 w_ring_int_norsz[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X263 o_result_ring[6] a_10975_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X266 VGND a_20083_10935# _60_.X VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X268 r_dly_store_ring[2] a_19367_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X272 VPWR net6 a_18703_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X277 a_14116_7119# a_13717_7119# a_13990_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X278 VGND a_19827_7637# a_19785_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X279 a_19878_8573# a_19605_8207# a_19793_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X280 a_18763_11445# r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X285 dbg_ring_sig[1] a_16771_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X288 o_result_ring[1] a_18151_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X293 VGND net7 a_9411_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X294 a_13795_11445# w_ring_buf[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X295 VGND a_10851_10357# dbg_ring_sig[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X296 VGND w_ring_norsz[10] w_ring_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X299 a_19651_10749# a_18869_10383# a_19567_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X301 _00_ r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X302 VGND a_12500_10357# net4 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X309 o_result_ring[2] a_19991_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X310 r_dly_store_ring[3] a_19827_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X314 a_15887_7485# a_15189_7119# a_15630_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X315 a_18961_7669# a_18795_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X318 VGND net7 a_10975_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X324 a_20004_11471# a_19605_11471# a_19878_11837# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X327 r_dly_store_ctr[1] a_20471_11739# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X330 VGND a_14158_7231# a_14116_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X331 w_ring_buf[11] a_16403_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X335 VGND a_9747_7093# dbg_ring_sig[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X336 VPWR a_17659_11623# _08_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X339 a_17210_7663# a_16771_7669# a_17125_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X340 VGND a_18887_7119# dbg_ring_sig[3] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
R3 VGND net13 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X345 _04_ net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X346 w_ring_int_norsz[3] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X347 net3 a_12224_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X350 VGND w_ring_int_norsz[13] w_ring_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X351 a_11923_10927# a_11141_10933# a_11839_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X355 VGND a_13323_10058# w_ring_buf[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X356 a_13714_12015# a_13275_12021# a_13629_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X363 a_11540_11305# a_11141_10933# a_11414_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X367 VGND a_12875_10357# dbg_ring_sig[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X368 w_ring_norsz[4] net3 a_15109_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X374 a_17336_8041# a_16937_7669# a_17210_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X379 a_18057_12335# a_18015_12247# _02_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.195 ps=1.9 w=0.65 l=0.15
X383 VPWR a_12875_10357# dbg_ring_sig[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X386 VGND w_ring_buf[0] a_15943_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X389 a_17033_9839# w_ring_buf[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X397 a_19973_8573# a_19439_8207# a_19878_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X398 a_15887_7485# a_15023_7119# a_15630_7231# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X399 VGND r_dly_store_ctr[2] a_20175_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X400 a_12985_10927# w_ring_buf[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X407 VGND a_14563_9295# dbg_ring_sig[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X409 VPWR i_stop a_9814_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X411 a_19402_7637# a_19234_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X427 o_result_ctr[2] a_20175_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X429 a_9850_9839# a_9577_9845# a_9765_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X436 a_15076_11471# _01_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X437 VGND w_ring_norsz[8] a_14103_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X445 a_19310_11989# a_19142_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X447 w_ring_norsz[4] w_ring_int_norsz[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X448 a_9765_9839# w_ring_buf[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X450 dbg_ring_sig[2] a_17783_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X453 a_19142_12015# a_18869_12021# a_19057_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X457 VPWR r_dly_store_ring[9] a_21279_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X459 VPWR r_ring_ctr[1] a_19531_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X460 a_19567_10749# a_18703_10383# a_19310_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X463 a_19237_10749# a_18703_10383# a_19142_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X464 VPWR a_11863_10357# o_result_ring[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X465 VPWR w_ring_int_norsz[12] a_14729_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X468 VPWR w_ring_int_norsz[11] a_16293_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X469 a_9850_8751# a_9577_8757# a_9765_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X472 VPWR a_13795_11445# dbg_ring_sig[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X474 VPWR a_16677_10625# a_16567_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
R4 VGND net11 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X482 VGND a_10018_8725# a_9976_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X486 a_15462_7485# a_15023_7119# a_15377_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X489 VPWR a_14103_10927# o_result_ring[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X492 a_11858_7637# a_11690_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X496 a_19310_10495# a_19142_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X498 r_dly_store_ring[14] a_10443_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X499 o_result_ctr[1] a_20911_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X501 VPWR r_dly_store_ring[10] a_21279_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X503 VPWR r_dly_store_ring[1] a_18151_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X504 a_11417_7669# a_11251_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X505 dbg_ring_sig[10] a_18027_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X508 a_16555_10383# a_16109_10383# a_16459_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X509 w_ring_int_norsz[8] net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X513 a_11509_10927# a_10975_10933# a_11414_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X514 VPWR a_19439_9295# dbg_ring_sig[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X516 w_ring_norsz[0] net4 a_12717_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X517 VGND a_21279_9839# o_result_ring[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X518 a_19605_11471# a_19439_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X521 VPWR a_15911_11445# a_15898_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X522 a_10275_7663# a_9411_7669# a_10018_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X524 VGND net3 w_ring_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X527 VGND r_dly_store_ring[0] a_14747_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X529 VPWR a_19991_9295# o_result_ring[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X533 a_15588_7119# a_15189_7119# a_15462_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X535 w_ring_int_norsz[14] net13 a_11901_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X543 VPWR a_14839_6575# o_result_ring[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X548 r_ring_ctr[1] a_15911_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X549 a_19402_7637# a_19234_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X558 w_ring_int_norsz[15] w_ring_norsz[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X564 dbg_ring_sig[2] a_17783_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X567 a_13809_12015# a_13275_12021# a_13714_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X568 VGND a_12723_7663# o_result_ring[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X570 a_10310_591# a_10133_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X573 VGND a_15630_7231# a_15588_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X575 VGND dbg_reset a_12355_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X576 VPWR _07_ a_18015_12247# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X581 dbg_ring_sig[9] a_19439_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X582 VGND net3 w_ring_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R5 VPWR stg01_16.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X587 VPWR w_ring_int_norsz[6] a_12613_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X592 a_15076_11471# _01_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X593 a_16677_10625# a_16459_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X594 VPWR net6 a_19347_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X597 w_ring_buf[3] a_18703_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X601 VPWR a_10443_7637# a_10359_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X603 a_17180_11721# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X604 VGND w_ring_buf[9] a_19439_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X607 a_20046_8319# a_19878_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X608 VPWR net7 a_9411_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X609 a_20046_8319# a_19878_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X610 _03_ net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X612 o_result_ring[2] a_19991_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X615 VGND w_ring_buf[0] a_14655_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X616 _06_ a_17180_11721# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X617 a_17659_11623# _06_ a_17833_11499# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X622 dbg_ring_ctr[1] a_19531_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X623 a_14944_10217# a_14545_9845# a_14818_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X624 a_11858_7637# a_11690_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X628 a_19057_12015# r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X629 VPWR a_18763_11445# dbg_ring_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X636 a_10851_10357# w_ring_buf[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X637 a_18141_11471# r_ring_ctr[1] _07_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X641 a_16109_10383# a_15943_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X643 VGND net6 a_18703_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X646 dbg_ring_sig[8] a_14563_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X649 a_15377_7119# w_ring_buf[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X652 dbg_ring_sig[4] a_13735_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X654 o_result_ctr[1] a_20911_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X661 a_13070_10927# a_12631_10933# a_12985_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
R6 VGND net8 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X662 a_16567_10749# a_15943_10383# a_16459_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X663 VPWR a_19735_11989# a_19651_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X666 VPWR r_dly_store_ring[8] a_16127_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X672 VPWR a_12723_7663# o_result_ring[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X673 VPWR w_ring_norsz[10] a_17415_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X676 VPWR r_dly_store_ctr[1] a_20911_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X678 a_15898_11837# a_14821_11471# a_15736_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X681 VPWR a_10379_9460# w_ring_buf[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X682 a_13905_7119# w_ring_buf[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X684 a_19605_8207# a_19439_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X686 r_dly_store_ring[2] a_19367_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X688 VPWR a_10699_7119# o_result_ring[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X692 dbg_reset a_11895_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X694 a_18774_8751# a_18335_8757# a_18689_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X697 a_15937_9545# w_ring_norsz[9] a_15853_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X698 VGND w_ring_buf[5] a_11619_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X699 a_16209_8751# net4 w_ring_norsz[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X700 a_12875_10357# w_ring_buf[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X703 a_13257_8457# w_ring_norsz[4] a_13173_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X706 w_ring_int_norsz[14] w_ring_norsz[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X708 a_19268_10383# a_18869_10383# a_19142_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X712 VGND a_11863_10357# o_result_ring[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X714 r_dly_store_ctr[0] a_19735_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X715 a_9839_9269# w_ring_buf[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X719 dbg_ring_sig[12] a_15115_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X723 VPWR a_18027_8181# dbg_ring_sig[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X726 w_ring_int_norsz[11] net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X730 VGND a_14747_12015# o_result_ring[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X732 net4 a_12500_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X733 _60_.X a_20083_10935# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X736 a_18900_9129# a_18501_8757# a_18774_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X738 VGND i_stop a_9814_591# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X750 a_19659_7663# a_18961_7669# a_19402_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X754 a_9577_7669# a_9411_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X757 VPWR net7 a_14379_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X761 VPWR a_20303_8573# a_20471_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X762 a_19199_8751# a_18501_8757# a_18942_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X769 a_14541_7119# a_13551_7119# a_14415_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X776 VPWR a_20379_9813# a_20295_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X779 VGND a_18243_7663# o_result_ring[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X782 r_dly_store_ring[6] a_10443_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X785 dbg_ring_ctr[1] a_19531_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X787 a_19199_8751# a_18335_8757# a_18942_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X788 VPWR a_18303_11187# dbg_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X791 a_19693_12393# a_18703_12021# a_19567_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X799 VGND a_10699_7119# o_result_ring[13] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X802 a_19605_8207# a_19439_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X805 VGND w_ring_norsz[4] a_13643_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X809 VGND a_19531_10927# dbg_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
R7 g_ring3[9].stg01_15.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X815 o_result_ring[3] a_20267_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X816 a_12529_8751# net3 w_ring_norsz[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X817 VPWR net2 a_10133_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X818 VPWR a_10851_10357# dbg_ring_sig[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X820 VPWR a_19439_9295# dbg_ring_sig[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X821 VPWR w_ring_norsz[14] a_9135_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X822 a_14158_7231# a_13990_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X824 VGND net4 w_ring_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X825 VGND net5 _05_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X828 o_result_ring[15] a_14103_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X830 a_15389_11713# a_15171_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X834 VGND a_15243_9839# a_15411_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X836 VGND net7 a_12631_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X837 dbg_ring_sig[12] a_15115_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X839 VGND w_ring_buf[3] a_18887_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X845 a_20211_9839# a_19513_9845# a_19954_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X846 VPWR a_14839_6575# o_result_ring[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X851 a_12115_7663# a_11251_7669# a_11858_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X853 VGND w_ring_int_norsz[9] w_ring_norsz[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X854 dbg_reset a_11895_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X857 VGND r_dly_store_ring[6] a_10975_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
R8 g_ring3[11].stg01_10.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X862 a_10401_10217# a_9411_9845# a_10275_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X865 VPWR a_19367_8725# a_19283_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X869 a_15911_11445# a_15736_11471# a_16090_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X871 a_18961_7669# a_18795_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X875 VPWR w_dly_stop[2] a_11895_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X878 a_13449_7663# net12 w_ring_int_norsz[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X879 VGND a_20175_12015# o_result_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X884 a_18869_12021# a_18703_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X886 a_11690_7663# a_11251_7669# a_11605_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X888 VGND net7 a_9411_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X891 VPWR a_12875_10357# dbg_ring_sig[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X898 VGND a_19735_10651# a_19693_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X899 VGND a_14563_9295# dbg_ring_sig[8] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X901 VPWR a_18243_7663# o_result_ring[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X908 VGND a_9556_8181# net7 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X909 VGND w_ring_norsz[10] a_17415_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X910 VGND a_19991_9295# o_result_ring[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X912 VPWR a_13735_6575# dbg_ring_sig[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X917 o_result_ctr[0] a_20175_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X923 dbg_ring_ctr[0] a_18303_11187# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X927 a_11816_8041# a_11417_7669# a_11690_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X930 VGND a_10379_9460# w_ring_buf[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X934 o_result_ring[3] a_20267_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X935 VPWR a_12283_7637# a_12199_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X939 VGND a_17783_8751# dbg_ring_sig[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X942 r_dly_store_ctr[2] a_19735_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X945 a_18027_8181# w_ring_buf[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X949 VPWR a_18303_11187# dbg_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X957 VGND r_dly_store_ring[12] a_16495_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X963 VGND a_18303_11187# dbg_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X964 VGND a_19531_10927# dbg_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X965 VPWR net6 a_16771_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X966 VGND a_11759_8372# w_ring_buf[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X969 a_17543_9839# a_16845_9845# a_17286_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X971 VGND a_15115_7663# dbg_ring_sig[12] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X975 a_16293_12021# a_16127_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X978 a_12115_7663# a_11417_7669# a_11858_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X979 o_result_ring[0] a_14747_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X982 VPWR a_17199_10357# a_17186_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X983 o_result_ring[15] a_14103_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X985 r_dly_store_ring[12] a_16055_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X988 a_15911_11445# _04_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X993 a_13840_12393# a_13441_12021# a_13714_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X994 a_16861_11989# a_16643_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1001 a_17118_9839# a_16845_9845# a_17033_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1002 dbg_ring_sig[14] a_9963_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1011 dbg_ring_sig[6] a_9839_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1015 a_13649_9545# w_ring_norsz[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1018 r_dly_store_ring[7] a_12007_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1019 dbg_ring_sig[1] a_16771_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1022 dbg_ring_sig[7] a_10851_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1023 VGND a_10443_8725# a_10401_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1024 a_10593_591# a_10416_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1026 o_result_ring[11] a_18243_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1031 dbg_ring_sig[12] a_15115_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1033 VPWR net6 a_16679_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1034 VPWR r_dly_store_ring[4] a_14839_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1036 a_20303_11837# a_19439_11471# a_20046_11583# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1038 VPWR a_17635_7663# a_17803_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1044 VGND net15 w_ring_int_norsz[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1047 a_9747_7093# w_ring_buf[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1048 VGND w_ring_norsz[14] a_9135_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1050 a_17719_7663# a_16937_7669# a_17635_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1053 a_17383_12319# _05_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1054 VPWR a_17783_8751# dbg_ring_sig[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1055 a_17833_11499# _07_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X1058 VPWR a_20046_8319# a_19973_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1060 VGND w_ring_int_norsz[5] w_ring_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1061 VGND a_12868_11445# _59_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1062 a_11863_10357# r_dly_store_ring[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1065 VGND a_20267_7663# o_result_ring[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1066 r_dly_store_ring[0] a_14307_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1067 a_11417_7669# a_11251_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1070 r_dly_store_ring[0] a_14307_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1071 a_15305_9545# w_ring_norsz[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1072 dbg_ring_sig[9] a_19439_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1077 VGND a_14415_7485# a_14583_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1080 a_10018_7637# a_9850_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1081 VGND _04_ a_15433_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1082 a_20046_11583# a_19878_11837# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1085 VPWR a_17286_9813# a_17213_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1091 VPWR a_20046_11583# a_19973_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1092 VPWR r_dly_store_ctr[0] a_20175_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
R9 VGND net10 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1098 VPWR a_15115_7663# dbg_ring_sig[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1100 VGND a_13663_10901# a_13621_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1104 w_ring_int_norsz[6] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1105 a_13085_9839# w_ring_norsz[15] a_13001_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1111 dbg_ring_ctr[0] a_18303_11187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1112 VGND net3 w_ring_norsz[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1116 o_result_ring[4] a_14839_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1117 a_9556_8181# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1118 a_9850_8751# a_9411_8757# a_9765_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1119 VGND r_ring_ctr[0] _00_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1120 VPWR w_ring_norsz[2] a_17783_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1124 a_14986_9813# a_14818_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1125 r_dly_store_ring[12] a_16055_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1126 a_12257_8751# w_ring_norsz[5] a_12173_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1127 VGND w_ring_norsz[8] w_ring_norsz[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1129 r_dly_store_ring[10] a_20471_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1130 dbg_ring_sig[14] a_9963_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1132 a_17213_9839# a_16679_9845# a_17118_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1133 a_12357_9545# w_ring_int_norsz[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1137 o_result_ring[5] a_12723_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1147 VPWR w_ring_norsz[1] a_16495_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1150 VGND a_16127_9839# o_result_ring[8] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1158 a_9976_9129# a_9577_8757# a_9850_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1159 r_ring_ctr[2] a_17383_12319# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1160 VGND w_ring_buf[0] a_16127_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1162 a_9850_7663# a_9411_7669# a_9765_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1165 VPWR a_18763_11445# dbg_ring_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1168 a_18303_11187# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X1169 o_result_ring[11] a_18243_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1173 a_17186_10749# a_16109_10383# a_17024_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1174 dbg_ring_sig[12] a_15115_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1176 a_12985_10927# w_ring_buf[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1178 o_result_ring[2] a_19991_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1183 VGND net2 a_10133_591# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1184 VPWR w_dly_stop[1] a_11619_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1185 VGND w_ring_norsz[11] a_16403_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1186 w_ring_int_norsz[4] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1188 w_dly_stop[2] a_11619_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1195 VGND net7 a_9411_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1198 a_14499_7485# a_13717_7119# a_14415_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1203 VGND a_12500_11445# _99_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1204 r_dly_store_ring[7] a_12007_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1205 VGND net6 a_16679_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1210 a_12809_9545# w_ring_norsz[14] a_12725_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1211 net1 a_12355_591# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X1212 a_9976_8041# a_9577_7669# a_9850_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1213 VPWR a_20267_7663# o_result_ring[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1214 VGND r_dly_store_ring[10] a_21279_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1216 VPWR a_11839_10927# a_12007_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1221 dbg_ring_sig[2] a_17783_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1226 VPWR r_dly_store_ring[13] a_10699_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1229 VGND a_14839_6575# o_result_ring[4] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1234 VPWR net2 a_15667_7671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1237 a_15071_11146# _08_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1239 a_20337_10217# a_19347_9845# a_20211_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1246 a_10018_7637# a_9850_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1247 a_15243_9839# a_14379_9845# a_14986_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1248 VGND a_19367_8725# a_19325_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1249 a_19567_12015# a_18869_12021# a_19310_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1250 r_dly_store_ring[1] a_17711_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1252 o_result_ctr[1] a_20911_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1253 VGND r_ring_ctr[1] a_17180_11721# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1255 VPWR a_9963_8207# dbg_ring_sig[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1258 VGND net4 _03_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1263 _59_.X a_12868_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1269 VPWR a_14139_12015# a_14307_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1270 VPWR w_ring_int_norsz[10] a_16293_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1272 VGND a_14139_12015# a_14307_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1273 o_result_ring[5] a_12723_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1277 a_17024_10383# a_16109_10383# a_16677_10625# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1279 VPWR w_ring_buf[2] a_17783_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1281 a_19954_9813# a_19786_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1282 a_18501_8757# a_18335_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1286 net3 a_12224_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1290 a_16364_10383# _00_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1292 VGND net1 w_ring_int_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1293 o_result_ring[13] a_10699_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1295 VGND a_9839_9269# dbg_ring_sig[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1297 a_14139_12015# a_13275_12021# a_13882_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1300 w_ring_norsz[4] net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1303 VGND a_13882_11989# a_13840_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1304 a_18869_10383# a_18703_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1308 net6 a_15667_7671# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1309 VPWR a_10275_7663# a_10443_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1313 net7 a_9556_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1316 VGND a_18243_7663# o_result_ring[11] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1322 VPWR a_20175_10383# o_result_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1326 VGND a_15115_7663# dbg_ring_sig[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1328 a_14361_9545# w_ring_norsz[0] a_14277_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1329 VPWR a_10310_591# a_10416_591# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X1331 a_10275_9839# a_9577_9845# a_10018_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1334 o_result_ring[3] a_20267_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1335 VGND a_16127_9839# o_result_ring[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1339 VPWR r_dly_store_ring[2] a_19991_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1340 VPWR a_15411_9813# a_15327_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1348 VPWR a_19659_7663# a_19827_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1350 dbg_ring_sig[2] a_17783_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1352 VGND a_20379_9813# a_20337_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1355 VPWR r_dly_store_ctr[2] a_20175_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1356 o_result_ring[14] a_10975_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1361 VGND a_17635_7663# a_17803_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1362 a_13196_11305# a_12797_10933# a_13070_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1364 dbg_ring_sig[4] a_13735_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1369 w_ring_norsz[2] w_ring_int_norsz[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1372 a_9577_7669# a_9411_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1374 a_17669_10217# a_16679_9845# a_17543_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1375 w_ring_norsz[3] net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1378 VPWR w_ring_norsz[4] a_13643_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1379 a_16090_11471# _04_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1380 o_result_ring[1] a_18151_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1381 VGND a_9963_8207# dbg_ring_sig[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1383 dbg_ring_sig[13] a_9747_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1387 a_18689_8751# w_ring_buf[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1388 a_11391_10548# w_ring_norsz[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1389 a_19701_9839# w_ring_buf[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1390 a_13717_7119# a_13551_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1391 VPWR w_ring_buf[4] a_13735_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1392 o_result_ring[11] a_18243_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1394 VGND a_11839_10927# a_12007_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1395 VGND a_10975_9839# o_result_ring[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1397 VGND w_ring_norsz[2] a_17783_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1399 a_10563_8372# w_ring_norsz[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1405 VPWR a_20083_10935# _60_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1406 r_ring_ctr[0] a_17199_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1407 a_10275_9839# a_9411_9845# a_10018_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1409 o_result_ring[13] a_10699_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1411 VGND a_19310_10495# a_19268_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1415 VGND a_19439_9295# dbg_ring_sig[9] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1417 a_17286_9813# a_17118_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1420 VGND w_ring_int_norsz[12] w_ring_norsz[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1421 a_15381_8457# net11 w_ring_int_norsz[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1423 a_15845_11471# a_14655_11471# a_15736_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1424 VGND a_11582_10901# a_11540_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1425 VPWR a_12224_9813# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1426 VGND w_ring_norsz[1] a_16495_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1429 VGND a_19991_9295# o_result_ring[2] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1432 o_result_ring[6] a_10975_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1435 o_result_ctr[1] a_20911_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1437 a_10275_8751# a_9577_8757# a_10018_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1438 a_17286_9813# a_17118_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1444 a_16673_8751# w_ring_norsz[10] a_16589_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1449 w_ring_norsz[8] w_ring_int_norsz[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1451 VGND a_12355_12015# net5 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1452 VGND a_18763_11445# dbg_ring_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1453 a_19954_9813# a_19786_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1454 VPWR a_18243_7663# o_result_ring[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1457 VPWR a_15115_7663# dbg_ring_sig[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1459 a_11605_7663# w_ring_buf[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1460 w_ring_int_norsz[10] net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1461 dbg_ring_sig[4] a_13735_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1462 a_10275_8751# a_9411_8757# a_10018_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1464 VGND w_dly_stop[1] a_11619_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1468 o_result_ring[3] a_20267_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1472 w_dly_stop[2] a_11619_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1475 a_16364_10383# _00_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
R10 g_ring2[8].stg01_8.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1476 o_result_ctr[0] a_20175_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1480 dbg_reset a_11895_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1485 o_result_ring[14] a_10975_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1488 a_10275_7663# a_9577_7669# a_10018_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1490 dbg_ring_sig[5] a_11619_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1492 VGND net6 a_18703_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1493 VGND a_17711_9813# a_17669_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1496 a_15841_8751# net1 w_ring_int_norsz[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1499 dbg_ring_sig[9] a_19439_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1504 VPWR a_14103_10927# o_result_ring[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1508 VGND a_17378_7637# a_17336_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1509 a_13717_8457# w_ring_norsz[12] a_13633_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1511 VPWR r_dly_store_ring[0] a_14747_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1514 VGND w_ring_norsz[3] a_18703_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1517 VPWR a_10443_9813# a_10359_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1522 VPWR a_20211_9839# a_20379_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1527 o_result_ring[7] a_11863_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1528 a_19149_7663# w_ring_buf[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1531 a_13717_7119# a_13551_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1532 r_dly_store_ring[8] a_15411_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1533 a_12797_10933# a_12631_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1535 w_ring_norsz[11] w_ring_norsz[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1537 o_result_ring[11] a_18243_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1541 w_ring_buf[12] a_14747_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1543 a_11809_9545# w_ring_norsz[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1545 o_result_ring[2] a_19991_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1550 VPWR a_11759_8372# w_ring_buf[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1551 dbg_ring_sig[14] a_9963_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1552 a_14821_11471# a_14655_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1553 VGND w_ring_norsz[12] w_ring_int_norsz[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1554 a_16209_9545# net4 w_ring_norsz[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1561 VGND a_20471_11739# a_20429_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1564 a_15736_11471# a_14821_11471# a_15389_11713# VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1568 VPWR dbg_reset a_12355_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1569 a_18942_8725# a_18774_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1570 VPWR a_10443_8725# a_10359_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1573 o_result_ring[0] a_14747_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1574 VPWR net7 a_9411_9845# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1579 a_17543_9839# a_16679_9845# a_17286_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1580 VGND w_ring_norsz[6] w_ring_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1583 a_18942_8725# a_18774_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1585 a_9577_9845# a_9411_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1586 a_20211_9839# a_19347_9845# a_19954_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1587 VGND a_14839_6575# o_result_ring[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1588 VPWR a_20175_12015# o_result_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1590 VPWR w_ring_norsz[3] a_14369_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1595 VPWR a_16771_9295# dbg_ring_sig[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1596 w_ring_int_norsz[2] net1 a_15305_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1605 VPWR a_16055_7387# a_15971_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1607 a_12224_9813# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1609 dbg_ring_sig[5] a_11619_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1613 VGND net6 a_16771_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1614 a_15171_11471# a_14821_11471# a_15076_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1616 a_19142_10749# a_18869_10383# a_19057_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1617 a_13921_9545# w_ring_int_norsz[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1618 VPWR a_19199_8751# a_19367_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1619 dbg_ring_sig[7] a_10851_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1620 VGND a_20267_7663# o_result_ring[3] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1622 VGND a_10275_7663# a_10443_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R11 net9 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1624 a_19057_12015# r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1626 VGND w_ring_norsz[7] w_ring_int_norsz[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1627 w_ring_norsz[1] net3 a_14005_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1631 VGND a_13238_10901# a_13196_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1635 a_10359_7663# a_9577_7669# a_10275_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1638 VGND a_10975_8751# o_result_ring[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1639 dbg_ring_sig[7] a_10851_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1641 w_ring_norsz[7] net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1646 a_11839_10927# a_10975_10933# a_11582_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1649 VGND a_13735_6575# dbg_ring_sig[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1650 w_ring_norsz[3] w_ring_int_norsz[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1653 w_ring_norsz[6] w_ring_norsz[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1656 VPWR a_17711_9813# a_17627_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1658 VGND a_19659_7663# a_19827_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 dbg_reset a_11895_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1663 dbg_ring_sig[14] a_9963_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1666 VPWR a_9747_7093# dbg_ring_sig[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1667 VPWR net6 a_18795_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1668 a_11391_10548# w_ring_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1672 a_11414_10927# a_11141_10933# a_11329_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1674 VGND net14 w_ring_int_norsz[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1675 VGND net1 w_ring_int_norsz[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1680 VGND r_dly_store_ring[15] a_14103_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1687 a_16643_12393# a_16293_12021# a_16548_12381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1688 o_result_ring[9] a_21279_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1694 VPWR a_12115_7663# a_12283_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1696 VPWR a_12355_591# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1698 VPWR a_15736_11471# a_15911_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1699 net2 a_9814_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1702 VPWR net6 a_15023_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1703 w_ring_norsz[13] w_ring_norsz[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1707 _99_.X a_12500_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1709 a_17125_7663# w_ring_buf[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1710 VGND a_10310_591# a_10416_591# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1711 o_result_ring[12] a_16495_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1713 VPWR a_10975_9839# o_result_ring[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1718 a_15109_8457# w_ring_norsz[11] a_15025_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1719 a_13714_12015# a_13441_12021# a_13629_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1721 VPWR w_ring_buf[11] a_16863_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1725 o_result_ctr[2] a_20175_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1726 VGND w_ring_norsz[4] w_ring_int_norsz[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1727 a_17761_8041# a_16771_7669# a_17635_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1729 a_9577_8757# a_9411_8757# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1731 a_17208_12393# a_16127_12021# a_16861_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1737 a_19878_8573# a_19439_8207# a_19793_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1740 VPWR a_13735_6575# dbg_ring_sig[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1744 VPWR a_20267_7663# o_result_ring[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1745 a_9765_7663# w_ring_buf[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1746 a_20387_11837# a_19605_11471# a_20303_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1747 VGND w_ring_norsz[15] w_ring_norsz[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1752 w_ring_norsz[15] net3 a_12441_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1753 VGND w_ring_buf[8] a_14563_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1756 VPWR w_ring_norsz[11] a_16403_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1762 a_19310_10495# a_19142_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1764 VPWR r_ring_ctr[0] _07_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1765 VPWR a_10975_8751# o_result_ring[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1766 a_16643_12393# a_16127_12021# a_16548_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1769 VPWR a_17208_12393# a_17383_12319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1770 _05_ net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1771 VPWR a_11619_7119# dbg_ring_sig[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1775 VGND a_19735_11989# a_19693_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1776 VGND a_19439_9295# dbg_ring_sig[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1784 a_18869_8751# a_18335_8757# a_18774_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1787 VPWR w_ring_buf[14] a_9963_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1789 a_10018_9813# a_9850_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1791 a_20004_8207# a_19605_8207# a_19878_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1792 a_19743_7663# a_18961_7669# a_19659_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1796 o_result_ctr[2] a_20175_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1798 a_15171_11471# a_14655_11471# a_15076_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1800 a_14385_8751# w_ring_norsz[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
R12 VGND net12 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1802 w_ring_int_norsz[0] w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1806 VGND a_15911_11445# a_15845_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1808 _03_ net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1810 VPWR w_ring_buf[1] a_16771_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1811 dbg_ring_sig[10] a_18027_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1819 VPWR a_11858_7637# a_11785_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1821 VPWR a_13495_10927# a_13663_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1823 VPWR a_9963_8207# dbg_ring_sig[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1827 VGND net6 a_15023_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1828 a_14733_9839# w_ring_buf[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1834 a_13990_7485# a_13717_7119# a_13905_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1836 VPWR a_9747_7093# dbg_ring_sig[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1841 a_14729_8457# w_ring_norsz[3] a_14645_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1843 a_18763_11445# r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1844 a_13495_10927# a_12631_10933# a_13238_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1847 a_19234_7663# a_18795_7669# a_19149_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1849 VPWR a_19310_11989# a_19237_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1850 VGND a_10443_9813# a_10401_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1851 a_13165_10927# a_12631_10933# a_13070_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1852 a_11785_7663# a_11251_7669# a_11690_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1858 a_17118_9839# a_16679_9845# a_17033_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1859 o_result_ring[4] a_14839_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1861 VPWR a_19735_10651# a_19651_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1864 VPWR a_12500_10357# net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1865 a_14001_8457# net1 w_ring_int_norsz[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1867 VGND w_ring_norsz[10] w_ring_int_norsz[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1868 a_14733_9839# w_ring_buf[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1871 VPWR a_14415_7485# a_14583_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1879 a_16721_10383# a_16677_10625# a_16555_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1882 VGND i_start a_12355_591# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X1885 o_result_ring[14] a_10975_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1886 VGND a_11619_7119# dbg_ring_sig[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1893 a_19360_8041# a_18961_7669# a_19234_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1894 VPWR a_11895_11471# dbg_reset VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1895 VPWR a_13238_10901# a_13165_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1896 VGND a_20211_9839# a_20379_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1900 a_12717_9839# w_ring_norsz[7] a_12633_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1901 a_13323_10058# w_ring_norsz[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1903 a_14545_9845# a_14379_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1905 a_16845_9845# a_16679_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1908 w_ring_norsz[7] w_ring_int_norsz[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1911 r_dly_store_ring[10] a_20471_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1913 a_16013_7119# a_15023_7119# a_15887_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1914 VPWR net7 a_11251_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1918 dbg_ring_sig[0] a_13795_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1919 a_18501_8757# a_18335_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1920 a_9850_9839# a_9411_9845# a_9765_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1922 VPWR w_ring_norsz[11] a_15381_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1924 a_13629_12015# w_ring_buf[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1925 a_19793_8207# w_ring_buf[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1926 a_18413_12335# r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1928 w_ring_buf[8] a_14103_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1929 a_17221_8751# net10 w_ring_int_norsz[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1933 a_11533_9545# w_ring_norsz[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1934 VGND a_9963_8207# dbg_ring_sig[14] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1936 dbg_ring_sig[13] a_9747_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1938 a_13882_11989# a_13714_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1939 net5 a_12355_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X1943 VGND net2 a_20083_10935# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1945 VPWR w_ring_buf[12] a_15115_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1951 a_17133_10383# a_15943_10383# a_17024_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1952 VGND a_15667_7671# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1953 VGND net2 a_15667_7671# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1955 o_result_ring[6] a_10975_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1956 a_10563_8372# w_ring_norsz[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1957 w_ring_norsz[10] w_ring_norsz[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1962 w_ring_norsz[14] net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1965 a_15630_7231# a_15462_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1968 VGND a_12224_9813# net3 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1969 w_ring_norsz[2] net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1970 o_result_ring[5] a_12723_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1974 VPWR a_16495_6575# o_result_ring[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1976 dbg_ring_sig[15] a_12875_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1978 VGND a_13495_10927# a_13663_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1979 dbg_ring_sig[1] a_16771_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1981 VGND a_12115_7663# a_12283_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1990 a_12199_7663# a_11417_7669# a_12115_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1994 VGND a_17199_10357# a_17133_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1995 VGND a_17286_9813# a_17244_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1998 o_result_ring[14] a_10975_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2000 VGND _03_ a_16721_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2005 a_18303_11187# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2010 VGND a_18303_11187# dbg_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2017 VGND a_14103_10927# o_result_ring[15] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2020 a_19878_11837# a_19605_11471# a_19793_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2026 VPWR r_dly_store_ring[5] a_12723_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
R13 g_ring3[13].stg01_12.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2027 dbg_ring_sig[5] a_11619_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2029 a_11329_10927# w_ring_buf[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2031 VPWR a_9839_9269# dbg_ring_sig[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2032 dbg_ring_sig[9] a_19439_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2034 VGND w_ring_buf[2] a_17783_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2035 VGND a_18942_8725# a_18900_9129# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2037 a_15736_11471# a_14655_11471# a_15389_11713# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2038 VGND r_dly_store_ring[1] a_18151_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2040 o_result_ring[12] a_16495_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2042 VPWR a_17378_7637# a_17305_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2046 a_18015_12247# _07_ a_18413_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X2047 VPWR w_ring_norsz[3] a_18703_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2048 a_13795_11445# w_ring_buf[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2050 VPWR a_11895_11471# dbg_reset VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2051 VGND a_20046_11583# a_20004_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2052 a_11141_10933# a_10975_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2059 a_9747_7093# w_ring_buf[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2062 VGND a_18027_8181# dbg_ring_sig[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2064 w_ring_norsz[0] net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2066 o_result_ring[7] a_11863_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2067 a_15243_9839# a_14545_9845# a_14986_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2075 VGND a_19199_8751# a_19367_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2077 VPWR a_15243_9839# a_15411_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2078 dbg_ring_sig[0] a_13795_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2080 a_19693_10383# a_18703_10383# a_19567_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2082 a_17305_7663# a_16771_7669# a_17210_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2084 VGND a_17659_11623# _08_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2085 VPWR net6 a_19439_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2091 VGND a_17803_7637# a_17761_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2092 dbg_ring_sig[6] a_9839_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2093 a_13081_9545# net8 w_ring_int_norsz[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2098 VPWR a_15071_11146# _01_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2099 VGND a_18151_9839# o_result_ring[1] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2100 o_result_ring[5] a_12723_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2102 VGND r_ring_ctr[2] a_18057_12335# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2103 o_result_ring[7] a_11863_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2104 w_ring_buf[12] a_14747_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2106 o_result_ring[8] a_16127_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2110 VPWR a_16771_9295# dbg_ring_sig[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2113 a_13441_12021# a_13275_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2115 a_15377_7119# w_ring_buf[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2116 VGND a_11858_7637# a_11816_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2121 a_16937_7669# a_16771_7669# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2123 a_19142_12015# a_18703_12021# a_19057_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2124 VGND a_20175_10383# o_result_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2127 a_9945_7663# a_9411_7669# a_9850_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2130 dbg_ring_sig[11] a_16863_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2132 o_result_ring[10] a_21279_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2134 a_15433_11471# a_15389_11713# a_15267_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2138 a_18689_8751# w_ring_buf[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2139 VGND a_19567_10749# a_19735_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R14 net16 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2148 a_10310_591# a_10133_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X2149 VGND a_10975_8751# o_result_ring[14] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2152 dbg_ring_sig[5] a_11619_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2165 a_18869_12021# a_18703_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2166 VGND a_19402_7637# a_19360_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2172 VPWR a_16861_11989# a_16751_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2173 dbg_ring_ctr[1] a_19531_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2174 a_10018_9813# a_9850_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2180 dbg_ring_sig[4] a_13735_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2184 VPWR a_14158_7231# a_14085_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2186 VPWR r_dly_store_ring[6] a_10975_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2187 VPWR a_14747_12015# o_result_ring[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2189 VPWR w_ring_buf[9] a_19439_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2190 dbg_ring_sig[7] a_10851_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2192 a_11717_9839# w_ring_norsz[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2193 a_13785_10548# w_ring_norsz[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2194 a_16845_9845# a_16679_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2202 w_ring_int_norsz[1] w_ring_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2204 o_result_ring[9] a_21279_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2205 a_11605_7663# w_ring_buf[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2209 _06_ a_17180_11721# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2220 a_14085_7485# a_13551_7119# a_13990_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2221 w_ring_norsz[14] w_ring_int_norsz[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2223 VPWR a_10975_9839# o_result_ring[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2224 VGND r_dly_store_ring[13] a_10699_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2225 a_10018_8725# a_9850_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
R15 VPWR g_ring3[10].stg01_9.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2229 _07_ r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2232 VPWR r_dly_store_ring[14] a_10975_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2233 _02_ a_18015_12247# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.36 ps=2.72 w=1 l=0.15
X2234 VPWR net7 a_10975_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2235 VPWR a_10275_9839# a_10443_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2236 r_dly_store_ring[4] a_14583_7387# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2241 dbg_ring_sig[11] a_16863_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2242 VGND a_12723_7663# o_result_ring[5] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2244 VPWR a_11391_10548# w_ring_buf[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2245 a_13001_9839# w_ring_int_norsz[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2247 a_10018_8725# a_9850_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2252 VGND w_ring_norsz[7] w_ring_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2254 o_result_ring[10] a_21279_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2256 w_ring_norsz[8] net3 a_13085_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2258 o_result_ctr[0] a_20175_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2260 a_19149_7663# w_ring_buf[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2264 w_ring_int_norsz[2] w_ring_norsz[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2267 VGND a_19310_11989# a_19268_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2268 VGND a_18151_9839# o_result_ring[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2269 VPWR r_dly_store_ring[11] a_18243_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2270 w_ring_int_norsz[9] net15 a_14385_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2271 VPWR a_10975_8751# o_result_ring[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2275 VGND net6 a_18795_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2282 VGND w_ring_norsz[2] w_ring_int_norsz[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2283 VPWR a_10275_8751# a_10443_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2285 o_result_ring[6] a_10975_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2286 VPWR net7 a_13275_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2293 VGND a_16055_7387# a_16013_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2296 a_15279_11837# _04_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2299 VGND net7 a_14379_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2301 a_20303_8573# a_19605_8207# a_20046_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2311 dbg_ring_sig[10] a_18027_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2312 net7 a_9556_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2313 a_9839_9269# w_ring_buf[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2318 a_12897_8751# net1 w_ring_int_norsz[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2319 VPWR a_16495_6575# o_result_ring[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2322 VPWR r_ring_ctr[0] _00_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2323 r_ring_ctr[1] a_15911_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2327 VGND net5 _04_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2330 VGND a_9839_9269# dbg_ring_sig[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2331 net4 a_12500_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2338 a_9577_8757# a_9411_8757# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2340 VGND a_10018_9813# a_9976_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2344 dbg_ring_ctr[1] a_19531_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2347 VGND a_17783_8751# dbg_ring_sig[2] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2349 w_dly_stop[1] a_11343_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2351 VGND a_17383_12319# a_17317_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2355 VPWR a_16863_7119# dbg_ring_sig[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2356 VPWR a_12723_7663# o_result_ring[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2358 a_16751_12015# _05_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2359 VPWR a_16127_9839# o_result_ring[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2360 a_19793_11471# r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2361 VPWR a_19567_10749# a_19735_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2362 a_15971_7485# a_15189_7119# a_15887_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2368 VPWR a_17543_9839# a_17711_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2373 a_16751_12015# a_16127_12021# a_16643_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2374 o_result_ring[0] a_14747_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2378 a_19785_8041# a_18795_7669# a_19659_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2381 a_20303_8573# a_19439_8207# a_20046_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2382 VGND a_21279_8751# o_result_ring[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2387 a_19325_9129# a_18335_8757# a_19199_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2388 VPWR w_ring_norsz[10] a_17221_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2394 w_ring_int_norsz[12] net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2395 w_ring_norsz[8] net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2400 o_result_ring[12] a_16495_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2406 a_11582_10901# a_11414_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2410 VPWR net5 _05_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2412 a_10851_10357# w_ring_buf[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2413 o_result_ring[8] a_16127_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2415 a_13990_7485# a_13551_7119# a_13905_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2416 a_12500_10357# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2419 a_17125_7663# w_ring_buf[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2422 r_dly_store_ring[13] a_10443_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2426 VPWR a_12355_12015# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2429 dbg_ring_sig[3] a_18887_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2430 VGND a_13735_6575# dbg_ring_sig[4] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2438 a_13785_10548# w_ring_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2439 VGND net16 w_ring_int_norsz[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2440 a_15369_10217# a_14379_9845# a_15243_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2444 _00_ r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2446 VPWR w_ring_int_norsz[9] a_14361_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2449 VPWR net4 _03_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2452 a_19651_12015# a_18869_12021# a_19567_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2457 VPWR a_21279_9839# o_result_ring[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2459 a_15389_11713# a_15171_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2461 a_13882_11989# a_13714_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2462 VGND r_dly_store_ctr[1] a_20911_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2464 VPWR a_17783_8751# dbg_ring_sig[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2465 r_dly_store_ring[15] a_13663_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2466 VGND a_16863_7119# dbg_ring_sig[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2467 VPWR a_20471_11739# a_20387_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2468 a_9765_7663# w_ring_buf[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2469 VPWR a_20471_8475# a_20387_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2470 w_ring_norsz[5] w_ring_norsz[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2472 a_12500_10357# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2475 dbg_ring_sig[0] a_13795_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2478 a_15557_7485# a_15023_7119# a_15462_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2484 VPWR r_dly_store_ring[15] a_14103_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2487 a_17635_7663# a_16771_7669# a_17378_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2491 a_15071_11146# _08_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2492 a_14986_9813# a_14818_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2493 VGND w_ring_norsz[9] w_ring_norsz[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2494 VGND a_11391_10548# w_ring_buf[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2497 _04_ net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2498 a_12875_10357# w_ring_buf[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2500 a_13579_10927# a_12797_10933# a_13495_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2503 VGND r_dly_store_ring[9] a_21279_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2507 a_16548_12381# _02_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2510 VPWR a_20911_11471# o_result_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2511 VGND net7 a_11251_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2513 VGND a_16771_9295# dbg_ring_sig[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2514 VPWR a_21279_8751# o_result_ring[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2520 VGND a_15887_7485# a_16055_7387# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2521 a_18774_8751# a_18501_8757# a_18689_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2529 dbg_ring_sig[15] a_12875_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2530 a_14415_7485# a_13717_7119# a_14158_7231# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2533 a_11965_11305# a_10975_10933# a_11839_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2536 a_10359_9839# a_9577_9845# a_10275_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2540 a_17024_10383# a_15943_10383# a_16677_10625# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2543 a_19567_10749# a_18869_10383# a_19310_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2546 a_19513_9845# a_19347_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2547 a_17244_10217# a_16845_9845# a_17118_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2548 r_dly_store_ring[9] a_20379_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2550 a_19701_9839# w_ring_buf[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2552 dbg_ring_sig[15] a_12875_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2560 VGND a_21279_9839# o_result_ring[9] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2561 dbg_ring_sig[3] a_18887_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2562 a_14158_7231# a_13990_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2565 VGND a_15411_9813# a_15369_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2568 VPWR _06_ a_17659_11623# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2569 VPWR a_11619_7119# dbg_ring_sig[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2572 w_ring_norsz[3] net4 a_16673_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2573 VPWR w_ring_norsz[7] a_13081_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2578 VPWR a_17024_10383# a_17199_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2579 VPWR r_dly_store_ring[3] a_20267_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2580 VGND a_18027_8181# dbg_ring_sig[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2584 VPWR a_17803_7637# a_17719_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2586 VGND a_20046_8319# a_20004_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2587 a_19513_9845# a_19347_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2589 VGND w_ring_norsz[9] w_ring_int_norsz[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2593 a_10359_8751# a_9577_8757# a_10275_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2595 a_18165_12015# _07_ _02_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X2597 VPWR a_10018_7637# a_9945_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2598 dbg_ring_sig[8] a_14563_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2606 a_11690_7663# a_11417_7669# a_11605_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2607 w_ring_buf[10] a_17415_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2613 VPWR w_ring_buf[0] a_15943_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2614 a_10379_9460# w_ring_norsz[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2616 VPWR a_18942_8725# a_18869_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2617 VPWR a_19567_12015# a_19735_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2618 VGND a_19567_12015# a_19735_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2619 a_9976_10217# a_9577_9845# a_9850_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2620 w_dly_stop[1] a_11343_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2622 a_13905_7119# w_ring_buf[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2623 a_13238_10901# a_13070_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2624 a_17199_10357# a_17024_10383# a_17378_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2633 dbg_ring_sig[11] a_16863_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2634 a_12241_8041# a_11251_7669# a_12115_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2637 dbg_ring_ctr[2] a_18763_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2642 dbg_ring_sig[6] a_9839_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2645 a_19567_12015# a_18703_12021# a_19310_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2647 VGND w_ring_int_norsz[11] w_ring_norsz[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2648 VGND r_dly_store_ring[4] a_14839_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2651 a_19237_12015# a_18703_12021# a_19142_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2653 a_10593_591# a_10416_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X2654 r_dly_store_ring[15] a_13663_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2655 o_result_ring[7] a_11863_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2656 a_9765_9839# w_ring_buf[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2658 a_19234_7663# a_18961_7669# a_19149_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2660 VPWR a_19531_10927# dbg_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2661 VPWR a_20175_10383# o_result_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2666 dbg_ring_sig[0] a_13795_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2667 VGND a_11895_11471# dbg_reset VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2669 o_result_ring[10] a_21279_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2670 VPWR a_12007_10901# a_11923_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2672 a_14821_11471# a_14655_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2677 w_ring_int_norsz[0] net16 a_11717_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2678 o_result_ring[15] a_14103_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2681 VGND w_ring_buf[12] a_15115_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2684 VPWR net6 a_18335_8757# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2688 VGND a_11619_7119# dbg_ring_sig[5] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2690 a_9577_9845# a_9411_9845# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2692 w_ring_int_norsz[7] w_ring_norsz[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2694 VPWR a_20911_11471# o_result_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2695 VGND a_16495_6575# o_result_ring[12] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2698 VPWR a_12868_11445# _59_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2699 VGND w_dly_stop[2] a_11895_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2702 VGND w_ring_norsz[11] w_ring_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2707 VGND a_11863_10357# o_result_ring[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2708 VGND w_ring_buf[11] a_16863_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2710 a_9765_8751# w_ring_buf[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2713 a_20295_9839# a_19513_9845# a_20211_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2715 o_result_ring[9] a_21279_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2718 VPWR a_16127_9839# o_result_ring[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2720 VGND a_13795_11445# dbg_ring_sig[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2721 dbg_ring_sig[1] a_16771_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2722 a_16293_8751# w_ring_norsz[2] a_16209_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2726 VPWR w_ring_int_norsz[13] a_13257_8457# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2728 VGND net13 w_ring_int_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2734 VPWR a_14307_11989# a_14223_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2735 a_14277_9545# net3 w_ring_norsz[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2737 w_ring_norsz[0] w_ring_int_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2740 VPWR r_ring_ctr[2] a_18165_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.105 ps=1.21 w=1 l=0.15
X2743 a_17262_11721# r_ring_ctr[0] a_17180_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2745 VGND net6 a_19347_9845# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2748 a_16937_7669# a_16771_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2750 a_19793_11471# r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2753 a_13621_11305# a_12631_10933# a_13495_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2754 a_14005_9545# w_ring_norsz[8] a_13921_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2755 VPWR a_19402_7637# a_19329_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2756 w_ring_buf[4] a_13643_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2758 o_result_ring[9] a_21279_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2762 r_dly_store_ring[13] a_10443_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2764 VPWR a_14747_12015# o_result_ring[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2767 VGND a_10275_8751# a_10443_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2769 a_19329_7663# a_18795_7669# a_19234_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2773 dbg_ring_sig[11] a_16863_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2778 VGND w_ring_buf[14] a_9963_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2780 a_19605_11471# a_19439_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2781 a_17199_10357# _03_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2784 o_result_ring[12] a_16495_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2786 w_ring_buf[14] a_9135_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2790 VGND a_20303_11837# a_20471_11739# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2791 VGND r_dly_store_ring[5] a_12723_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2792 VGND w_ring_int_norsz[6] w_ring_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2805 dbg_ring_sig[3] a_18887_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2807 VPWR r_dly_store_ring[12] a_16495_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2808 o_result_ring[10] a_21279_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2815 VPWR w_ring_norsz[5] a_12897_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2818 a_19283_8751# a_18501_8757# a_19199_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2819 a_19057_10383# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2822 a_11582_10901# a_11414_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2823 VPWR net2 a_20083_10935# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2826 r_dly_store_ring[5] a_12283_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2828 dbg_ring_ctr[2] a_18763_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2829 VPWR net7 a_12631_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2830 VPWR net7 a_13551_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2831 a_19786_9839# a_19513_9845# a_19701_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2835 dbg_ring_sig[6] a_9839_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2836 w_ring_norsz[12] w_ring_norsz[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2837 VPWR a_12500_11445# _99_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2838 VPWR a_10851_10357# dbg_ring_sig[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2840 net1 a_12355_591# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X2842 a_15189_7119# a_15023_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2844 a_19268_12393# a_18869_12021# a_19142_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2849 a_15025_8457# w_ring_int_norsz[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2850 VPWR w_ring_norsz[2] a_15841_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2851 VPWR a_19531_10927# dbg_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2852 a_16589_8751# w_ring_int_norsz[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2855 o_result_ring[4] a_14839_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2857 VPWR a_14563_9295# dbg_ring_sig[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2859 a_15630_7231# a_15462_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2860 a_12613_8751# w_ring_norsz[13] a_12529_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2861 VGND a_11895_11471# dbg_reset VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2863 w_ring_int_norsz[5] net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2864 a_17210_7663# a_16937_7669# a_17125_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2873 w_ring_buf[10] a_17415_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2875 o_result_ring[15] a_14103_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2876 a_11329_10927# w_ring_buf[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2880 a_14265_12393# a_13275_12021# a_14139_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2882 a_13323_10058# w_ring_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2883 VPWR r_ring_ctr[1] a_17262_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2886 VPWR w_ring_buf[0] a_14655_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2887 VGND a_10563_8372# w_ring_buf[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2888 _59_.X a_12868_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2892 a_9850_7663# a_9577_7669# a_9765_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2893 a_10379_9460# w_ring_norsz[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2900 a_19786_9839# a_19347_9845# a_19701_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2903 a_12224_9813# net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2906 VGND a_10018_7637# a_9976_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2908 a_11863_10357# r_dly_store_ring[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2909 w_ring_int_norsz[7] net1 a_11809_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2912 a_12868_11445# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2913 dbg_ring_sig[13] a_9747_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2916 a_16109_10383# a_15943_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2917 VPWR a_19954_9813# a_19881_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2920 VPWR net6 a_18703_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2921 dbg_ring_sig[3] a_18887_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2922 VPWR a_16863_7119# dbg_ring_sig[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2924 VPWR a_20175_12015# o_result_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2925 VGND a_21279_8751# o_result_ring[10] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2927 VGND net4 w_ring_norsz[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2928 a_13629_12015# w_ring_buf[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2929 a_17370_12015# a_16293_12021# a_17208_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2931 a_13633_8457# net3 w_ring_norsz[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2932 VGND r_dly_store_ctr[0] a_20175_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2933 a_11759_8372# w_ring_norsz[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2940 net5 a_12355_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X2942 w_ring_int_norsz[13] net12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2949 VGND net7 a_13551_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2952 a_19881_9839# a_19347_9845# a_19786_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2956 a_12868_11445# net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2958 a_15189_7119# a_15023_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2962 o_result_ring[0] a_14747_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2963 _60_.X a_20083_10935# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2968 w_ring_norsz[15] w_ring_int_norsz[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2969 VPWR a_15389_11713# a_15279_11837# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2974 VPWR net6 a_19439_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2975 w_ring_buf[8] a_14103_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2981 VGND a_20175_12015# o_result_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2983 a_19878_11837# a_19439_11471# a_19793_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2985 a_16739_12393# a_16293_12021# a_16643_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2986 a_14818_9839# a_14545_9845# a_14733_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2990 VGND a_14307_11989# a_14265_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2991 a_14545_9845# a_14379_9845# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2992 a_15853_9545# w_ring_int_norsz[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2995 a_13173_8457# net3 w_ring_norsz[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2996 VGND r_dly_store_ring[14] a_10975_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3001 VGND w_ring_buf[4] a_13735_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3002 VPWR a_21279_9839# o_result_ring[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3006 r_dly_store_ring[4] a_14583_7387# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3008 a_17383_12319# a_17208_12393# a_17562_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3018 a_15267_11471# a_14821_11471# a_15171_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3019 VGND w_ring_norsz[12] a_14747_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3021 VGND a_12283_7637# a_12241_8041# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3022 w_ring_buf[9] a_18887_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3023 VPWR a_20303_11837# a_20471_11739# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3024 a_13238_10901# a_13070_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3026 VGND r_ring_ctr[1] a_19531_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3029 o_result_ring[13] a_10699_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3030 a_11839_10927# a_11141_10933# a_11582_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3032 a_11414_10927# a_10975_10933# a_11329_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3033 a_13070_10927# a_12797_10933# a_12985_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3034 dbg_ring_ctr[0] a_18303_11187# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3036 w_ring_buf[14] a_9135_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3040 VGND r_dly_store_ring[11] a_18243_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3046 VGND a_16863_7119# dbg_ring_sig[11] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3047 VPWR a_19310_10495# a_19237_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3048 VGND w_ring_norsz[14] w_ring_norsz[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3051 r_dly_store_ctr[0] a_19735_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3052 VPWR net7 a_9411_7669# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3054 VGND a_16495_6575# o_result_ring[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3055 VGND a_16771_9295# dbg_ring_sig[1] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3056 VPWR a_21279_8751# o_result_ring[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3057 VGND net3 w_ring_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3058 a_9945_9839# a_9411_9845# a_9850_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3059 VPWR a_18151_9839# o_result_ring[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3064 VGND a_19954_9813# a_19912_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3067 VPWR a_13785_10548# w_ring_buf[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3072 a_17659_11623# _07_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X3073 VGND a_14103_10927# o_result_ring[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3075 r_dly_store_ring[11] a_17803_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3079 a_20429_8207# a_19439_8207# a_20303_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3080 VPWR a_14986_9813# a_14913_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3081 VPWR a_9839_9269# dbg_ring_sig[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3082 a_17405_9545# net9 w_ring_int_norsz[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3085 VPWR a_18887_7119# dbg_ring_sig[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3088 w_ring_buf[2] a_17783_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3095 a_10401_9129# a_9411_8757# a_10275_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3097 VPWR a_11582_10901# a_11509_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3098 VGND a_14986_9813# a_14944_10217# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3101 a_16905_12381# a_16861_11989# a_16739_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3102 VGND net6 a_19439_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3103 VGND w_ring_int_norsz[10] w_ring_norsz[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3105 a_9945_8751# a_9411_8757# a_9850_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3108 VGND a_12007_10901# a_11965_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R16 g_ring3[14].stg01_13.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3114 VGND a_10851_10357# dbg_ring_sig[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3115 a_14913_9839# a_14379_9845# a_14818_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3117 w_ring_buf[1] a_16495_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3121 o_result_ctr[2] a_20175_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3124 a_17378_7637# a_17210_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3126 dbg_ring_sig[8] a_14563_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3127 r_dly_store_ring[5] a_12283_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3131 VPWR w_ring_norsz[12] a_13449_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3138 dbg_ring_sig[15] a_12875_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3140 VPWR w_ring_buf[5] a_11619_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3144 o_result_ring[13] a_10699_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3146 a_10401_8041# a_9411_7669# a_10275_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3150 a_17378_10383# _03_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3152 w_ring_buf[11] a_16403_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3154 VPWR a_13882_11989# a_13809_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3155 a_16293_12021# a_16127_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3156 VGND w_ring_norsz[5] w_ring_int_norsz[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3157 o_result_ring[1] a_18151_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3160 w_ring_norsz[9] w_ring_norsz[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3168 VGND r_dly_store_ring[2] a_19991_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3169 w_ring_norsz[14] net3 a_12257_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3178 a_12441_9545# w_ring_norsz[6] a_12357_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3181 VGND a_12875_10357# dbg_ring_sig[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3184 VGND a_17543_9839# a_17711_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3185 a_19659_7663# a_18795_7669# a_19402_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3187 a_15279_11837# a_14655_11471# a_15171_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3192 a_19057_10383# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3195 VGND a_18887_7119# dbg_ring_sig[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3197 VGND a_20471_8475# a_20429_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3199 a_20303_11837# a_19605_11471# a_20046_11583# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3203 a_16567_10749# _03_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3210 a_16548_12381# _02_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
R17 VPWR g_ring3[15].stg01_14.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3214 dbg_ring_ctr[0] a_18303_11187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3218 VPWR net7 a_11343_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3219 a_13495_10927# a_12797_10933# a_13238_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3223 r_dly_store_ring[8] a_15411_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3225 VGND w_ring_norsz[3] w_ring_int_norsz[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3228 r_ring_ctr[2] a_17383_12319# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3233 VGND _05_ a_16905_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3234 r_ring_ctr[0] a_17199_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3235 dbg_ring_ctr[2] a_18763_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3236 VGND net6 a_19439_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3240 w_ring_norsz[7] net3 a_12809_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3249 a_20046_11583# a_19878_11837# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3250 dbg_ring_sig[13] a_9747_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X3253 a_15327_9839# a_14545_9845# a_15243_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3257 a_15462_7485# a_15189_7119# a_15377_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3258 a_14645_8457# net4 w_ring_norsz[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3262 VPWR a_13663_10901# a_13579_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3264 VPWR a_19827_7637# a_19743_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3267 a_17378_7637# a_17210_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3270 w_ring_int_norsz[15] net14 a_11533_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3271 w_ring_int_norsz[1] net1 a_13649_9545# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3273 a_17317_12393# a_16127_12021# a_17208_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3274 VPWR w_ring_buf[3] a_18887_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3276 a_19310_11989# a_19142_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3277 VGND a_13795_11445# dbg_ring_sig[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3278 w_ring_buf[9] a_18887_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3286 VPWR a_10699_7119# o_result_ring[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3287 a_18015_12247# r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.365 ps=1.73 w=1 l=0.15
X3288 VPWR a_11863_10357# o_result_ring[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3290 VPWR a_15887_7485# a_16055_7387# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3291 VPWR a_13795_11445# dbg_ring_sig[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3296 _99_.X a_12500_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3301 VPWR a_15667_7671# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3302 VGND net6 a_18335_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3303 a_12633_9839# w_ring_int_norsz[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3305 VGND a_20911_11471# o_result_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3309 VGND a_13785_10548# w_ring_buf[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3311 VPWR w_ring_buf[0] a_16127_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3312 a_14818_9839# a_14379_9845# a_14733_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3313 w_ring_buf[4] a_13643_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3314 a_17033_9839# w_ring_buf[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3318 VPWR w_ring_norsz[9] a_18887_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3324 a_14139_12015# a_13441_12021# a_13882_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3326 VGND r_dly_store_ring[3] a_20267_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3328 w_ring_buf[2] a_17783_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3330 VPWR a_9556_8181# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3332 VPWR a_15630_7231# a_15557_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3336 dbg_ring_sig[10] a_18027_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3338 VPWR w_ring_buf[8] a_14563_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3339 VGND net4 w_ring_norsz[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3342 w_ring_int_norsz[9] w_ring_norsz[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3343 VGND w_ring_norsz[5] w_ring_norsz[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3347 r_dly_store_ring[11] a_17803_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 i_start VGND 0.76f
C1 i_stop VGND 0.85f
C2 o_result_ring[12] VGND 3.64f
C3 o_result_ring[4] VGND 3.28f
C4 dbg_ring_sig[4] VGND 3.37f
C5 dbg_ring_sig[3] VGND 3.44f
C6 dbg_ring_sig[11] VGND 3.54f
C7 dbg_ring_sig[5] VGND 3.49f
C8 o_result_ring[13] VGND 3.45f
C9 dbg_ring_sig[13] VGND 5.02f
C10 o_result_ring[3] VGND 3.63f
C11 o_result_ring[11] VGND 3.79f
C12 dbg_ring_sig[12] VGND 3.63f
C13 o_result_ring[5] VGND 3.63f
C14 dbg_ring_sig[10] VGND 4.11f
C15 dbg_ring_sig[14] VGND 5.45f
C16 o_result_ring[10] VGND 5.34f
C17 dbg_ring_sig[2] VGND 4.29f
C18 o_result_ring[14] VGND 5.53f
C19 o_result_ring[2] VGND 5.82f
C20 dbg_ring_sig[9] VGND 5.89f
C21 dbg_ring_sig[1] VGND 4.88f
C22 dbg_ring_sig[8] VGND 4.5f
C23 dbg_ring_sig[6] VGND 4.94f
C24 o_result_ring[9] VGND 5.14f
C25 o_result_ring[1] VGND 4.54f
C26 o_result_ring[8] VGND 4.5f
C27 o_result_ring[6] VGND 5.61f
C28 o_result_ctr[0] VGND 4.38f
C29 dbg_ring_sig[15] VGND 4.22f
C30 o_result_ring[7] VGND 6.15f
C31 dbg_ring_sig[7] VGND 5.55f
C32 dbg_ring_ctr[1] VGND 4.17f
C33 dbg_ring_ctr[0] VGND 4.38f
C34 o_result_ring[15] VGND 4.04f
C35 o_result_ctr[1] VGND 5.23f
C36 dbg_ring_ctr[2] VGND 3.83f
C37 dbg_ring_sig[0] VGND 3.92f
C38 o_result_ctr[2] VGND 3.63f
C39 o_result_ring[0] VGND 3.62f
C40 dbg_reset VGND 5.64f
C41 VPWR VGND 2.81p
C42 a_10593_591# VGND 0.227f $ **FLOATING
C43 a_12355_591# VGND 0.698f $ **FLOATING
C44 a_10416_591# VGND 0.498f $ **FLOATING
C45 a_10310_591# VGND 0.578f $ **FLOATING
C46 a_10133_591# VGND 0.5f $ **FLOATING
C47 a_9814_591# VGND 0.535f $ **FLOATING
C48 a_16495_6575# VGND 1.2f $ **FLOATING
C49 a_14839_6575# VGND 1.2f $ **FLOATING
C50 a_13735_6575# VGND 1.2f $ **FLOATING
C51 r_dly_store_ring[12] VGND 0.879f $ **FLOATING
C52 a_15377_7119# VGND 0.23f $ **FLOATING
C53 a_18887_7119# VGND 1.2f $ **FLOATING
C54 a_16863_7119# VGND 1.2f $ **FLOATING
C55 a_15887_7485# VGND 0.609f $ **FLOATING
C56 a_16055_7387# VGND 0.817f $ **FLOATING
C57 a_15462_7485# VGND 0.626f $ **FLOATING
C58 a_15630_7231# VGND 0.581f $ **FLOATING
C59 a_15189_7119# VGND 1.43f $ **FLOATING
C60 a_15023_7119# VGND 1.81f $ **FLOATING
C61 r_dly_store_ring[4] VGND 0.794f $ **FLOATING
C62 a_13905_7119# VGND 0.23f $ **FLOATING
C63 a_14415_7485# VGND 0.609f $ **FLOATING
C64 a_14583_7387# VGND 0.817f $ **FLOATING
C65 a_13990_7485# VGND 0.626f $ **FLOATING
C66 a_14158_7231# VGND 0.581f $ **FLOATING
C67 a_13717_7119# VGND 1.43f $ **FLOATING
C68 a_13551_7119# VGND 1.81f $ **FLOATING
C69 a_11619_7119# VGND 1.2f $ **FLOATING
C70 a_10699_7119# VGND 1.2f $ **FLOATING
C71 a_9747_7093# VGND 1.2f $ **FLOATING
C72 a_19149_7663# VGND 0.23f $ **FLOATING
C73 a_17125_7663# VGND 0.23f $ **FLOATING
C74 w_ring_buf[4] VGND 1.49f $ **FLOATING
C75 a_11605_7663# VGND 0.23f $ **FLOATING
C76 r_dly_store_ring[13] VGND 0.866f $ **FLOATING
C77 a_9765_7663# VGND 0.23f $ **FLOATING
C78 a_20267_7663# VGND 1.2f $ **FLOATING
C79 r_dly_store_ring[3] VGND 0.696f $ **FLOATING
C80 a_19659_7663# VGND 0.609f $ **FLOATING
C81 a_19827_7637# VGND 0.817f $ **FLOATING
C82 a_19234_7663# VGND 0.626f $ **FLOATING
C83 a_19402_7637# VGND 0.581f $ **FLOATING
C84 a_18961_7669# VGND 1.43f $ **FLOATING
C85 a_18795_7669# VGND 1.81f $ **FLOATING
C86 a_18243_7663# VGND 1.2f $ **FLOATING
C87 r_dly_store_ring[11] VGND 0.696f $ **FLOATING
C88 a_17635_7663# VGND 0.609f $ **FLOATING
C89 a_17803_7637# VGND 0.817f $ **FLOATING
C90 a_17210_7663# VGND 0.626f $ **FLOATING
C91 a_17378_7637# VGND 0.581f $ **FLOATING
C92 a_16937_7669# VGND 1.43f $ **FLOATING
C93 a_16771_7669# VGND 1.81f $ **FLOATING
C94 a_15667_7671# VGND 0.648f $ **FLOATING
C95 a_15115_7663# VGND 1.2f $ **FLOATING
C96 w_ring_buf[12] VGND 1.58f $ **FLOATING
C97 a_14747_7663# VGND 0.524f $ **FLOATING
C98 a_13643_7663# VGND 0.524f $ **FLOATING
C99 a_12723_7663# VGND 1.2f $ **FLOATING
C100 r_dly_store_ring[5] VGND 0.696f $ **FLOATING
C101 a_12115_7663# VGND 0.609f $ **FLOATING
C102 a_12283_7637# VGND 0.817f $ **FLOATING
C103 a_11690_7663# VGND 0.626f $ **FLOATING
C104 a_11858_7637# VGND 0.581f $ **FLOATING
C105 a_11417_7669# VGND 1.43f $ **FLOATING
C106 a_11251_7669# VGND 1.81f $ **FLOATING
C107 a_10275_7663# VGND 0.609f $ **FLOATING
C108 a_10443_7637# VGND 0.817f $ **FLOATING
C109 a_9850_7663# VGND 0.626f $ **FLOATING
C110 a_10018_7637# VGND 0.581f $ **FLOATING
C111 a_9577_7669# VGND 1.43f $ **FLOATING
C112 a_9411_7669# VGND 1.81f $ **FLOATING
C113 a_19793_8207# VGND 0.23f $ **FLOATING
C114 a_20303_8573# VGND 0.609f $ **FLOATING
C115 a_20471_8475# VGND 0.817f $ **FLOATING
C116 a_19878_8573# VGND 0.626f $ **FLOATING
C117 a_20046_8319# VGND 0.581f $ **FLOATING
C118 a_19605_8207# VGND 1.43f $ **FLOATING
C119 a_19439_8207# VGND 1.81f $ **FLOATING
C120 w_ring_buf[3] VGND 1.64f $ **FLOATING
C121 w_ring_buf[11] VGND 1.87f $ **FLOATING
C122 w_ring_buf[5] VGND 1.61f $ **FLOATING
C123 w_ring_buf[13] VGND 1.94f $ **FLOATING
C124 a_18703_8207# VGND 0.524f $ **FLOATING
C125 a_18027_8181# VGND 1.2f $ **FLOATING
C126 a_16403_8207# VGND 0.524f $ **FLOATING
C127 w_ring_int_norsz[4] VGND 0.878f $ **FLOATING
C128 w_ring_int_norsz[12] VGND 1.04f $ **FLOATING
C129 w_ring_int_norsz[5] VGND 0.844f $ **FLOATING
C130 w_ring_norsz[12] VGND 2.65f $ **FLOATING
C131 w_ring_int_norsz[13] VGND 0.897f $ **FLOATING
C132 w_ring_norsz[4] VGND 2.81f $ **FLOATING
C133 a_11759_8372# VGND 0.524f $ **FLOATING
C134 a_10563_8372# VGND 0.524f $ **FLOATING
C135 a_9963_8207# VGND 1.2f $ **FLOATING
C136 a_9556_8181# VGND 0.648f $ **FLOATING
C137 a_18689_8751# VGND 0.23f $ **FLOATING
C138 w_ring_buf[10] VGND 2.19f $ **FLOATING
C139 a_21279_8751# VGND 1.2f $ **FLOATING
C140 r_dly_store_ring[10] VGND 1.09f $ **FLOATING
C141 a_19199_8751# VGND 0.609f $ **FLOATING
C142 a_19367_8725# VGND 0.817f $ **FLOATING
C143 a_18774_8751# VGND 0.626f $ **FLOATING
C144 a_18942_8725# VGND 0.581f $ **FLOATING
C145 a_18501_8757# VGND 1.43f $ **FLOATING
C146 a_18335_8757# VGND 1.81f $ **FLOATING
C147 a_17783_8751# VGND 1.2f $ **FLOATING
C148 a_17415_8751# VGND 0.524f $ **FLOATING
C149 net10 VGND 0.822f $ **FLOATING
C150 net11 VGND 1.17f $ **FLOATING
C151 g_ring3[11].stg01_10.HI VGND 0.415f $ **FLOATING
C152 w_ring_norsz[3] VGND 3.89f $ **FLOATING
C153 w_ring_norsz[11] VGND 2.31f $ **FLOATING
C154 w_ring_int_norsz[3] VGND 0.917f $ **FLOATING
C155 w_ring_int_norsz[11] VGND 0.995f $ **FLOATING
C156 g_ring3[12].stg01_11.HI VGND 0.415f $ **FLOATING
C157 g_ring3[13].stg01_12.HI VGND 0.415f $ **FLOATING
C158 net12 VGND 1.27f $ **FLOATING
C159 g_ring3[14].stg01_13.HI VGND 0.415f $ **FLOATING
C160 a_9765_8751# VGND 0.23f $ **FLOATING
C161 w_ring_int_norsz[6] VGND 0.722f $ **FLOATING
C162 w_ring_norsz[5] VGND 2.92f $ **FLOATING
C163 w_ring_int_norsz[14] VGND 0.722f $ **FLOATING
C164 net13 VGND 1.49f $ **FLOATING
C165 w_ring_norsz[13] VGND 3.28f $ **FLOATING
C166 a_10975_8751# VGND 1.2f $ **FLOATING
C167 r_dly_store_ring[14] VGND 0.735f $ **FLOATING
C168 a_10275_8751# VGND 0.609f $ **FLOATING
C169 a_10443_8725# VGND 0.817f $ **FLOATING
C170 a_9850_8751# VGND 0.626f $ **FLOATING
C171 a_10018_8725# VGND 0.581f $ **FLOATING
C172 a_9577_8757# VGND 1.43f $ **FLOATING
C173 w_ring_buf[14] VGND 1.73f $ **FLOATING
C174 a_9411_8757# VGND 1.81f $ **FLOATING
C175 a_9135_8751# VGND 0.524f $ **FLOATING
C176 w_ring_buf[2] VGND 1.52f $ **FLOATING
C177 w_ring_norsz[10] VGND 2.25f $ **FLOATING
C178 a_19991_9295# VGND 1.2f $ **FLOATING
C179 r_dly_store_ring[2] VGND 0.957f $ **FLOATING
C180 a_19439_9295# VGND 1.2f $ **FLOATING
C181 a_18887_9295# VGND 0.524f $ **FLOATING
C182 a_17783_9295# VGND 0.524f $ **FLOATING
C183 w_ring_norsz[2] VGND 2.9f $ **FLOATING
C184 a_16771_9295# VGND 1.2f $ **FLOATING
C185 a_16495_9295# VGND 0.524f $ **FLOATING
C186 w_ring_int_norsz[10] VGND 1.16f $ **FLOATING
C187 net9 VGND 1.79f $ **FLOATING
C188 g_ring3[10].stg01_9.HI VGND 0.415f $ **FLOATING
C189 g_ring3[15].stg01_14.HI VGND 0.415f $ **FLOATING
C190 w_ring_int_norsz[2] VGND 0.839f $ **FLOATING
C191 w_ring_norsz[9] VGND 3.95f $ **FLOATING
C192 w_ring_norsz[1] VGND 2.68f $ **FLOATING
C193 a_14563_9295# VGND 1.2f $ **FLOATING
C194 w_ring_int_norsz[9] VGND 0.897f $ **FLOATING
C195 w_ring_int_norsz[1] VGND 0.722f $ **FLOATING
C196 w_ring_int_norsz[7] VGND 1.02f $ **FLOATING
C197 w_ring_int_norsz[15] VGND 1.14f $ **FLOATING
C198 net1 VGND 8.63f $ **FLOATING
C199 net14 VGND 0.97f $ **FLOATING
C200 w_ring_norsz[14] VGND 3.66f $ **FLOATING
C201 w_ring_norsz[6] VGND 2.98f $ **FLOATING
C202 a_10379_9460# VGND 0.524f $ **FLOATING
C203 a_9839_9269# VGND 1.2f $ **FLOATING
C204 a_19701_9839# VGND 0.23f $ **FLOATING
C205 a_17033_9839# VGND 0.23f $ **FLOATING
C206 net15 VGND 1.44f $ **FLOATING
C207 a_14733_9839# VGND 0.23f $ **FLOATING
C208 a_21279_9839# VGND 1.2f $ **FLOATING
C209 r_dly_store_ring[9] VGND 0.891f $ **FLOATING
C210 a_20211_9839# VGND 0.609f $ **FLOATING
C211 a_20379_9813# VGND 0.817f $ **FLOATING
C212 a_19786_9839# VGND 0.626f $ **FLOATING
C213 a_19954_9813# VGND 0.581f $ **FLOATING
C214 a_19513_9845# VGND 1.43f $ **FLOATING
C215 w_ring_buf[9] VGND 1.67f $ **FLOATING
C216 a_19347_9845# VGND 1.81f $ **FLOATING
C217 a_18151_9839# VGND 1.2f $ **FLOATING
C218 r_dly_store_ring[1] VGND 0.696f $ **FLOATING
C219 a_17543_9839# VGND 0.609f $ **FLOATING
C220 a_17711_9813# VGND 0.817f $ **FLOATING
C221 a_17118_9839# VGND 0.626f $ **FLOATING
C222 a_17286_9813# VGND 0.581f $ **FLOATING
C223 a_16845_9845# VGND 1.43f $ **FLOATING
C224 w_ring_buf[1] VGND 1.58f $ **FLOATING
C225 a_16679_9845# VGND 1.81f $ **FLOATING
C226 a_16127_9839# VGND 1.2f $ **FLOATING
C227 r_dly_store_ring[8] VGND 0.813f $ **FLOATING
C228 a_15243_9839# VGND 0.609f $ **FLOATING
C229 a_15411_9813# VGND 0.817f $ **FLOATING
C230 a_14818_9839# VGND 0.626f $ **FLOATING
C231 a_14986_9813# VGND 0.581f $ **FLOATING
C232 a_14545_9845# VGND 1.43f $ **FLOATING
C233 w_ring_buf[8] VGND 1.55f $ **FLOATING
C234 a_14379_9845# VGND 1.81f $ **FLOATING
C235 a_14103_9839# VGND 0.524f $ **FLOATING
C236 g_ring3[9].stg01_15.HI VGND 0.415f $ **FLOATING
C237 w_ring_norsz[8] VGND 2.57f $ **FLOATING
C238 net8 VGND 1.51f $ **FLOATING
C239 a_13323_10058# VGND 0.524f $ **FLOATING
C240 net3 VGND 6.53f $ **FLOATING
C241 w_ring_int_norsz[8] VGND 0.923f $ **FLOATING
C242 a_12224_9813# VGND 0.648f $ **FLOATING
C243 g_ring2[8].stg01_8.HI VGND 0.415f $ **FLOATING
C244 w_ring_int_norsz[0] VGND 0.987f $ **FLOATING
C245 a_9765_9839# VGND 0.23f $ **FLOATING
C246 w_ring_norsz[15] VGND 2.57f $ **FLOATING
C247 a_10975_9839# VGND 1.2f $ **FLOATING
C248 r_dly_store_ring[6] VGND 0.735f $ **FLOATING
C249 a_10275_9839# VGND 0.609f $ **FLOATING
C250 a_10443_9813# VGND 0.817f $ **FLOATING
C251 a_9850_9839# VGND 0.626f $ **FLOATING
C252 a_10018_9813# VGND 0.581f $ **FLOATING
C253 a_9577_9845# VGND 1.43f $ **FLOATING
C254 w_ring_buf[6] VGND 1.64f $ **FLOATING
C255 a_9411_9845# VGND 1.81f $ **FLOATING
C256 a_19057_10383# VGND 0.23f $ **FLOATING
C257 a_20175_10383# VGND 1.2f $ **FLOATING
C258 r_dly_store_ctr[0] VGND 0.696f $ **FLOATING
C259 a_19567_10749# VGND 0.609f $ **FLOATING
C260 a_19735_10651# VGND 0.817f $ **FLOATING
C261 a_19142_10749# VGND 0.626f $ **FLOATING
C262 a_19310_10495# VGND 0.581f $ **FLOATING
C263 a_18869_10383# VGND 1.43f $ **FLOATING
C264 a_18703_10383# VGND 1.81f $ **FLOATING
C265 stg01_16.HI VGND 0.415f $ **FLOATING
C266 a_16567_10749# VGND 0.168f $ **FLOATING
C267 a_16364_10383# VGND 0.259f $ **FLOATING
C268 a_17024_10383# VGND 0.736f $ **FLOATING
C269 a_17199_10357# VGND 0.971f $ **FLOATING
C270 a_16459_10383# VGND 0.714f $ **FLOATING
C271 a_16677_10625# VGND 0.653f $ **FLOATING
C272 a_16109_10383# VGND 1.57f $ **FLOATING
C273 a_15943_10383# VGND 1.92f $ **FLOATING
C274 net16 VGND 2.03f $ **FLOATING
C275 w_ring_norsz[0] VGND 2.95f $ **FLOATING
C276 a_13785_10548# VGND 0.524f $ **FLOATING
C277 a_12875_10357# VGND 1.2f $ **FLOATING
C278 a_12500_10357# VGND 0.648f $ **FLOATING
C279 a_11863_10357# VGND 1.2f $ **FLOATING
C280 w_ring_norsz[7] VGND 2.9f $ **FLOATING
C281 a_11391_10548# VGND 0.524f $ **FLOATING
C282 a_10851_10357# VGND 1.2f $ **FLOATING
C283 _60_.X VGND 0.226f $ **FLOATING
C284 _00_ VGND 1.44f $ **FLOATING
C285 _03_ VGND 1.68f $ **FLOATING
C286 a_12985_10927# VGND 0.23f $ **FLOATING
C287 r_dly_store_ring[7] VGND 0.932f $ **FLOATING
C288 a_11329_10927# VGND 0.23f $ **FLOATING
C289 a_20083_10935# VGND 0.648f $ **FLOATING
C290 net2 VGND 10.8f $ **FLOATING
C291 a_19531_10927# VGND 1.2f $ **FLOATING
C292 a_18303_11187# VGND 1.2f $ **FLOATING
C293 net4 VGND 7.57f $ **FLOATING
C294 a_15071_11146# VGND 0.524f $ **FLOATING
C295 a_14103_10927# VGND 1.2f $ **FLOATING
C296 r_dly_store_ring[15] VGND 0.696f $ **FLOATING
C297 a_13495_10927# VGND 0.609f $ **FLOATING
C298 a_13663_10901# VGND 0.817f $ **FLOATING
C299 a_13070_10927# VGND 0.626f $ **FLOATING
C300 a_13238_10901# VGND 0.581f $ **FLOATING
C301 a_12797_10933# VGND 1.43f $ **FLOATING
C302 w_ring_buf[15] VGND 1.69f $ **FLOATING
C303 a_12631_10933# VGND 1.81f $ **FLOATING
C304 a_11839_10927# VGND 0.609f $ **FLOATING
C305 a_12007_10901# VGND 0.817f $ **FLOATING
C306 a_11414_10927# VGND 0.626f $ **FLOATING
C307 a_11582_10901# VGND 0.581f $ **FLOATING
C308 a_11141_10933# VGND 1.43f $ **FLOATING
C309 w_ring_buf[7] VGND 1.43f $ **FLOATING
C310 a_10975_10933# VGND 1.81f $ **FLOATING
C311 a_19793_11471# VGND 0.23f $ **FLOATING
C312 a_20911_11471# VGND 1.2f $ **FLOATING
C313 r_dly_store_ctr[1] VGND 0.696f $ **FLOATING
C314 a_20303_11837# VGND 0.609f $ **FLOATING
C315 a_20471_11739# VGND 0.817f $ **FLOATING
C316 a_19878_11837# VGND 0.626f $ **FLOATING
C317 a_20046_11583# VGND 0.581f $ **FLOATING
C318 a_19605_11471# VGND 1.43f $ **FLOATING
C319 a_19439_11471# VGND 1.81f $ **FLOATING
C320 _08_ VGND 1.89f $ **FLOATING
C321 _06_ VGND 0.904f $ **FLOATING
C322 a_15279_11837# VGND 0.168f $ **FLOATING
C323 a_15076_11471# VGND 0.259f $ **FLOATING
C324 a_18763_11445# VGND 1.2f $ **FLOATING
C325 r_ring_ctr[0] VGND 4.45f $ **FLOATING
C326 r_ring_ctr[1] VGND 3.37f $ **FLOATING
C327 a_17659_11623# VGND 0.56f $ **FLOATING
C328 a_17180_11721# VGND 0.502f $ **FLOATING
C329 a_15736_11471# VGND 0.736f $ **FLOATING
C330 a_15911_11445# VGND 0.971f $ **FLOATING
C331 a_15171_11471# VGND 0.714f $ **FLOATING
C332 _04_ VGND 1.61f $ **FLOATING
C333 a_15389_11713# VGND 0.653f $ **FLOATING
C334 a_14821_11471# VGND 1.57f $ **FLOATING
C335 _01_ VGND 1.08f $ **FLOATING
C336 a_14655_11471# VGND 1.92f $ **FLOATING
C337 a_13795_11445# VGND 1.2f $ **FLOATING
C338 _59_.X VGND 0.226f $ **FLOATING
C339 a_12868_11445# VGND 0.648f $ **FLOATING
C340 _99_.X VGND 0.226f $ **FLOATING
C341 a_12500_11445# VGND 0.648f $ **FLOATING
C342 a_11895_11471# VGND 1.2f $ **FLOATING
C343 w_dly_stop[2] VGND 0.681f $ **FLOATING
C344 a_11619_11471# VGND 0.524f $ **FLOATING
C345 w_dly_stop[1] VGND 0.683f $ **FLOATING
C346 a_11343_11471# VGND 0.524f $ **FLOATING
C347 a_19057_12015# VGND 0.23f $ **FLOATING
C348 a_18057_12335# VGND 0.211f $ **FLOATING
C349 a_16751_12015# VGND 0.168f $ **FLOATING
C350 a_16548_12381# VGND 0.259f $ **FLOATING
C351 a_13629_12015# VGND 0.23f $ **FLOATING
C352 net5 VGND 5.54f $ **FLOATING
C353 a_20175_12015# VGND 1.2f $ **FLOATING
C354 r_dly_store_ctr[2] VGND 0.696f $ **FLOATING
C355 a_19567_12015# VGND 0.609f $ **FLOATING
C356 a_19735_11989# VGND 0.817f $ **FLOATING
C357 a_19142_12015# VGND 0.626f $ **FLOATING
C358 a_19310_11989# VGND 0.581f $ **FLOATING
C359 a_18869_12021# VGND 1.43f $ **FLOATING
C360 a_18703_12021# VGND 1.81f $ **FLOATING
C361 net6 VGND 10.5f $ **FLOATING
C362 r_ring_ctr[2] VGND 2.38f $ **FLOATING
C363 _07_ VGND 1.92f $ **FLOATING
C364 a_18015_12247# VGND 0.706f $ **FLOATING
C365 a_17208_12393# VGND 0.736f $ **FLOATING
C366 a_17383_12319# VGND 0.971f $ **FLOATING
C367 a_16643_12393# VGND 0.714f $ **FLOATING
C368 _05_ VGND 1.77f $ **FLOATING
C369 a_16861_11989# VGND 0.653f $ **FLOATING
C370 a_16293_12021# VGND 1.57f $ **FLOATING
C371 _02_ VGND 1.56f $ **FLOATING
C372 a_16127_12021# VGND 1.92f $ **FLOATING
C373 a_14747_12015# VGND 1.2f $ **FLOATING
C374 r_dly_store_ring[0] VGND 0.696f $ **FLOATING
C375 a_14139_12015# VGND 0.609f $ **FLOATING
C376 a_14307_11989# VGND 0.817f $ **FLOATING
C377 a_13714_12015# VGND 0.626f $ **FLOATING
C378 a_13882_11989# VGND 0.581f $ **FLOATING
C379 a_13441_12021# VGND 1.43f $ **FLOATING
C380 w_ring_buf[0] VGND 5.17f $ **FLOATING
C381 a_13275_12021# VGND 1.81f $ **FLOATING
C382 net7 VGND 11.7f $ **FLOATING
C383 a_12355_12015# VGND 0.698f $ **FLOATING
.ends
