* PEX produced on Fri Mar 22 11:45:11 AM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tdc_ring.ext - technology: sky130A

.subckt tdc_ring dbg_delay_stop dbg_dly_sig[0] dbg_dly_sig[11] dbg_dly_sig[13] dbg_dly_sig[2]
+ dbg_dly_sig[4] dbg_dly_sig[5] dbg_dly_sig[6] dbg_dly_sig[7] dbg_dly_sig[8] dbg_dly_sig[9]
+ dbg_ring_ctr[0] dbg_ring_ctr[1] dbg_ring_ctr[2] i_start i_stop o_result_ctr[0] o_result_ctr[2]
+ o_result_ring[0] o_result_ring[10] o_result_ring[12] o_result_ring[13] o_result_ring[14]
+ o_result_ring[15] o_result_ring[2] o_result_ring[5] o_result_ring[8] o_result_ring[7]
+ o_result_ring[4] o_result_ring[1] dbg_dly_sig[10] dbg_dly_sig[15] o_result_ring[9]
+ o_result_ring[6] o_result_ring[11] o_result_ctr[1] o_result_ring[3] dbg_dly_sig[12]
+ dbg_dly_sig[14] dbg_dly_sig[1] dbg_dly_sig[3] dbg_start_pulse VGND VPWR
X0 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 r_dly_store_ring[12] a_24887_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_14082_9661# a_13809_9295# a_13997_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 VPWR clknet_1_1__leaf_i_stop a_22015_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 VGND r_dly_store_ring[0] a_16127_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X16 net3 clknet_2_2__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_22470_7119# a_22155_7271# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X18 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 VPWR clknet_0_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 _04_ a_13054_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 net22 w_dly_sig2_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X30 r_dly_store_ring[2] a_14675_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X31 net7 clknet_2_2__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR net79 _06_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X34 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 o_result_ring[6] a_16127_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X37 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 a_12415_10357# clknet_1_0__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[5] net35 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X40 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X41 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X42 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X44 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X45 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X48 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X49 VPWR a_18795_10927# o_result_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X50 VGND net65 a_24837_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X51 o_result_ring[0] a_16127_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X52 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X53 VPWR clknet_0_w_dly_stop a_14278_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X54 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X57 a_9861_10927# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X58 a_12040_9813# clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X60 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X61 a_22879_10749# a_22181_10383# a_22622_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X62 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[2] net25 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X64 a_12035_6183# a_12131_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X66 VGND clknet_0_w_dly_stop a_11045_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X67 a_22454_10749# a_22015_10383# a_22369_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X69 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X70 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X71 a_23903_9447# a_23999_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X72 a_14909_12533# clknet_0_w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X73 a_17493_9295# net73 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X74 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X75 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X76 net6 clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X77 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X78 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X81 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X83 VPWR a_13059_11187# o_result_ring[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X87 _86_.X a_12040_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X89 a_14457_4399# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X90 a_15427_10927# a_14729_10933# a_15170_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X91 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X92 a_22443_8181# r_dly_store_ring[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X94 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X98 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X99 a_17314_5487# clknet_0_w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X101 VGND a_14462_8181# a_14391_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X102 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X103 VGND clknet_1_0__leaf_i_stop a_9595_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X104 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X105 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X106 VGND clknet_0_w_dly_sig1_n_ana_[11] a_23202_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X107 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X109 VPWR w_dly_sig2_n_ana_[11] net58 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X110 VGND a_13059_11187# o_result_ring[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X114 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[3] net27 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X115 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X117 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X118 a_15925_6031# a_15759_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X119 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X120 VPWR a_17746_8319# a_17673_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X121 a_18773_8181# clknet_0_w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X123 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X124 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X129 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X130 VPWR clknet_2_0__leaf_w_dly_stop net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X131 a_15553_4943# a_14563_4943# a_15427_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X134 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X137 dbg_start_pulse w_strt_pulse_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X138 VPWR clknet_2_3__leaf_w_dly_stop net11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X139 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[12] net63 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X140 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[8] net49 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X142 a_12415_6005# clknet_1_0__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X143 VPWR w_dly_sig1_n_ana_[15] a_16565_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X144 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X145 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[9] net52 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X149 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X150 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X151 a_16210_6575# clknet_0_w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X153 VGND a_21150_10495# a_21108_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X154 VGND clknet_2_0__leaf_w_dly_stop dbg_delay_stop VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X155 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X156 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X157 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X160 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X161 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X162 VPWR a_14250_9407# a_14177_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X164 VGND a_11863_6835# o_result_ring[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X165 VGND net74 a_12539_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X166 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X168 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X170 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X171 o_result_ring[4] a_11863_9011# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X174 VPWR a_14988_12233# a_14998_12137# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X175 VGND clknet_2_3__leaf_w_dly_stop net15 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X177 VGND clknet_0_w_dly_sig1_n_ana_[6] a_18878_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X179 VGND w_dly_sig2_n_ana_[1] net18 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X180 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X181 a_14278_7663# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X182 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X184 a_17673_8573# a_17139_8207# a_17578_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X185 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X190 VGND clknet_0_w_dly_sig1_n_ana_[1] a_16854_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X191 VPWR clknet_0_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X192 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X193 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X196 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X197 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X198 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X199 _03_ a_13743_12131# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X200 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X201 net39 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X202 net40 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X203 a_19047_13335# a_19215_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X205 a_14967_4399# a_14103_4405# a_14710_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X207 o_result_ring[13] a_22995_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X208 VPWR _00_ a_15562_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0672 ps=0.74 w=0.42 l=0.15
X209 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X210 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X211 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X212 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X213 a_13971_8181# a_14255_8181# a_14190_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X215 VPWR a_15170_10901# a_15097_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X216 VGND net46 w_dly_sig2_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X218 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X221 VGND a_17714_12812# r_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X224 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X225 a_24639_9295# a_24419_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X229 w_dly_sig2_n_ana_[7] net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X231 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X232 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X233 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X235 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X236 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X238 a_9849_7093# clknet_0_w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X239 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X240 a_15170_5055# a_15002_5309# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X241 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X244 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X245 net2 clknet_2_2__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X246 a_15002_10927# a_14563_10933# a_14917_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X247 VPWR net29 a_12969_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X248 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X250 a_21270_11471# clknet_0_w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X251 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X252 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X253 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X255 a_21362_9839# clknet_0_w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X256 net53 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X258 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X259 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X260 VGND a_13643_7119# dbg_dly_sig[3] VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X261 o_result_ctr[2] a_23119_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X263 VGND a_18003_8573# a_18171_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X269 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X270 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X272 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X273 a_11045_10901# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X274 VPWR r_dly_store_ring[14] a_22383_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X275 VGND net59 a_25409_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X276 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X279 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X280 a_12622_6005# a_12415_6005# a_12798_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X283 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X284 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X286 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X288 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X289 a_15851_11721# _06_ _01_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X291 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X292 a_13875_8359# a_13971_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X293 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X294 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X295 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X296 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X297 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X298 net61 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X299 VPWR net58 a_9861_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X300 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X301 a_12438_6575# w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X303 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X304 a_24490_9269# a_24290_9569# a_24639_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X305 net49 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X306 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[9] net51 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X309 r_dly_store_ring[6] a_15135_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X311 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X313 VPWR a_18171_9563# a_18087_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X314 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X316 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X317 VPWR a_22443_8181# o_result_ring[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X318 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X319 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X320 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X322 a_19855_13469# a_19635_13481# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X323 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X324 VPWR w_ring_ctr_clk a_17682_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X325 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X326 _08_ r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X327 VGND a_12622_10357# a_12551_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X328 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X329 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X330 a_12771_6031# a_12551_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X331 VGND r_dly_store_ring[10] a_21279_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X332 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X333 VPWR a_22383_9295# o_result_ring[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X334 a_21362_8751# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X335 VPWR net3 w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X337 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X338 VGND a_20322_6549# a_20280_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X340 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X341 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X343 a_19430_11471# clknet_0_w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X345 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X347 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X348 _05_ a_15116_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.229 ps=1.75 w=1 l=0.15
X349 a_11517_11721# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X350 VGND a_12415_10357# a_12422_10657# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X351 o_result_ring[13] a_22995_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X353 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X354 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X356 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X357 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X358 VGND a_11672_10357# dbg_dly_sig[0] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X359 o_result_ring[0] a_16127_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X362 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X364 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X366 a_17118_13103# a_16845_13109# a_17033_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X367 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X370 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X371 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X372 a_24837_9295# a_24283_9269# a_24490_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X375 a_24209_8207# net61 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X377 VGND clknet_0_w_ring_ctr_clk a_20626_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X378 VGND w_ring_ctr_clk a_17682_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X379 VGND clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X380 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X381 net35 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X385 a_19949_13812# _09_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X388 a_16565_11445# w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X389 o_result_ctr[0] a_18795_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X390 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X391 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X392 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X393 VPWR a_11863_6835# o_result_ring[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X394 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X395 a_22493_7485# a_22155_7271# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X397 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X399 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X400 a_12622_6005# a_12422_6305# a_12771_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X401 _00_ a_15575_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X402 a_13059_11187# r_dly_store_ring[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X403 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X404 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X405 VPWR clknet_0_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X406 a_16366_6143# a_16198_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X407 VPWR clknet_1_1__leaf_i_stop a_19715_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X408 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X409 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X410 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X411 VGND a_13059_11187# o_result_ring[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X413 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X414 a_9049_9839# net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X417 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X420 VPWR net6 w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X421 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X423 net58 w_dly_sig2_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X424 VGND w_dly_sig2_n_ana_[3] net26 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X425 VGND clknet_0_w_dly_sig1_n_ana_[4] a_11689_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X426 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X434 VGND w_dly_sig2_n_ana_[7] net42 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X435 dbg_start_pulse w_strt_pulse_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X436 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X437 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X441 VPWR clknet_0_w_dly_stop a_11689_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X443 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[6] net39 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X445 a_18087_8573# a_17305_8207# a_18003_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X447 r_dly_store_ring[9] a_18999_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X448 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X449 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X451 _07_ a_18506_13423# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X453 VPWR a_23989_11471# dbg_ring_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X454 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X455 VGND r_dly_store_ring[2] a_16403_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X456 a_17025_8725# i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X457 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X458 a_14923_12381# a_14350_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.12 ps=1.41 w=0.42 l=0.15
X459 w_dly_sig2_n_ana_[13] clknet_2_1__leaf_w_dly_stop a_10981_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X461 VPWR clknet_0_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X463 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X464 a_15382_8207# w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X465 a_19793_12015# r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X468 a_15562_12393# a_14998_12137# a_15192_12292# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0662 ps=0.735 w=0.42 l=0.15
X469 VPWR clknet_1_1__leaf_i_stop a_17139_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X470 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X473 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X474 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X475 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X476 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X477 VPWR a_23903_9447# r_dly_store_ring[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X478 a_12131_6005# a_12422_6305# a_12373_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X480 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X483 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X484 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X486 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X487 a_14917_10927# net77 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X488 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X489 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X490 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X491 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X492 a_20069_6575# net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X493 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X495 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X497 a_24490_9269# a_24283_9269# a_24666_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X498 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X499 VGND a_16127_5487# o_result_ring[6] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X500 a_22369_10383# r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X501 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X502 VGND a_16916_7637# dbg_dly_sig[15] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X504 a_22465_6895# net14 w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X507 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X511 a_19982_6031# w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X515 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X516 a_12798_10749# a_12551_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X517 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X520 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X522 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X524 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X528 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X529 net77 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X530 a_21362_7663# w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X534 a_18574_6549# a_18406_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X535 _00_ a_15575_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X536 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X537 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X538 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X539 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X541 a_11689_9269# clknet_0_w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X544 a_22671_7119# a_22535_7093# a_22251_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X545 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X549 a_15093_4777# a_14103_4405# a_14967_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X551 a_20626_8207# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X552 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X554 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X556 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X557 a_24666_9661# a_24419_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X559 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X560 VPWR clknet_0_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X562 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X566 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[8] net47 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X567 VPWR a_12415_6005# a_12422_6305# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X568 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X569 a_15185_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X570 a_23202_7663# clknet_0_w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X571 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X572 a_14081_5461# clknet_0_w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X574 VPWR net70 a_11517_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X575 a_13743_12131# a_13551_12375# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X576 o_result_ctr[1] a_21831_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X577 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X578 o_result_ring[14] a_22383_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X579 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X580 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X581 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X582 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X584 _01_ _06_ a_15851_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X585 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X586 net9 clknet_2_2__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X588 VPWR w_dly_sig1_n_ana_[10] a_21362_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X590 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X591 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X592 VPWR clknet_1_0__leaf_i_stop a_15759_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X593 a_20579_6575# a_19715_6581# a_20322_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X595 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X596 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X597 VGND clknet_0_w_dly_sig1_n_ana_[7] a_17038_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X598 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X602 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X603 a_14700_11989# a_14988_12233# a_14923_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.066 ps=0.745 w=0.36 l=0.15
X605 net13 clknet_2_3__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X606 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X607 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X608 o_result_ring[6] a_16127_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X609 a_12438_6575# w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X610 a_18966_11721# r_ring_ctr[1] _06_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X611 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X615 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X616 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X619 VGND a_14103_10927# w_strt_pulse_n VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X620 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X621 a_22535_7093# clknet_1_1__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X622 o_result_ring[15] a_20359_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X623 net16 clknet_2_3__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X624 VGND clknet_0_w_dly_sig1_n_ana_[12] a_18589_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X625 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X626 VPWR a_11987_7671# dbg_dly_sig[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X627 VPWR clknet_0_w_dly_stop a_14278_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X628 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X629 o_result_ring[10] a_21279_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X631 VGND clknet_2_2__leaf_w_dly_stop net4 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X632 VPWR clknet_0_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X634 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X635 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X637 net43 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X638 VPWR a_17286_12695# a_17220_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X641 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X642 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X646 VPWR a_20471_11989# a_20387_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X647 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X648 w_dly_sig1_n_ana_[0] dbg_start_pulse VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X649 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X650 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X651 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X653 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X654 _09_ a_21281_12117# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.13 ps=1.11 w=0.65 l=0.15
X655 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X656 a_24218_9295# a_23903_9447# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X657 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X658 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X659 VGND clknet_0_w_ring_ctr_clk a_20626_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X660 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[11] net60 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X661 VGND net71 a_18049_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X665 net55 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X666 a_18506_13423# r_ring_ctr[0] a_18420_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X667 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X668 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X669 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X673 VPWR clknet_0_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X674 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X675 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X676 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X679 net48 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X680 w_ring_ctr_clk a_13551_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X682 VPWR clknet_0_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X683 w_dly_sig2_n_ana_[3] clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X684 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X685 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X686 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X687 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X688 VGND a_21891_6835# o_result_ring[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X689 a_14250_9407# a_14082_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X690 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X691 a_18786_12559# clknet_0_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X695 a_24837_9295# a_24290_9569# a_24490_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X696 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X697 a_21150_10495# a_20982_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X698 a_21281_12117# _07_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X699 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X700 VGND a_23903_9447# r_dly_store_ring[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X701 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X702 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X704 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X705 VPWR w_dly_sig1_n_ana_[14] a_18773_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X706 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X708 a_16210_6575# clknet_0_w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X709 net26 w_dly_sig2_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X710 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X712 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X716 a_19605_12021# a_19439_12021# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X721 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X722 VGND net66 w_dly_sig2_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X724 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X725 VPWR a_21831_12015# o_result_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X726 VPWR clknet_0_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X727 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X728 a_17305_8207# a_17139_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X732 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X733 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X734 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X736 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X738 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X739 VPWR a_20747_6549# a_20663_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X740 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X741 o_result_ring[8] a_20635_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X742 VPWR clknet_2_3__leaf_w_dly_stop net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X743 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X745 a_19430_10927# w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X746 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X747 VGND clknet_0_w_dly_sig1_n_ana_[10] a_18773_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X749 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X750 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X751 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X752 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X753 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X754 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X758 VGND a_24490_9269# a_24419_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X759 a_22155_7271# a_22251_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X760 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X761 dbg_ring_ctr[0] a_13955_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X762 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X763 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X764 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X765 a_22995_9269# r_dly_store_ring[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X766 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X768 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X769 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X770 VPWR w_dly_sig1_n_ana_[9] a_19982_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X771 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X773 a_17033_12559# _01_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.109 ps=1.36 w=0.42 l=0.15
X774 VGND net1 a_13551_12375# VGND sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X775 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X779 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X782 a_15128_11305# a_14729_10933# a_15002_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X783 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X784 VGND r_ring_ctr[0] a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X786 a_10689_9839# clknet_2_0__leaf_w_dly_stop w_dly_sig2_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X787 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[3] net28 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X788 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[10] net56 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X790 VPWR a_15192_12292# a_15121_12393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X791 a_12040_9813# clknet_2_0__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X792 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X794 a_13997_9295# net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X797 VGND a_22995_9269# o_result_ring[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X798 VPWR a_15427_5309# a_15595_5211# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X799 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X800 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X802 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X803 a_12551_6031# a_12422_6305# a_12131_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X804 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X806 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net80 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X807 net71 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X808 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X809 a_24803_8573# a_24021_8207# a_24719_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X810 VPWR a_19499_13321# a_19506_13225# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X811 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X813 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net76 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X814 VPWR a_14350_11989# r_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X815 a_21362_9839# clknet_0_w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X816 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X818 a_12438_7663# w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X819 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X820 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X822 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X824 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X825 VPWR a_13144_11989# _46_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X826 a_18321_6575# net49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X828 a_18773_9269# w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X830 a_22535_7093# clknet_1_1__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X832 a_14350_11989# a_14700_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X833 a_17038_10927# clknet_0_w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X836 net47 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X837 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[4] net33 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X838 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X841 net15 clknet_2_3__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X842 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X843 VGND net29 a_12969_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X844 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X845 a_23202_9839# clknet_0_w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X846 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X847 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X852 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X854 a_10981_11721# net62 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X855 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X856 VPWR a_22622_10495# a_22549_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X857 a_23999_9269# a_24283_9269# a_24218_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X859 VGND a_19860_7093# dbg_dly_sig[14] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X861 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X862 a_15014_10383# clknet_0_w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X863 VPWR a_21575_10651# a_21491_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X864 a_18773_8181# clknet_0_w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X866 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X867 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X868 a_14507_9661# a_13643_9295# a_14250_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X870 a_18831_6575# a_18133_6581# a_18574_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X871 VPWR r_ring_ctr[1] a_18929_13647# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X872 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X873 w_strt_pulse_n a_14103_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X874 VPWR w_dly_sig1_n_ana_[3] a_12438_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X875 a_19860_7093# net68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X876 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X879 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X880 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X881 VPWR w_dly_sig2_n_ana_[14] net70 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X883 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X884 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X885 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X886 net34 w_dly_sig2_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X887 VGND clknet_0_w_dly_sig1_n_ana_[7] a_17038_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X888 a_21362_8751# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X891 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X892 dbg_dly_sig[15] a_16916_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X893 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X894 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X896 VPWR w_dly_sig1_n_ana_[1] a_15382_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X897 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[10] net55 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X899 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X901 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X905 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net81 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X906 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X907 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X908 VGND r_dly_store_ring[3] a_16127_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X909 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X912 VGND clknet_0_w_dly_sig1_n_ana_[12] a_18589_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X915 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X916 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X917 r_dly_store_ring[9] a_18999_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X918 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X920 VGND w_dly_sig1_n_ana_[15] a_16565_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X921 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X924 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X926 VGND net30 w_dly_sig2_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X927 a_17305_8207# a_17139_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X928 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X930 VPWR clknet_1_0__leaf_w_ring_ctr_clk a_16679_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X931 VPWR a_17714_12812# r_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X932 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X933 a_18506_13423# r_ring_ctr[2] a_18337_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X934 VGND a_23047_10651# a_23005_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X935 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X937 dbg_ring_ctr[0] a_13955_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X938 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X939 VGND clknet_1_0__leaf_i_stop a_16679_13109# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X941 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X942 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[6] net41 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X944 o_result_ring[8] a_20635_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X946 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X947 net74 w_dly_sig2_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X948 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X949 a_18049_13647# net16 w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X950 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X952 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X953 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X959 VPWR net40 a_16679_5495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X961 VGND a_13955_10357# dbg_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X962 VGND r_dly_store_ring[15] a_20359_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X963 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X964 a_9849_8181# clknet_0_w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X967 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X968 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X969 VGND clknet_0_w_dly_sig1_n_ana_[4] a_11689_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X972 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X973 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X975 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X976 a_18786_12559# clknet_0_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X977 VGND clknet_0_w_dly_stop a_20626_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X980 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X981 a_18773_10357# clknet_0_w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X982 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X985 a_12425_9813# clknet_0_w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X986 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X987 a_24389_8573# a_23855_8207# a_24294_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X988 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X990 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X991 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X993 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X994 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X995 net27 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X996 a_22891_7119# a_22671_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X997 VGND clknet_0_w_dly_sig1_n_ana_[11] a_23202_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X998 a_9849_7093# clknet_0_w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X999 VGND clknet_0_w_dly_sig1_n_ana_[13] a_16749_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1000 VPWR a_14675_9563# a_14591_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1001 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1002 VPWR clknet_0_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1003 VPWR a_21831_12015# o_result_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1004 a_11689_8181# clknet_0_w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1005 a_15382_8207# w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1008 VPWR clknet_0_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1009 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1011 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1012 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1013 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1014 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1015 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1016 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1017 net62 w_dly_sig2_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1018 a_14729_10933# a_14563_10933# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1022 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1023 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1024 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1026 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1027 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1029 VGND a_17284_6005# dbg_dly_sig[8] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1030 r_dly_store_ring[14] a_21575_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1031 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1032 net14 clknet_2_3__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1033 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1035 a_20626_12559# clknet_0_w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1036 a_11689_7093# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1038 VPWR clknet_0_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1039 a_16854_10383# clknet_0_w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1040 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1042 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1043 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1044 VGND a_16127_5487# o_result_ring[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1045 VPWR a_18929_13647# dbg_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1048 VGND a_20359_9839# o_result_ring[15] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1049 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1050 VGND a_24719_8573# a_24887_8475# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1051 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1052 _06_ net79 a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1053 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1054 net44 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1056 VPWR a_13696_5461# dbg_dly_sig[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1057 a_14278_7663# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1058 VPWR a_21279_6575# o_result_ring[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1059 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1060 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1061 a_22742_7093# a_22542_7393# a_22891_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1062 a_19215_13335# a_19499_13321# a_19434_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1063 a_12425_8725# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1065 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1066 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1067 VGND net51 a_22097_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1068 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1069 net19 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1071 VPWR net34 a_9309_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1072 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1073 VPWR net7 w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1074 VGND a_18112_6005# dbg_dly_sig[9] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1076 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1077 VGND w_dly_sig1_n_ana_[5] a_14278_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1078 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1079 net59 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1080 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1081 a_24021_8207# a_23855_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1082 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1083 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1084 a_20982_10749# a_20709_10383# a_20897_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1086 a_22369_10383# r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1087 VGND w_dly_sig1_ana_[1] a_14011_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1088 VGND clknet_0_i_stop a_21362_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1089 a_20626_8207# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1091 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1092 VGND a_23356_8181# dbg_dly_sig[12] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1093 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1094 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1097 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1099 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1100 o_result_ctr[2] a_23119_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1102 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1103 a_14809_8207# a_14255_8181# a_14462_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1104 a_23202_7663# clknet_0_w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1105 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1106 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1107 VPWR net65 a_24837_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1108 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1110 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1111 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1113 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1116 VGND clknet_1_0__leaf_w_ring_ctr_clk a_16679_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1117 VGND clknet_1_1__leaf_i_stop a_19715_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1118 VGND a_19706_13380# a_19635_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1122 a_17493_9295# net73 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1123 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1125 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1126 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1127 VPWR a_13054_11445# _04_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X1128 VPWR w_dly_sig2_n_ana_[2] net22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1129 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1131 a_19434_13469# a_19047_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1132 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1133 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1135 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1136 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1137 VGND clknet_2_3__leaf_w_dly_stop net17 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1138 VPWR clknet_1_0__leaf_i_stop a_13643_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1139 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1140 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1142 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1143 a_13713_6005# clknet_0_w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1144 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1145 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1146 a_18929_13647# r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1147 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1149 VPWR a_15170_5055# a_15097_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1150 a_17284_6005# net44 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1152 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1153 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1154 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1155 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1157 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1160 VPWR a_16623_6397# a_16791_6299# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1162 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1163 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1164 a_18878_8751# clknet_0_w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1165 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1166 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1168 w_dly_sig1_n_ana_[6] net35 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1169 VPWR r_dly_store_ring[0] a_16127_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1170 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1171 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1173 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1175 VGND a_15170_10901# a_15128_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1176 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1177 a_18406_6575# a_17967_6581# a_18321_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1179 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1180 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1184 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1185 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1186 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1187 a_14278_6575# w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1189 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1190 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1191 net23 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1192 a_19982_6031# w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1194 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1196 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1197 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1198 a_18112_6005# net48 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1199 a_14931_13103# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1200 VPWR w_dly_strt_ana_[2] a_12263_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1201 VGND clknet_0_w_dly_sig1_n_ana_[12] a_23202_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1203 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[4] net31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1205 r_ring_ctr[1] a_17714_12812# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X1206 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1209 a_22918_7485# a_22671_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1211 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1213 VGND a_13955_10357# dbg_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1214 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1215 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1216 a_22580_10383# a_22181_10383# a_22454_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1217 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1218 a_17284_6005# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1220 a_16749_9813# clknet_0_w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1221 net10 clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1222 a_15511_10927# a_14729_10933# a_15427_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1223 VPWR a_17711_13077# a_17627_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1224 net11 clknet_2_3__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1225 a_14638_8573# a_14391_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1226 VGND a_12035_6183# r_dly_store_ring[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1227 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1229 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1230 a_11425_10633# clknet_2_0__leaf_w_dly_stop w_dly_sig2_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1239 VPWR w_dly_sig1_n_ana_[14] a_18773_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1240 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1241 a_18532_6953# a_18133_6581# a_18406_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1243 VPWR a_21281_12117# _09_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1244 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[2] net24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1245 o_result_ring[5] a_11863_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1246 VPWR a_14156_12533# _88_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1247 a_19878_12015# a_19439_12021# a_19793_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1248 a_21362_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1250 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1251 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1253 a_12539_11471# net74 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1254 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1255 net42 w_dly_sig2_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1256 VPWR a_18703_7119# o_result_ring[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1259 VPWR net8 w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1261 o_result_ring[15] a_20359_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1262 VPWR clknet_0_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1264 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1265 a_18112_6005# net48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1266 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1267 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1268 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1269 VGND clknet_0_w_dly_stop a_14278_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1270 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1271 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[2] net24 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1272 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1273 a_24021_8207# a_23855_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1274 w_dly_sig1_n_ana_[5] net31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1276 o_result_ring[8] a_20635_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1278 net54 w_dly_sig2_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1279 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1280 o_result_ctr[0] a_18795_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1281 VPWR clknet_2_0__leaf_w_dly_stop net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1283 VGND clknet_0_w_dly_sig1_n_ana_[10] a_18773_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1284 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1285 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1286 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1287 VPWR w_dly_sig1_n_ana_[12] a_20613_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1288 net80 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1289 VPWR a_19706_13380# a_19635_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1290 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1293 VPWR a_18831_6575# a_18999_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1294 a_14278_9839# w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1295 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[1] net21 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1296 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1299 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1300 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1303 VPWR net17 a_23119_8759# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1304 VGND clknet_0_w_dly_sig1_n_ana_[13] a_21362_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1305 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1307 a_20626_12559# clknet_0_w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1308 VGND a_21407_10749# a_21575_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1309 VPWR a_18296_7093# _85_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1311 a_18703_11471# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1312 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1314 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1315 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1317 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1319 VPWR net63 w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1322 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1323 VGND a_20359_9839# o_result_ring[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1324 a_24283_9269# clknet_1_1__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1325 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1326 dbg_ring_ctr[1] a_18929_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1327 a_18325_13647# r_ring_ctr[0] _08_ VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1328 VGND a_22995_9269# o_result_ring[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1329 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1331 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1332 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1333 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1334 a_14729_4943# a_14563_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1336 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1340 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1344 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1346 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1348 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1349 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1351 net3 clknet_2_2__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1354 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1355 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1357 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1358 VPWR clknet_0_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1361 VPWR clknet_2_0__leaf_w_dly_stop net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1362 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1367 VGND a_17711_13077# a_17669_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1368 VPWR w_dly_sig2_n_ana_[6] net38 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1370 a_14809_8207# a_14262_8481# a_14462_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1371 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1372 VPWR clknet_0_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1373 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1374 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1376 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1377 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1378 a_23202_9839# clknet_0_w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1380 w_dly_sig2_n_ana_[11] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1381 a_14278_7663# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1384 VGND clknet_0_w_dly_sig1_n_ana_[11] a_21270_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1385 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1386 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1390 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1391 VPWR clknet_0_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1393 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1394 a_20626_4943# clknet_0_w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1395 dbg_dly_sig[10] a_19216_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1399 VPWR r_ring_ctr[2] _08_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1400 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[1] net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1403 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1404 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1405 VPWR w_dly_sig1_n_ana_[3] a_12438_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1407 VPWR a_12622_6005# a_12551_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X1409 VPWR clknet_0_w_dly_stop a_11045_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1410 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1411 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1412 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1414 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1415 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1418 a_13144_11989# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1419 net60 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1420 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1422 a_14710_4373# a_14542_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1424 VPWR a_15116_13103# _05_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1425 VGND clknet_0_w_dly_sig1_n_ana_[4] a_9849_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1427 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1428 a_23356_8181# net60 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1429 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1430 VGND r_ring_ctr[2] a_23989_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1431 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1432 VPWR clknet_0_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1433 a_14190_8207# a_13875_8359# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1434 a_10141_9071# net27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1435 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1436 VGND a_13875_8359# r_dly_store_ring[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1437 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1438 net66 w_dly_sig2_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1439 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1443 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1444 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1445 a_14988_12233# clknet_1_0__leaf_w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1446 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1447 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1452 w_dly_sig1_n_ana_[1] net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1453 VPWR w_dly_sig2_ana_[1] a_11425_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1454 VPWR clknet_0_i_stop a_12425_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1455 a_22671_7119# a_22542_7393# a_22251_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1456 VGND a_18703_7119# o_result_ring[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1458 a_17127_12925# a_16679_12559# a_17033_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1460 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1461 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1462 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1463 dbg_ring_ctr[2] a_23989_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1464 r_dly_store_ring[0] a_15595_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1465 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1466 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1467 VPWR a_18003_8573# a_18171_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1469 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1470 VGND clknet_0_w_dly_stop a_11689_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1471 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1472 a_16854_10383# clknet_0_w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1473 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1475 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1476 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1477 a_19705_5807# net12 w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1481 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[7] net45 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1483 o_result_ring[8] a_20635_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1484 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1485 w_dly_sig2_n_ana_[14] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1486 o_result_ring[4] a_11863_9011# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1487 VPWR clknet_2_2__leaf_w_dly_stop net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1488 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1489 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1491 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1494 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[15] net79 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1495 o_result_ring[10] a_21279_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1496 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1497 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1498 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1500 a_14710_4373# a_14542_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1501 a_24719_8573# a_24021_8207# a_24462_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1504 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1506 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1508 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1509 net37 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1510 VGND a_19584_6005# dbg_dly_sig[11] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1511 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1512 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1513 o_result_ring[9] a_19255_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1515 a_15427_10927# a_14563_10933# a_15170_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1517 o_result_ring[13] a_22995_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1521 VGND r_ring_ctr[1] a_16109_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X1523 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1524 VGND clknet_0_w_dly_stop a_20626_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1525 a_14967_4399# a_14269_4405# a_14710_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1526 r_dly_store_ring[10] a_20747_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1527 a_21362_8751# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1528 a_15097_10927# a_14563_10933# a_15002_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1530 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1531 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1532 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1533 a_13233_12724# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1534 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1536 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1537 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1538 a_21362_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1539 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1542 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1543 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1545 a_17578_9661# a_17305_9295# a_17493_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1546 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1548 _88_.X a_14156_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1549 a_11689_8181# clknet_0_w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1550 a_24462_8319# a_24294_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1551 VPWR w_dly_stop a_14278_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1552 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1553 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1556 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1562 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1563 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1564 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1566 net24 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1567 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[10] net57 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1568 a_20322_6549# a_20154_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1569 a_23089_7119# a_22535_7093# a_22742_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1570 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1571 r_dly_store_ring[2] a_14675_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1572 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1574 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[4] net32 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1576 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1578 a_22181_10383# a_22015_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1579 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1580 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1582 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1583 a_11689_7093# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1584 VPWR clknet_0_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1585 net30 w_dly_sig2_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1586 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1589 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1590 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1593 w_dly_strt_ana_[3] a_12263_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1594 VPWR clknet_0_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1595 net17 clknet_2_3__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1597 w_dly_sig2_ana_[1] w_dly_sig2_n_ana_[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1599 a_18703_11471# r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
X1600 w_dly_sig1_n_ana_[2] net9 a_11337_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1601 _86_.X a_12040_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1602 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1603 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1606 VPWR net2 w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1610 VGND w_dly_sig1_n_ana_[1] a_15382_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1611 a_20303_12015# a_19605_12021# a_20046_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1612 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1614 VGND net81 a_13054_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1615 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1617 a_20046_11989# a_19878_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1618 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1619 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1621 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1622 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1623 dbg_dly_sig[7] a_16679_5495# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1624 VGND r_dly_store_ctr[1] a_21831_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1625 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1626 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1627 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1628 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1629 VGND w_dly_sig1_n_ana_[5] a_14278_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1630 a_11863_6835# r_dly_store_ring[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X1631 VPWR w_dly_sig1_n_ana_[2] a_14278_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1632 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1634 VPWR w_dly_sig1_n_ana_[9] a_19982_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1635 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1637 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1638 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1640 r_ring_ctr[0] a_14350_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.185 ps=1.87 w=0.65 l=0.15
X1642 VGND a_17543_12925# a_17714_12812# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1643 VPWR clknet_0_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1644 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1646 w_dly_sig1_n_ana_[8] net3 a_18053_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1647 a_19584_6005# net56 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1648 VPWR clknet_0_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1649 _87_.X a_23119_8759# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1651 a_17627_12925# a_16845_12559# a_17543_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X1652 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1653 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1656 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1657 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1658 VPWR w_dly_sig1_n_ana_[0] w_dly_sig1_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1661 VGND w_dly_strt_ana_[3] a_13743_12131# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1665 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1666 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1667 net38 w_dly_sig2_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1669 a_14278_9839# w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1670 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1674 VPWR a_11672_7637# dbg_dly_sig[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1675 o_result_ring[11] a_21891_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1677 net46 w_dly_sig2_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1679 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[14] net73 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1680 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1681 net18 w_dly_sig2_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1682 a_16623_6397# a_15759_6031# a_16366_6143# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1683 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1684 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1687 net68 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1688 a_18296_7093# clknet_1_1__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1690 VPWR a_17746_9407# a_17673_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1691 a_18773_9269# w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1692 VGND clknet_2_3__leaf_w_dly_stop net13 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1693 VPWR a_21407_10749# a_21575_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1696 w_dly_sig1_n_ana_[7] net39 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1697 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1698 VPWR a_11863_6835# o_result_ring[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1699 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1700 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net75 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1702 w_dly_sig1_n_ana_[0] net75 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1703 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1704 o_result_ring[9] a_19255_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1705 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1706 a_9493_10633# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1708 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1710 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1712 a_18773_4917# clknet_0_w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1713 r_ring_ctr[1] a_17714_12812# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1714 VPWR w_dly_sig2_n_ana_[10] net54 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1716 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[13] net67 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1717 a_19584_6005# net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1718 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1719 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1720 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1721 VGND a_20635_8751# o_result_ring[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1722 VPWR clknet_0_w_ring_ctr_clk a_14909_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1723 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1725 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1726 a_18773_8181# clknet_0_w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1727 w_dly_sig1_n_ana_[10] net15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1729 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1730 VGND dbg_start_pulse w_dly_sig1_n_ana_[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1731 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1733 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1735 net64 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1736 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1738 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[9] net52 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1739 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1740 a_14278_8751# w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1743 a_17673_9661# a_17139_9295# a_17578_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1746 dbg_dly_sig[12] a_23356_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1748 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1750 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1751 a_18605_4719# net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1753 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1754 VGND a_13955_10357# dbg_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1755 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1756 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1759 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1762 a_14269_4405# a_14103_4405# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1764 VPWR _05_ a_15575_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1765 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1767 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1768 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1769 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1770 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1771 dbg_dly_sig[9] a_18112_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1772 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1773 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1774 a_16623_6397# a_15925_6031# a_16366_6143# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1776 o_result_ring[10] a_21279_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1778 a_13955_10357# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1779 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1780 a_14213_8573# a_13875_8359# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1781 VGND w_dly_sig1_n_ana_[10] a_21362_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1782 net79 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1783 VGND clknet_1_0__leaf_i_stop a_14563_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1784 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1786 a_9849_8181# clknet_0_w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1787 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1789 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1791 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[3] net29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1792 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1793 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1794 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1795 net65 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1797 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1798 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1799 o_result_ring[3] a_16127_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1802 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1804 a_14946_12015# a_14350_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0913 pd=0.855 as=0.122 ps=1.42 w=0.42 l=0.15
X1805 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1806 a_20322_6549# a_20154_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1807 a_12425_9813# clknet_0_w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1808 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1809 VPWR a_16791_6299# a_16707_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1811 a_13997_9295# net21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1812 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1813 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1814 a_10473_9460# w_dly_stop_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1815 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1816 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1817 net12 clknet_2_3__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1818 a_9849_7093# clknet_0_w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1820 VGND clknet_0_w_dly_stop a_14278_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1821 VGND a_22383_9295# o_result_ring[14] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1822 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1823 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1824 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1827 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1830 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1831 VPWR clknet_0_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1832 a_15427_5309# a_14563_4943# a_15170_5055# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1834 VPWR w_dly_sig1_n_ana_[12] a_20613_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1836 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1837 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1838 dbg_dly_sig[0] a_11672_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1840 a_14542_4399# a_14103_4405# a_14457_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1841 net32 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1843 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1845 a_12438_7663# w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1846 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[6] net40 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1849 a_22963_10749# a_22181_10383# a_22879_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1850 VPWR clknet_2_2__leaf_w_dly_stop net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1851 VPWR clknet_0_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1852 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1854 VGND clknet_1_1__leaf_i_stop a_22015_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1855 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1856 VGND w_dly_sig1_n_ana_[4] a_12438_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1857 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1858 VPWR clknet_2_2__leaf_w_dly_stop net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1861 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1862 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1863 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1866 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[14] net71 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1868 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1869 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1870 a_19499_13321# clknet_1_1__leaf_w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1871 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1873 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1875 VPWR a_23119_10927# o_result_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1876 VPWR a_20359_9839# o_result_ring[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1877 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1878 VGND a_22443_8181# o_result_ring[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1883 VGND w_dly_sig1_n_ana_[13] a_19430_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1884 VGND w_dly_sig2_n_ana_[9] net50 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1885 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1886 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1887 VPWR a_21279_6575# o_result_ring[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1888 dbg_dly_sig[2] a_11304_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1889 VGND _05_ a_15575_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1890 a_12425_8725# clknet_0_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1893 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1898 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[14] net72 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1899 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1900 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1901 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1903 a_13054_11445# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.107 ps=1 w=0.42 l=0.15
X1905 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1906 VGND a_22155_7271# r_dly_store_ring[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1907 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1908 VPWR a_20579_6575# a_20747_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1909 a_20579_6575# a_19881_6581# a_20322_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1910 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1912 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1915 a_18421_13647# r_ring_ctr[1] a_18325_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1916 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1921 a_14668_4777# a_14269_4405# a_14542_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1923 VPWR clknet_0_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1924 VPWR a_12040_9813# _86_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1925 VPWR a_20635_8751# o_result_ring[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1928 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1929 VPWR net46 a_9493_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1930 VGND a_11863_9011# o_result_ring[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1931 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1933 VPWR clknet_0_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1934 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1935 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1936 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1937 a_14391_8207# a_14255_8181# a_13971_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1938 a_15170_5055# a_15002_5309# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1939 VGND clknet_0_w_dly_sig1_n_ana_[14] a_15185_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1943 w_dly_sig1_ana_[1] w_dly_sig1_n_ana_[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1944 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1945 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1946 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1947 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1948 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1950 net43 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1951 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1952 VPWR clknet_1_1__leaf_i_stop a_23855_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1953 a_11672_7637# net32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1954 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1955 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1957 a_15192_12292# a_14998_12137# a_15368_12381# VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.0687 ps=0.76 w=0.36 l=0.15
X1958 VPWR a_14103_10927# w_strt_pulse_n VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1959 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1960 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1962 a_20626_4943# clknet_0_w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1963 net57 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1964 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1965 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1966 VGND clknet_0_w_dly_sig1_n_ana_[9] a_21362_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1967 VPWR a_22995_9269# o_result_ring[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1968 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1969 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1973 net69 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1976 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1977 VGND clknet_1_1__leaf_i_stop a_17139_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1978 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1982 a_17286_12695# a_17127_12925# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.149 ps=1.22 w=0.64 l=0.15
X1983 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1984 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1985 VPWR w_ring_ctr_clk a_17682_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1986 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1987 VPWR a_15595_5211# a_15511_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1991 a_21407_10749# a_20709_10383# a_21150_10495# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1992 VGND clknet_1_0__leaf_i_stop a_14103_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1993 a_19433_5807# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1994 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1997 VGND clknet_0_w_dly_sig1_n_ana_[15] a_18786_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1998 VGND a_16127_9839# o_result_ring[0] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1999 VPWR clknet_0_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2000 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2002 net75 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2003 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2004 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2005 a_18087_9661# a_17305_9295# a_18003_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2008 a_10137_9839# clknet_2_0__leaf_w_dly_stop w_dly_sig2_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2009 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2010 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2012 net48 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2014 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2015 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2016 net21 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2017 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2018 VGND a_21891_6835# o_result_ring[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2019 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2021 VPWR clknet_0_w_ring_ctr_clk a_14909_12533# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2023 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2024 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2025 r_dly_store_ring[10] a_20747_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2026 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2027 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2029 o_result_ring[3] a_16127_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2031 a_16845_12559# a_16679_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2032 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2033 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2036 o_result_ring[1] a_13059_11187# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2037 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2038 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2039 a_14255_8181# clknet_1_0__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2040 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2041 VGND a_13955_10357# dbg_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2042 a_14507_9661# a_13809_9295# a_14250_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2043 a_16845_13109# a_16679_13109# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2044 VGND clknet_0_w_dly_stop a_11689_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2045 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2046 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[6] net39 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2047 a_13713_6005# clknet_0_w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2050 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2051 _09_ a_21281_12117# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.151 ps=1.35 w=1 l=0.15
X2052 VPWR w_dly_sig2_n_ana_[15] net74 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2053 VGND net33 a_12969_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2057 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2058 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2060 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2061 a_17224_12559# a_16845_12559# a_17127_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X2062 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2063 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2064 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2065 a_15382_8207# w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2066 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2067 dbg_ring_ctr[0] a_13955_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2069 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2070 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2071 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2074 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2075 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2076 a_13693_18762# i_start VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2078 a_16565_11445# w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2079 a_12539_11471# w_strt_pulse_n w_dly_sig2_n_ana_[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2080 VPWR clknet_0_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2081 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2085 a_24419_9295# a_24290_9569# a_23999_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2086 VGND w_dly_sig1_n_ana_[3] a_12438_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2087 a_14278_6575# w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2089 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2091 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2093 VPWR clknet_1_0__leaf_i_stop a_14563_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2097 a_19430_10927# w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2098 VPWR r_dly_store_ring[6] a_16127_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2099 a_21362_8751# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2100 r_dly_store_ring[8] a_18171_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2102 a_18957_6953# a_17967_6581# a_18831_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2104 w_dly_sig2_n_ana_[4] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2105 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2106 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2107 VPWR a_22742_7093# a_22671_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2108 dbg_start_pulse w_strt_pulse_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X2109 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2111 a_18003_8573# a_17305_8207# a_17746_8319# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2114 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2115 dbg_dly_sig[4] a_11987_7671# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2118 a_19982_6031# w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2120 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2121 a_12425_9813# clknet_0_w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2122 VPWR clknet_0_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2125 VGND a_18999_6549# a_18957_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2126 net36 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2128 VPWR w_dly_sig2_n_ana_[12] net62 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2129 VPWR w_dly_stop a_14278_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2130 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2131 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2136 a_23999_9269# a_24290_9569# a_24241_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2138 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[11] net61 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2140 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2141 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2142 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2143 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2144 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[8] net49 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2146 VGND a_17714_12812# a_17672_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X2147 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2148 a_19973_12015# a_19439_12021# a_19878_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2149 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2150 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2151 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2152 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2153 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2155 a_17314_5487# clknet_0_w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2157 dbg_ring_ctr[1] a_18929_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2158 a_13551_11721# net75 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2159 net45 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2160 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2161 VPWR clknet_0_i_stop a_21362_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2163 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2164 VPWR clknet_0_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2165 VGND clknet_1_1__leaf_i_stop a_23855_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2166 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2167 VPWR clknet_0_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2168 a_22879_10749# a_22015_10383# a_22622_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2169 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2170 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[13] net68 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2172 a_17038_10927# clknet_0_w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2175 VPWR a_18929_13647# dbg_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2176 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2179 a_22549_10749# a_22015_10383# a_22454_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2180 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2181 VPWR a_23119_10927# o_result_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2185 VGND w_dly_sig1_n_ana_[13] a_19430_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2186 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[11] net59 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2187 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2188 a_19635_13481# a_19506_13225# a_19215_13335# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2189 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2192 net50 w_dly_sig2_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2194 VPWR a_11304_9269# dbg_dly_sig[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2195 a_11863_9011# r_dly_store_ring[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2196 VPWR w_dly_sig1_n_ana_[2] a_14278_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2197 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2199 a_13693_18762# i_start VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2201 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2202 net72 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2203 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2204 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2205 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2206 VGND a_17286_13077# a_17244_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2207 VPWR net59 w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2212 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2213 VPWR a_24283_9269# a_24290_9569# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2215 a_17543_13103# a_16845_13109# a_17286_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2216 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2218 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2219 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[15] net78 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2220 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2221 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2222 a_17746_9407# a_17578_9661# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2223 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2225 a_16845_12559# a_16679_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2226 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2227 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2228 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2229 VPWR a_15135_4373# a_15051_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2230 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2231 VPWR clknet_0_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2232 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2233 a_17746_9407# a_17578_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2234 a_24294_8573# a_24021_8207# a_24209_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2235 net2 clknet_2_2__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2236 VPWR a_21891_6835# o_result_ring[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2237 a_17286_13077# a_17118_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2238 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2240 a_14255_8181# clknet_1_0__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2241 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2243 VGND a_21279_6575# o_result_ring[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2244 a_22622_10495# a_22454_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2245 w_dly_sig1_n_ana_[6] net5 a_10417_7983# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2248 VGND a_14988_12233# a_14998_12137# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2251 VGND clknet_0_w_dly_stop a_11045_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2252 VGND a_15595_10901# a_15553_11305# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2253 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2255 VPWR clknet_0_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2256 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2257 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2258 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2260 a_20429_12393# a_19439_12021# a_20303_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2262 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2263 VGND a_23989_11471# dbg_ring_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2264 VGND w_dly_sig1_ana_[1] a_14809_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2266 a_18003_8573# a_17139_8207# a_17746_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2267 VPWR a_14011_7119# dbg_dly_sig[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2269 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2270 VGND a_16127_7663# o_result_ring[3] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2273 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2276 a_10473_9460# w_dly_stop_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2279 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2280 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[6] net41 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2283 o_result_ring[7] a_18703_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2285 dbg_ring_ctr[2] a_23989_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2286 VGND clknet_0_w_dly_sig1_n_ana_[4] a_9849_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2287 net61 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2288 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2289 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2290 a_14278_7663# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2292 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2294 VPWR a_24719_8573# a_24887_8475# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2296 VGND a_16127_9839# o_result_ring[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2297 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2298 a_12425_8725# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2299 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2300 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2304 a_19457_13103# a_19047_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2305 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2306 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2307 a_11045_10901# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2308 a_17305_9295# a_17139_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2309 a_20613_9269# w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2311 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[2] net25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2315 a_14156_12533# dbg_start_pulse VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2318 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2319 a_17682_12015# w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2320 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2322 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2323 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2324 VGND w_dly_sig2_n_ana_[5] net34 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2325 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2330 o_result_ring[1] a_13059_11187# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2331 VGND a_18795_10927# o_result_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2332 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2333 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2334 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2335 net35 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2339 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2341 VGND w_dly_sig1_ana_[1] a_11241_10159# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2342 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2343 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2344 a_21891_6835# r_dly_store_ring[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2345 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2346 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2347 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2348 VGND net55 a_22465_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2351 o_result_ring[1] a_13059_11187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2354 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2355 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2356 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2357 o_result_ring[12] a_22443_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2358 net25 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2359 VPWR a_12035_6183# r_dly_store_ring[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2360 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2361 dbg_dly_sig[3] a_13643_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2364 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[3] net27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2367 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2369 VGND a_16403_8751# o_result_ring[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2371 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2372 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2374 a_14082_9661# a_13643_9295# a_13997_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2376 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2377 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2378 VGND _08_ a_21436_12375# VGND sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0536 ps=0.675 w=0.42 l=0.15
X2379 a_23989_11471# r_ring_ctr[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2380 VGND r_dly_store_ctr[0] a_18795_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2381 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2382 o_result_ring[9] a_19255_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2383 VGND w_dly_sig1_n_ana_[9] a_19982_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2384 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2385 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2386 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2387 w_dly_sig2_n_ana_[0] w_strt_pulse_n a_12539_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2388 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2389 VPWR a_24462_8319# a_24389_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2390 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2391 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2392 VPWR w_dly_sig2_n_ana_[7] net42 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2393 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2394 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2395 o_result_ring[3] a_16127_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2396 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2398 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2400 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2401 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2403 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2404 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2409 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2410 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2412 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2413 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2414 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net80 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2415 a_14646_7119# clknet_0_w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2416 dbg_start_pulse w_strt_pulse_n VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2417 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2418 net81 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2419 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2420 net63 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2422 VPWR clknet_0_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2423 VGND a_12415_6005# a_12422_6305# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2424 VGND a_20579_6575# a_20747_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2425 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[11] net60 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2427 a_14611_8207# a_14391_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2428 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2430 VGND clknet_2_2__leaf_w_dly_stop net9 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2431 a_13696_5461# net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2433 _03_ a_13743_12131# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X2434 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[13] net69 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2435 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2437 a_20004_12393# a_19605_12021# a_19878_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2438 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2441 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2442 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2444 a_12373_10749# a_12035_10535# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2445 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2446 a_17578_8573# a_17139_8207# a_17493_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2447 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2448 VGND a_20471_11989# a_20429_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2449 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2450 a_14208_9295# a_13809_9295# a_14082_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2453 a_17543_12925# a_16679_12559# a_17286_12695# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2454 VGND clknet_1_0__leaf_i_stop a_15759_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2455 a_18133_6581# a_17967_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2456 VGND w_dly_sig1_n_ana_[4] a_12438_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2458 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2460 VPWR net66 a_11241_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2461 a_12035_10535# a_12131_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2462 net15 clknet_2_3__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2463 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2464 a_16486_7119# w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2466 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2468 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2469 a_19860_7093# net68 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2470 VGND a_14011_7119# dbg_dly_sig[1] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2472 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2473 net4 clknet_2_2__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2475 VPWR a_20359_9839# o_result_ring[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2478 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2479 a_19154_7663# w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2481 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2482 o_result_ring[7] a_18703_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2484 VPWR a_16127_7663# o_result_ring[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2486 VGND r_dly_store_ctr[2] a_23119_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2487 dbg_ring_ctr[0] a_13955_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2488 dbg_delay_stop clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2489 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2490 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2492 a_20613_9269# w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2493 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2494 VGND r_ring_ctr[1] a_18929_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2496 VPWR _02_ a_20053_13481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2497 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2498 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2500 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2501 a_14462_8181# a_14262_8481# a_14611_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2502 a_12969_10383# a_12415_10357# a_12622_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2503 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2504 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2506 VGND net42 w_dly_sig2_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2507 a_12551_10383# a_12422_10657# a_12131_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2508 a_11337_9071# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2510 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2516 VGND net54 w_dly_sig2_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2517 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2518 a_17704_8207# a_17305_8207# a_17578_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2519 a_19430_11471# clknet_0_w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2520 VGND clknet_0_w_dly_sig1_n_ana_[14] a_15185_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2521 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2522 VGND w_dly_sig1_n_ana_[1] a_15382_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2523 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2524 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[10] net55 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2525 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2526 VGND a_14250_9407# a_14208_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2529 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2530 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2531 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2532 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2533 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2537 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2538 net78 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2539 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2541 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2543 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[9] net51 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2546 net9 clknet_2_2__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2548 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2550 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2551 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2552 a_11672_10357# net76 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2553 VPWR a_22995_9269# o_result_ring[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2555 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2556 a_25409_9071# net13 w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2565 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2567 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2568 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2570 VPWR net80 a_15116_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.75 as=0.0609 ps=0.71 w=0.42 l=0.15
X2571 a_20053_13481# a_19499_13321# a_19706_13380# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2572 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2574 dbg_ring_ctr[2] a_23989_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2575 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2578 net13 clknet_2_3__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2580 VGND w_dly_sig2_n_ana_[13] net66 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2581 VPWR a_13875_8359# r_dly_store_ring[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2583 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2584 o_result_ring[9] a_19255_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2585 a_15562_12393# a_14988_12233# a_15192_12292# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2587 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2588 VPWR r_ring_ctr[1] a_15851_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X2589 a_14278_9839# w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2590 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2592 VPWR a_16403_8751# o_result_ring[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2593 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2596 a_21270_11471# clknet_0_w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2598 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2599 VGND a_17746_8319# a_17704_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2600 VGND a_14967_4399# a_15135_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2601 a_18129_9295# a_17139_9295# a_18003_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2603 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2604 VGND a_23989_11471# dbg_ring_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2605 a_9849_8181# clknet_0_w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2606 a_20337_7093# w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2607 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2608 VGND r_ring_ctr[0] a_13955_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2609 VPWR clknet_1_1__leaf_i_stop a_20543_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2610 a_11689_9269# clknet_0_w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2611 o_result_ring[3] a_16127_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2614 r_dly_store_ring[0] a_15595_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2615 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2616 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2617 VGND clknet_0_w_dly_sig1_n_ana_[7] a_17314_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2620 a_17682_12015# w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2625 a_14081_5461# clknet_0_w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2626 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2627 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2631 a_11672_10357# net76 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2632 a_22742_7093# a_22535_7093# a_22918_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2633 VGND a_18795_10927# o_result_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2634 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2635 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2638 a_17213_13103# a_16679_13109# a_17118_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2639 a_18773_4917# clknet_0_w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2640 net51 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2641 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2645 a_15851_11721# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2646 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2647 a_11689_8181# clknet_0_w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2648 a_15382_8207# w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2649 VPWR a_22988_8181# dbg_dly_sig[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2652 a_21362_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2653 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2655 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2659 a_14462_8181# a_14255_8181# a_14638_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2660 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2663 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2664 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2665 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2666 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2667 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2668 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2670 a_15368_12381# a_15121_12393# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.149 ps=1.22 w=0.42 l=0.15
X2671 VGND w_dly_sig1_n_ana_[3] a_12438_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2672 a_14278_8751# w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2673 net76 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2674 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2675 VGND clknet_0_w_dly_sig1_n_ana_[1] a_12425_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2676 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2678 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2680 VGND clknet_0_w_dly_sig1_n_ana_[6] a_13713_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2683 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2684 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2685 VGND a_18929_13647# dbg_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2686 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2687 a_14081_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2688 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2689 a_18773_10357# clknet_0_w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2691 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2692 VPWR clknet_0_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2693 VPWR a_17286_13077# a_17213_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2694 VPWR clknet_0_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2696 o_result_ring[10] a_21279_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2699 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net77 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2700 VGND clknet_1_0__leaf_i_stop a_13643_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2701 VGND clknet_0_i_stop a_12425_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2704 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2705 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2706 a_13551_12375# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X2707 dbg_start_pulse w_strt_pulse_n VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X2708 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2712 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2713 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2714 a_17314_5487# clknet_0_w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2715 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2717 a_17314_7663# w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2718 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2721 net31 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2722 VGND w_dly_sig2_n_ana_[4] net30 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2723 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2727 a_16109_11471# r_ring_ctr[0] _01_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X2729 VGND w_dly_sig2_n_ana_[0] w_dly_sig2_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2730 VGND a_12040_9813# _86_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2731 VPWR clknet_0_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2732 VPWR r_dly_store_ring[8] a_20635_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2734 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2735 VPWR a_16916_7637# dbg_dly_sig[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2736 w_dly_sig1_n_ana_[11] net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2738 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2740 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2741 VGND net57 a_23089_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2742 a_17493_8207# net45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2743 VGND _04_ a_13551_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2744 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2745 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2746 VGND a_20747_6549# a_20705_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2747 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2748 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2749 VPWR a_12035_10535# r_dly_store_ring[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2750 a_14909_12533# clknet_0_w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2751 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2753 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2755 a_20626_4943# clknet_0_w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2756 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2757 a_18878_8751# clknet_0_w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2758 VPWR r_dly_store_ring[9] a_19255_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2760 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2762 VGND a_14350_11989# r_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X2764 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2765 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2767 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2768 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2769 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2771 VPWR clknet_2_0__leaf_w_dly_stop dbg_delay_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2772 VPWR a_24490_9269# a_24419_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2773 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2774 a_13233_12724# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2777 a_13713_6005# clknet_0_w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2778 a_18915_6575# a_18133_6581# a_18831_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2782 a_18929_13647# r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2783 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2786 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2787 VGND a_18171_9563# a_18129_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2788 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2789 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2790 VPWR a_21150_10495# a_21077_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2791 a_18589_9813# clknet_0_w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2792 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2794 w_dly_sig2_n_ana_[0] net74 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2795 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2797 VPWR net33 a_12969_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2798 w_dly_sig2_n_ana_[8] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2799 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2800 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2801 VGND a_22443_8181# o_result_ring[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2802 VGND a_15135_4373# a_15093_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2804 VGND w_dly_sig2_n_ana_[8] net46 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2805 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2806 o_result_ctr[2] a_23119_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2807 VPWR w_dly_sig2_n_ana_[1] net18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2808 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2809 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2812 VPWR clknet_0_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2813 VPWR clknet_0_i_stop a_12425_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2814 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2816 a_22251_7093# a_22542_7393# a_22493_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2818 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2819 o_result_ring[2] a_16403_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2821 a_17033_13103# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2824 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2825 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2826 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2827 r_dly_store_ring[14] a_21575_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2828 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2829 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2830 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2831 VGND net34 w_dly_sig2_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2832 VPWR a_19255_7119# o_result_ring[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2833 a_19982_6031# w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2834 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2835 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2837 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2838 a_17038_10927# clknet_0_w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2839 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2840 VPWR a_14011_7119# dbg_dly_sig[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2841 a_12969_10383# a_12422_10657# a_12622_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2842 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2843 VGND a_16127_7663# o_result_ring[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2846 VGND _03_ a_14103_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2848 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[4] net33 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2849 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2850 net47 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2852 VPWR a_17714_12812# r_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X2853 a_14917_4943# net25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2857 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2858 w_dly_stop_ana_[1] a_9595_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2860 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2861 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2864 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2867 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2869 VPWR clknet_0_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2871 a_21270_11471# clknet_0_w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2872 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2873 VPWR clknet_2_2__leaf_w_dly_stop net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2875 a_15002_5309# a_14563_4943# a_14917_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2876 a_17669_13481# a_16679_13109# a_17543_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2877 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[12] net64 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2878 net37 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2880 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2882 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2883 VGND w_dly_sig1_n_ana_[2] a_14278_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2884 VGND a_19499_13321# a_19506_13225# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2887 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2888 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2889 a_13955_10357# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2890 net56 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2891 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2892 a_24283_9269# clknet_1_1__leaf_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2893 net28 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2895 VPWR clknet_2_3__leaf_w_dly_stop net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2896 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2897 a_14391_8207# a_14262_8481# a_13971_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2899 a_12438_6575# w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2900 a_18420_13423# r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2901 a_15014_10383# clknet_0_w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2903 a_18337_13103# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2904 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2905 VPWR w_dly_sig1_n_ana_[6] a_16486_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2906 VPWR a_22535_7093# a_22542_7393# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2907 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2908 w_dly_sig1_n_ana_[3] net8 a_9589_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2911 VGND clknet_0_w_dly_sig1_n_ana_[12] a_23202_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2912 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2914 o_result_ring[15] a_20359_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2915 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2916 o_result_ring[12] a_22443_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2918 VPWR w_dly_sig1_n_ana_[8] a_19154_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2919 a_21362_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2920 VPWR clknet_0_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2922 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[7] net44 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2924 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2927 VGND clknet_0_w_dly_sig1_n_ana_[15] a_18786_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2928 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2930 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2931 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2934 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2935 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2937 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2939 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2940 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2941 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2943 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[9] net53 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2944 VPWR a_16679_5495# dbg_dly_sig[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2946 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2948 VGND a_13233_12724# w_dly_strt_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2949 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[12] net65 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2950 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2952 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2953 VGND a_18296_7093# _85_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2954 net20 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2955 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2956 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2961 o_result_ctr[1] a_21831_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2962 a_19430_11471# clknet_0_w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2963 a_14081_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2964 a_15185_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2965 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2966 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2967 VGND clknet_0_w_dly_sig1_n_ana_[8] a_18773_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2970 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2971 dbg_dly_sig[14] a_19860_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2972 dbg_ring_ctr[1] a_18929_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2973 a_16916_7637# net72 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2977 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2979 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2980 VGND a_11863_6835# o_result_ring[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2982 dbg_ring_ctr[1] a_18929_13647# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2985 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2986 VPWR a_11672_10357# dbg_dly_sig[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2987 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2992 VPWR w_dly_sig1_n_ana_[11] a_20337_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2994 a_14278_8751# w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2995 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2996 VPWR clknet_0_w_ring_ctr_clk a_20626_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2997 w_dly_sig2_n_ana_[10] clknet_2_1__leaf_w_dly_stop a_10337_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3000 VGND clknet_0_w_dly_sig1_n_ana_[1] a_16854_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3001 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3003 a_14700_11989# a_14998_12137# a_14946_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0913 ps=0.855 w=0.42 l=0.15
X3004 net22 w_dly_sig2_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3005 net5 clknet_2_2__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3006 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3009 VGND a_21831_12015# o_result_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3010 _04_ a_13054_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3011 a_14278_9839# w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3012 a_22988_8181# net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3013 a_16565_11445# w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3015 VGND a_23119_8759# _87_.X VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3018 VGND net70 w_dly_sig2_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3019 a_18703_11471# net79 _06_ VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3020 VGND w_dly_strt_ana_[2] a_12263_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3021 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3022 a_13809_9295# a_13643_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3024 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3025 VGND a_19255_7119# o_result_ring[9] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3027 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3028 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3029 a_16486_7119# w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3032 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3033 dbg_dly_sig[13] a_22988_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3034 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3035 VPWR net18 a_10689_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3036 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3037 o_result_ring[2] a_16403_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3038 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3039 VGND a_14011_7119# dbg_dly_sig[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3042 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3044 o_result_ring[11] a_21891_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3045 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3046 a_15427_5309# a_14729_4943# a_15170_5055# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3049 VGND clknet_0_w_dly_sig1_n_ana_[3] a_9849_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3051 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3052 VPWR a_22155_7271# r_dly_store_ring[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3053 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3054 VPWR w_dly_sig2_n_ana_[3] net26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3055 VPWR clknet_0_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3056 VPWR a_16127_7663# o_result_ring[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3058 a_14909_12533# clknet_0_w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3059 a_16749_6031# a_15759_6031# a_16623_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3061 r_ring_ctr[0] a_14350_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X3062 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3063 net14 clknet_2_3__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3064 VGND r_ring_ctr[2] a_18421_13647# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3065 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3066 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3067 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3072 a_16581_4943# net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3073 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3074 VGND clknet_0_w_dly_sig1_n_ana_[5] a_14081_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3075 a_20053_13481# a_19506_13225# a_19706_13380# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3076 _46_.X a_13144_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3077 a_20897_10383# net69 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3079 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[2] net23 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3082 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3083 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3084 a_14350_11989# a_14700_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.162 ps=1.33 w=1 l=0.15
X3085 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3087 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3088 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3089 VPWR a_18003_9661# a_18171_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3090 net8 clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3091 a_14457_4399# net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3093 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3094 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3095 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3096 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3097 VGND clknet_0_w_dly_sig1_n_ana_[2] a_11689_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3099 a_18773_4917# clknet_0_w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3100 VGND a_13696_5461# dbg_dly_sig[6] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X3101 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3102 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3103 VGND a_20635_8751# o_result_ring[8] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3106 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3107 a_24719_8573# a_23855_8207# a_24462_8319# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3110 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3111 w_dly_stop a_9871_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3113 VPWR a_12622_10357# a_12551_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3114 VGND a_21279_6575# o_result_ring[10] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3116 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3117 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3118 VGND clknet_2_0__leaf_w_dly_stop net10 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3119 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3120 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3122 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3123 a_12438_7663# w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3125 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3127 VGND w_dly_sig1_n_ana_[15] a_16565_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3128 VGND clknet_2_3__leaf_w_dly_stop net11 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3129 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[12] net63 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3130 VPWR a_19216_6005# dbg_dly_sig[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3131 o_result_ring[4] a_11863_9011# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3133 VGND a_22535_7093# a_22542_7393# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3134 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3135 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3136 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3139 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3141 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3142 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3143 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3144 net33 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3145 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3146 w_dly_sig2_n_ana_[6] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3147 a_11672_7637# net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3148 net70 w_dly_sig2_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3149 VPWR clknet_1_1__leaf_i_stop a_19439_12021# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3150 dbg_dly_sig[15] a_16916_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3155 a_16210_6575# clknet_0_w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3158 a_11241_10159# net10 w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3159 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3161 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[15] net79 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3162 a_21533_10383# a_20543_10383# a_21407_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3163 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3164 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3166 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3167 a_12425_8725# clknet_0_i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3168 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3170 dbg_dly_sig[8] a_17284_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3171 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3172 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3173 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3175 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3176 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3177 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3178 a_11689_9269# clknet_0_w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3180 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3181 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3182 VGND a_15192_12292# a_15121_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0989 ps=0.995 w=0.64 l=0.15
X3185 VGND clknet_0_w_dly_sig1_n_ana_[7] a_17314_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3186 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3188 a_13144_11989# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3189 VPWR w_dly_sig1_n_ana_[7] a_17314_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3192 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3194 a_14917_4943# net25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3195 a_14081_5461# clknet_0_w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3198 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3199 a_12035_10535# a_12131_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3200 VGND a_18003_9661# a_18171_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3202 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3203 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3208 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3210 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3211 dbg_dly_sig[5] a_11672_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3214 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3215 VGND clknet_0_w_dly_sig1_n_ana_[13] a_16749_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3217 a_11689_8181# clknet_0_w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3218 a_18133_6581# a_17967_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3219 a_18589_9813# clknet_0_w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3220 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3221 r_dly_store_ring[7] a_16791_6299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3224 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3225 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3226 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3228 VGND clknet_0_w_dly_sig1_n_ana_[9] a_20626_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3229 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3230 VPWR clknet_0_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3233 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3235 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3236 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3238 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3239 VGND net26 w_dly_sig2_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3240 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3242 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3243 VGND r_dly_store_ring[14] a_22383_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3244 VPWR a_24887_8475# a_24803_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3245 net41 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3246 VGND clknet_0_w_dly_sig1_n_ana_[6] a_13713_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3249 a_9861_9839# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3250 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3251 VGND clknet_2_2__leaf_w_dly_stop net3 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3252 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3253 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3254 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3255 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3256 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3259 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3260 net27 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3261 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3262 VGND _06_ _01_ VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3263 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3265 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3266 VGND a_16791_6299# a_16749_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3267 o_result_ring[11] a_21891_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3268 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3269 VGND a_18831_6575# a_18999_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3272 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3274 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3275 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3277 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3278 VGND a_16403_8751# o_result_ring[2] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3279 a_14646_7119# clknet_0_w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3281 VPWR net11 w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3283 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3284 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3285 a_12131_10357# a_12415_10357# a_12350_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3286 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3287 a_23089_7119# a_22542_7393# a_22742_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3288 VPWR a_18929_13647# dbg_ring_ctr[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3289 w_dly_sig1_n_ana_[0] dbg_start_pulse a_13551_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3290 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3292 VGND w_dly_sig1_n_ana_[9] a_19982_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3295 VPWR w_dly_sig1_n_ana_[13] a_19430_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3296 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3297 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3298 a_17314_7663# w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3303 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3304 dbg_dly_sig[1] a_14011_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3306 VPWR clknet_0_w_ring_ctr_clk a_20626_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3307 VGND a_20046_11989# a_20004_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3308 VPWR a_20635_8751# o_result_ring[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3309 VPWR r_dly_store_ctr[1] a_21831_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3310 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3311 clknet_1_0__leaf_i_stop a_12425_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3312 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3313 VGND a_21831_12015# o_result_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3314 w_dly_stop_ana_[1] a_9595_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3316 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3317 o_result_ring[15] a_20359_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3318 VPWR r_dly_store_ring[15] a_20359_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3319 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3320 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3321 a_18296_7093# clknet_1_1__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3322 VPWR r_dly_store_ring[10] a_21279_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3323 w_dly_sig2_n_ana_[15] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3324 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3325 net44 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3328 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3329 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3330 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3332 a_19154_7663# w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3333 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3334 a_20626_4943# clknet_0_w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3336 a_18786_12559# clknet_0_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3337 net29 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3338 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3340 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3341 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3343 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3345 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3347 net26 w_dly_sig2_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3348 a_14633_9295# a_13643_9295# a_14507_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3349 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3352 r_dly_store_ring[8] a_18171_8475# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3354 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3356 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3358 VGND net63 a_19705_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3359 dbg_dly_sig[6] a_13696_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3360 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3361 clknet_2_2__leaf_w_dly_stop a_14278_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3364 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3365 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3368 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3369 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3370 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3371 a_23570_8751# clknet_0_w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3372 a_22097_6031# net15 w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3373 a_9585_10927# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3375 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3376 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3377 a_13054_11445# net81 a_13269_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3381 o_result_ring[2] a_16403_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3382 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3383 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3386 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3387 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3388 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3389 dbg_ring_ctr[0] a_13955_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3390 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3391 VPWR a_19255_7119# o_result_ring[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3392 VPWR a_15427_10927# a_15595_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3393 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3394 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[5] net37 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3395 VGND clknet_2_0__leaf_w_dly_stop net6 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3396 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3397 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3400 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3401 dbg_dly_sig[12] a_23356_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3402 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3403 VGND clknet_0_i_stop a_21362_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3404 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3405 a_13825_12131# a_13551_12375# a_13743_12131# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3406 VGND a_24462_8319# a_24420_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3408 VGND a_23989_11471# dbg_ring_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3409 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3413 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3415 VGND clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3419 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3420 o_result_ctr[0] a_18795_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3422 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3423 w_dly_sig1_n_ana_[4] net27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3424 dbg_dly_sig[9] a_18112_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3427 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3430 net71 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3431 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3438 net79 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3440 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3441 a_11863_9011# r_dly_store_ring[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X3442 a_9849_8181# clknet_0_w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3444 a_20337_7093# w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3445 VGND w_dly_sig1_n_ana_[2] a_14278_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3446 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3447 VPWR a_14967_4399# a_15135_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3448 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3449 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3451 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3453 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3454 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3455 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3456 net23 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3460 net67 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3461 VPWR w_dly_sig1_n_ana_[6] a_16486_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3462 a_20069_6575# net53 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3464 VGND w_dly_sig2_n_ana_[11] net58 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3465 net73 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3466 VPWR a_16403_8751# o_result_ring[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3467 dbg_dly_sig[1] a_14011_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3468 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3469 VGND a_12035_10535# r_dly_store_ring[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3470 net36 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3473 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3475 VPWR a_13693_18762# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3478 net77 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3479 VPWR a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3481 VPWR w_strt_pulse_n dbg_start_pulse VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X3482 VGND a_14675_9563# a_14633_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3483 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3484 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3486 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3487 VPWR clknet_2_2__leaf_w_dly_stop net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3488 VGND net40 a_16679_5495# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3490 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3491 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3492 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[6] net40 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3497 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3499 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3503 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3505 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3506 VPWR r_dly_store_ring[7] a_18703_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3508 a_21364_12375# net78 a_21281_12117# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3509 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3510 a_15185_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3511 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3512 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3513 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3514 VGND clknet_0_w_dly_sig1_n_ana_[8] a_18773_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3518 a_19215_13335# a_19506_13225# a_19457_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3519 w_dly_stop a_9871_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3520 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3521 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3522 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3523 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3525 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net81 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3526 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3528 a_16198_6397# a_15759_6031# a_16113_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3531 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3532 VPWR a_14462_8181# a_14391_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3534 _01_ _06_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3536 o_result_ring[0] a_16127_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3539 VPWR w_dly_sig1_n_ana_[15] a_16565_11445# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3540 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3541 VPWR a_11863_9011# o_result_ring[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3542 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3543 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3545 a_24209_8207# net61 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3546 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3547 a_16707_6397# a_15925_6031# a_16623_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3548 net24 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3550 VPWR w_dly_sig1_n_ana_[13] a_19430_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3551 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3554 dbg_ring_ctr[0] a_13955_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3555 VGND r_ring_ctr[1] a_18703_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3557 net30 w_dly_sig2_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3558 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3559 w_dly_sig1_n_ana_[3] net23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3560 VPWR net4 w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3561 VGND a_19255_7119# o_result_ring[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3562 VPWR a_19047_13335# r_ring_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3563 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3565 VGND clknet_0_w_dly_sig1_n_ana_[1] a_12425_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3566 VPWR net9 w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3569 o_result_ring[2] a_16403_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3572 a_12438_6575# w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3573 VPWR net54 a_9585_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3574 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3575 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3577 VPWR a_13955_10357# dbg_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3579 VGND a_12622_6005# a_12551_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3581 VGND clknet_0_w_dly_sig1_n_ana_[11] a_21270_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3582 VGND a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3584 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3585 VPWR clknet_0_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3586 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3587 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3588 a_16324_6031# a_15925_6031# a_16198_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3589 a_18786_12559# clknet_0_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3590 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3591 VGND a_13693_18762# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3592 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3593 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3595 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3598 VPWR clknet_0_w_dly_stop a_11045_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3599 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3600 a_18773_10357# clknet_0_w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3601 _85_.X a_18296_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3605 VGND clknet_0_w_dly_sig1_n_ana_[5] a_14081_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3607 VPWR w_dly_strt_ana_[3] a_13825_12131# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3608 VGND clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3609 VPWR a_22383_9295# o_result_ring[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3610 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3611 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3612 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3616 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3617 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3618 o_result_ring[7] a_18703_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3619 net17 clknet_2_3__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3622 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3623 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3624 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3626 a_12373_6397# a_12035_6183# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3628 w_dly_sig1_n_ana_[9] net2 a_18605_4719# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3630 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3631 VGND clknet_0_w_dly_sig1_n_ana_[2] a_11689_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3633 a_17118_13103# a_16679_13109# a_17033_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3634 clknet_0_w_dly_stop a_14278_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3635 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3637 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3638 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3642 net21 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3643 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3644 dbg_dly_sig[11] a_19584_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3646 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3648 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3649 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3652 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3655 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3658 a_20897_10383# net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3659 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3660 net6 clknet_2_0__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3661 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3662 a_11045_10901# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3663 VGND a_15427_10927# a_15595_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3664 VGND w_dly_sig1_n_ana_[14] a_18773_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3665 net7 clknet_2_2__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3667 a_13713_6005# clknet_0_w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3668 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3669 VPWR clknet_2_3__leaf_w_dly_stop net13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3670 a_16854_10383# clknet_0_w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3671 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3672 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[5] net35 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3674 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3676 VGND a_16366_6143# a_16324_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3680 VGND clknet_1_0__leaf_i_stop a_14563_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3682 _06_ net79 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3683 VGND clknet_0_w_dly_sig1_n_ana_[14] a_19430_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3684 a_16210_6575# clknet_0_w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3685 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3686 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3687 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3688 _05_ a_15116_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X3689 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3690 a_12131_6005# a_12415_6005# a_12350_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3691 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3692 a_19154_7663# w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3693 w_dly_sig2_n_ana_[12] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3694 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3695 net66 w_dly_sig2_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3697 a_14637_4399# a_14103_4405# a_14542_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3699 a_20709_10383# a_20543_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3700 VGND a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3701 VGND clknet_2_3__leaf_w_dly_stop net12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3702 a_19881_6581# a_19715_6581# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3704 VPWR clknet_0_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3707 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3709 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3710 net19 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3712 a_20154_6575# a_19715_6581# a_20069_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3713 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3714 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3715 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3716 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3718 a_17627_13103# a_16845_13109# a_17543_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3719 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3720 a_22995_9269# r_dly_store_ring[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X3721 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3722 VPWR w_dly_sig1_n_ana_[7] a_17314_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3725 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3729 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3731 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3732 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3735 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3736 a_21436_12375# _07_ a_21364_12375# VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3737 VPWR r_dly_store_ctr[0] a_18795_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3738 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3739 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3742 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3743 VGND a_11045_10901# clknet_2_1__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3744 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3745 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3746 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3747 VPWR a_19949_13812# _02_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3749 VPWR w_dly_sig1_n_ana_[8] a_19154_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3750 w_dly_sig1_n_ana_[5] net6 a_11337_6895# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3751 net58 w_dly_sig2_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3752 w_dly_strt_ana_[2] a_11711_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3753 VPWR clknet_0_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3755 VGND clknet_0_w_dly_sig1_n_ana_[9] a_20626_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3756 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net76 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3757 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3760 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3762 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3763 a_12415_10357# clknet_1_0__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3764 VGND a_24283_9269# a_24290_9569# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3767 VPWR a_14507_9661# a_14675_9563# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3768 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3769 a_12551_6031# a_12415_6005# a_12131_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3770 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3771 VGND net24 a_13643_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3772 VPWR w_strt_pulse_n dbg_start_pulse VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3773 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3774 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3775 dbg_ring_ctr[1] a_18929_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3778 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3779 a_20280_6953# a_19881_6581# a_20154_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3781 _07_ a_18506_13423# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X3782 a_18773_9269# w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3784 net45 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3785 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3788 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3789 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3790 a_18321_6575# net49 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3791 VGND a_22622_10495# a_22580_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3792 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3793 VPWR i_stop a_17025_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3795 VGND a_18929_13647# dbg_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3797 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3798 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3799 o_result_ring[7] a_18703_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3802 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3803 a_15014_10383# clknet_0_w_dly_sig1_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3804 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3806 a_21491_10749# a_20709_10383# a_21407_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3808 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3809 net53 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3811 a_9585_9839# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3812 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[10] net57 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3814 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3815 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3817 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3818 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3820 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3821 a_16113_6031# net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3822 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3823 dbg_dly_sig[1] a_14011_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3827 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3829 VPWR r_dly_store_ctr[2] a_23119_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3831 a_15925_6031# a_15759_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3833 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3834 a_17305_9295# a_17139_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3836 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[15] net78 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3838 VPWR a_20303_12015# a_20471_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3840 a_18003_9661# a_17139_9295# a_17746_9407# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3841 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3842 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3843 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3844 VGND a_20303_12015# a_20471_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3845 w_dly_sig2_ana_[1] w_dly_sig2_n_ana_[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3846 VPWR a_13955_10357# dbg_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3847 a_12415_6005# clknet_1_0__leaf_i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3849 a_15938_11471# r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.185 ps=1.87 w=0.65 l=0.15
X3850 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3851 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3852 net10 clknet_2_0__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3854 a_14269_4405# a_14103_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3855 VPWR a_15595_10901# a_15511_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3856 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3857 r_ring_ctr[2] a_19047_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3861 net11 clknet_2_3__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3862 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3863 net49 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3865 net52 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3867 o_result_ctr[1] a_21831_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3868 VPWR a_23047_10651# a_22963_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3870 VGND a_14507_9661# a_14675_9563# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3871 VGND clknet_0_w_dly_sig1_n_ana_[3] a_9849_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3872 net32 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3873 VPWR w_dly_sig1_n_ana_[11] a_20337_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3874 net20 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3875 a_14278_8751# w_dly_sig1_n_ana_[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3876 VPWR w_dly_sig1_n_ana_[10] a_21362_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3877 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3878 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3882 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3886 VGND a_17714_12812# r_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X3888 a_20663_6575# a_19881_6581# a_20579_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3891 a_18589_9813# clknet_0_w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3893 r_ring_ctr[0] a_14350_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3894 a_20303_12015# a_19439_12021# a_20046_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3895 VPWR net74 w_dly_sig2_n_ana_[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3896 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3897 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3899 a_14156_12533# dbg_start_pulse VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3900 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3903 net74 w_dly_sig2_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3904 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3908 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3909 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3910 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3913 net54 w_dly_sig2_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3914 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3915 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3916 a_23570_8751# clknet_0_w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3917 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3918 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3920 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3921 a_21362_9839# clknet_0_w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3922 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[7] net43 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3924 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3925 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3927 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3928 a_17314_7663# w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3929 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3931 net68 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3932 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3936 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3937 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3938 a_15116_13103# a_14931_13103# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0767 ps=0.785 w=0.42 l=0.15
X3939 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3940 VGND r_dly_store_ring[8] a_20635_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3942 a_17682_12015# w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3944 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3945 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3946 VPWR r_ring_ctr[0] a_18966_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3947 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3948 a_23903_9447# a_23999_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3949 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3951 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3952 a_11304_9269# net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3953 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3955 a_17025_8725# i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3956 a_18773_4917# clknet_0_w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3957 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3959 VPWR _04_ a_13551_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3960 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3961 VGND a_11987_7671# dbg_dly_sig[4] VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3963 VPWR a_20046_11989# a_19973_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3964 VGND clknet_0_w_dly_sig1_n_ana_[14] a_19430_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3965 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3967 o_result_ring[5] a_11863_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X3968 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X3969 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3970 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3971 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X3972 dbg_dly_sig[3] a_13643_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3973 r_dly_store_ring[3] a_15595_5211# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3974 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3975 net62 w_dly_sig2_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3976 a_18878_8751# clknet_0_w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X3977 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[8] net48 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3978 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[5] net36 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3980 a_19499_13321# clknet_1_1__leaf_w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3981 VPWR a_16127_9839# o_result_ring[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3982 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3983 VGND clknet_0_w_dly_sig1_n_ana_[9] a_21362_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3984 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3985 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3986 a_24419_9295# a_24283_9269# a_23999_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3987 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3990 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3991 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3993 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3994 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3995 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3997 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3999 a_20626_12559# clknet_0_w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4001 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4003 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4006 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4007 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4009 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4012 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4013 VPWR net26 a_9861_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4014 dbg_dly_sig[1] a_14011_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X4015 a_15374_12015# a_15121_12393# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.179 ps=1.26 w=0.42 l=0.15
X4018 VGND clknet_0_i_stop a_12425_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4019 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4020 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4021 VPWR clknet_0_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4023 a_14646_7119# clknet_0_w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4025 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4027 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4028 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4030 o_result_ring[1] a_13059_11187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X4031 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4032 a_20982_10749# a_20543_10383# a_20897_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4033 r_dly_store_ring[3] a_15595_5211# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4035 VGND a_21281_12117# _09_ VGND sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X4036 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4037 net59 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4038 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4039 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4040 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4041 w_dly_sig1_n_ana_[8] net43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4042 r_dly_store_ctr[2] a_23047_10651# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4046 w_dly_sig2_n_ana_[7] clknet_2_1__leaf_w_dly_stop a_9049_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4047 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4048 o_result_ring[14] a_22383_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4049 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4050 VPWR w_strt_pulse_n dbg_start_pulse VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4051 VPWR a_12415_10357# a_12422_10657# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4052 a_22443_8181# r_dly_store_ring[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4054 VPWR a_18703_7119# o_result_ring[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4057 a_17672_12559# a_16679_12559# a_17543_12925# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X4058 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4060 VPWR w_dly_sig1_n_ana_[5] a_14278_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4061 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4065 a_16486_7119# w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4067 VPWR r_ring_ctr[2] a_23989_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4068 VGND net22 w_dly_sig2_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4069 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4070 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4071 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4072 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4074 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4076 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4077 a_20249_6575# a_19715_6581# a_20154_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4079 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4080 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4082 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4083 VPWR a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4084 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4085 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4086 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4087 a_15002_10927# a_14729_10933# a_14917_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4088 o_result_ring[0] a_16127_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4091 a_15121_12393# a_14988_12233# a_14700_11989# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4092 dbg_ring_ctr[2] a_23989_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4093 VGND a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4094 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4095 VGND w_dly_sig2_n_ana_[2] net22 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4096 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4097 VGND a_13054_11445# _04_ VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4098 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4100 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4101 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4103 a_16916_7637# net72 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4104 VGND a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4106 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4107 a_22454_10749# a_22181_10383# a_22369_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4108 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4112 a_21407_10749# a_20543_10383# a_21150_10495# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4114 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4116 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4117 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4119 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4120 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4122 net16 clknet_2_3__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4123 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4124 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4126 a_21077_10749# a_20543_10383# a_20982_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4127 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4131 a_11241_11721# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4133 VGND net17 a_23119_8759# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X4134 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4138 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[8] net47 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4141 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4142 VGND w_dly_sig1_n_ana_[8] a_19154_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4144 VGND clknet_0_w_dly_sig1_n_ana_[10] a_23570_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4145 VPWR clknet_2_3__leaf_w_dly_stop net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4148 o_result_ctr[2] a_23119_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4149 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4150 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[11] net61 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4151 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4153 net78 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4154 a_19430_10927# w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4155 VGND a_12425_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4156 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4158 VGND a_14350_11989# r_ring_ctr[0] VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4159 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4161 VGND _00_ a_15562_12393# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4162 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4165 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4167 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4168 net39 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4169 net40 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4170 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4172 VGND a_13144_11989# _46_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4173 a_14591_9661# a_13809_9295# a_14507_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4175 VPWR a_13233_12724# w_dly_strt_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4176 VPWR a_12425_8725# clknet_1_0__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4177 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4178 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4179 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4180 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4183 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4184 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4185 a_14278_6575# w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4187 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4189 r_ring_ctr[1] a_17714_12812# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X4190 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4191 a_21150_10495# a_20982_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4193 a_17038_10927# clknet_0_w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4194 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4195 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4198 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4200 VGND a_19949_13812# _02_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4201 VPWR _03_ a_14103_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4202 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4203 w_dly_strt_ana_[2] a_11711_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4207 a_17127_12925# a_16845_12559# a_17033_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X4208 VPWR a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4209 VGND a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4210 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4211 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4213 a_24845_8207# a_23855_8207# a_24719_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4214 a_20337_7093# w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4215 w_dly_sig2_n_ana_[1] clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4216 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4217 VPWR a_13643_7119# dbg_dly_sig[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4218 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4222 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4223 net57 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4225 VPWR net22 a_10137_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4226 a_21362_9839# clknet_0_w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4227 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4229 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4230 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4232 a_18406_6575# a_18133_6581# a_18321_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4233 a_17220_12925# a_16679_12559# a_17127_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0662 ps=0.735 w=0.42 l=0.15
X4234 a_15121_12393# a_14998_12137# a_14700_11989# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0657 ps=0.725 w=0.36 l=0.15
X4235 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4236 VGND w_dly_sig2_n_ana_[14] net70 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4237 a_19605_12021# a_19439_12021# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4239 VGND w_dly_sig1_n_ana_[14] a_18773_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4240 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4242 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4243 VPWR net28 a_11987_7671# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X4244 VGND a_14156_12533# _88_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4246 a_13971_8181# a_14262_8481# a_14213_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4247 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4248 VPWR net42 a_9769_10633# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4249 a_17682_12015# w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4250 _06_ r_ring_ctr[1] a_18966_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.175 ps=1.35 w=1 l=0.15
X4253 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4254 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4257 VGND a_22988_8181# dbg_dly_sig[13] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4260 a_14729_10933# a_14563_10933# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4263 VGND a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4264 VGND a_18703_7119# o_result_ring[7] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4266 VPWR a_10473_9460# w_dly_stop_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4267 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4271 a_18589_9813# clknet_0_w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4272 VGND w_ring_ctr_clk a_17682_12015# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4273 VGND w_dly_sig1_n_ana_[12] a_20613_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4275 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4276 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4278 a_15201_13469# a_14931_13103# a_15116_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4281 VGND a_22742_7093# a_22671_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4284 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4285 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4287 VPWR w_dly_sig2_n_ana_[5] net34 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4288 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4291 VGND r_ring_ctr[2] a_18506_13423# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X4292 clknet_2_1__leaf_w_dly_stop a_11045_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4295 VPWR a_17543_12925# a_17714_12812# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X4296 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4297 VGND a_17682_12015# clknet_0_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4298 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4299 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4301 a_20626_12559# clknet_0_w_ring_ctr_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4302 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4304 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4305 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4308 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4310 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4313 VPWR a_18171_8475# a_18087_8573# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4314 a_24462_8319# a_24294_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4317 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4318 VPWR a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4319 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4321 net46 w_dly_sig2_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4325 a_21362_7663# w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4327 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4329 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4330 VPWR a_14255_8181# a_14262_8481# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4333 o_result_ctr[0] a_18795_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4334 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4335 w_dly_sig2_n_ana_[13] net62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4336 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4338 VGND a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4339 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4341 VGND clknet_0_w_dly_sig1_n_ana_[8] a_18773_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4342 VPWR clknet_0_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4343 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net75 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4345 VPWR net75 a_13551_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X4346 VGND w_dly_sig2_n_ana_[6] net38 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4347 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4348 a_22622_10495# a_22454_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4350 VGND a_22879_10749# a_23047_10651# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4352 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4354 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4356 a_12771_10383# a_12551_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4357 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4358 dbg_dly_sig[4] a_11987_7671# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X4360 a_17286_12695# a_17127_12925# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4362 a_14177_9661# a_13643_9295# a_14082_9661# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4363 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4364 r_dly_store_ring[12] a_24887_8475# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4369 VPWR i_stop a_17025_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4370 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4371 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4373 VGND w_strt_pulse_n dbg_start_pulse VGND sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X4375 VPWR a_18574_6549# a_18501_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4376 VPWR clknet_2_3__leaf_w_dly_stop net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4377 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4378 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4381 a_22251_7093# a_22535_7093# a_22470_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4382 a_13551_11721# dbg_start_pulse w_dly_sig1_n_ana_[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4384 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4385 VGND r_dly_store_ring[9] a_19255_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X4387 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] a_12425_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4388 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4389 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4390 VGND w_dly_sig1_n_ana_[7] a_17314_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4391 net64 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4392 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[1] net19 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4393 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4394 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4395 VPWR clknet_2_2__leaf_w_dly_stop net9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4397 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4398 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4399 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] a_18773_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4400 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4401 a_19793_12015# r_ring_ctr[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4402 VPWR a_13955_10357# dbg_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4403 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4404 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4406 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4407 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4409 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4410 VGND a_24887_8475# a_24845_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4412 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4415 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[13] net68 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4416 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4417 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4420 a_9309_9839# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4421 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[3] net29 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4422 a_18501_6575# a_17967_6581# a_18406_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4424 a_13955_10357# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4425 VGND clknet_0_w_dly_sig1_n_ana_[6] a_18878_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4427 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4429 r_dly_store_ring[7] a_16791_6299# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4430 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4431 r_dly_store_ctr[2] a_23047_10651# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4432 a_19881_6581# a_19715_6581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4433 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4436 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4437 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4438 o_result_ring[4] a_11863_9011# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4441 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4444 VPWR clknet_1_0__leaf_i_stop a_16679_13109# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4445 a_16854_10383# clknet_0_w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4446 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4447 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4448 o_result_ring[6] a_16127_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4450 VPWR a_17543_13103# a_17711_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4451 VPWR clknet_1_0__leaf_i_stop a_17139_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4453 VGND clknet_1_1__leaf_i_stop a_20543_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4454 w_dly_sig1_n_ana_[2] net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4455 VGND a_17543_13103# a_17711_13077# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4457 VGND a_23119_10927# o_result_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4458 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4459 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4460 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4461 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4462 a_12798_6397# a_12551_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4463 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4464 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4465 net12 clknet_2_3__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4466 VGND a_15595_5211# a_15553_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4467 VGND net18 w_dly_sig2_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4469 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4470 VPWR clknet_0_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4471 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4472 VGND clknet_0_w_dly_sig1_n_ana_[3] a_14646_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4473 a_16749_9813# clknet_0_w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4474 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4477 a_11045_10901# clknet_0_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4478 VPWR net5 w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4482 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4483 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4485 a_17314_7663# w_dly_sig1_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4490 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4491 w_dly_sig1_n_ana_[12] net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4493 a_17543_13103# a_16679_13109# a_17286_13077# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4495 clknet_1_0__leaf_i_stop a_12425_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4496 net28 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4497 net56 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4498 net34 w_dly_sig2_n_ana_[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4499 a_20626_8207# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4501 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4503 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4504 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4506 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4508 VPWR r_ring_ctr[0] a_14931_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.109 ps=1.36 w=0.42 l=0.15
X4509 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4511 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4512 VGND w_dly_sig1_n_ana_[6] a_16486_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4513 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4514 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[14] net71 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4515 VGND a_14255_8181# a_14262_8481# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4516 VPWR a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4517 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4518 _88_.X a_14156_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4519 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4520 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4523 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4525 a_10417_7983# net35 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4526 VPWR w_dly_sig2_n_ana_[9] net50 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4527 a_19154_7663# w_dly_sig1_n_ana_[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4528 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4530 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4531 dbg_dly_sig[2] a_11304_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4532 VPWR clknet_0_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4533 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4538 VPWR a_16127_9839# o_result_ring[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4539 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4540 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4542 VPWR a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4543 a_12035_6183# a_12131_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4544 a_13269_11721# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.156 ps=1.36 w=0.42 l=0.15
X4545 a_13809_9295# a_13643_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4546 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4549 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4550 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4553 a_19882_13103# a_19635_13481# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4554 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4555 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4557 VGND a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4558 net41 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4559 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4560 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4562 a_16113_6031# net41 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4563 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4564 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[4] net31 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4567 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4569 a_21108_10383# a_20709_10383# a_20982_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4570 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4572 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4574 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4575 o_result_ring[11] a_21891_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4577 VPWR clknet_0_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4578 VPWR net55 w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4579 dbg_dly_sig[14] a_19860_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4581 VGND a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4582 a_23570_8751# clknet_0_w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4583 a_16366_6143# a_16198_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4586 VGND a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4587 dbg_ring_ctr[1] a_18929_13647# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4588 net25 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4589 o_result_ring[13] a_22995_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X4590 a_22988_8181# net64 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4591 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4593 VPWR a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4594 VGND clknet_2_3__leaf_w_dly_stop net16 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4596 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4599 a_12969_6031# a_12415_6005# a_12622_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X4602 VGND a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4603 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4604 VGND w_dly_sig1_n_ana_[11] a_20337_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4606 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4607 a_12969_6031# a_12422_6305# a_12622_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4614 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4616 a_15192_12292# a_14988_12233# a_15374_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0693 ps=0.75 w=0.42 l=0.15
X4617 VGND clknet_0_w_dly_sig1_n_ana_[15] a_14081_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4618 net69 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4619 o_result_ring[14] a_22383_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4620 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4621 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4622 a_20705_6953# a_19715_6581# a_20579_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4623 VPWR net71 w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4624 a_19706_13380# a_19499_13321# a_19882_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4625 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4626 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4627 a_13059_11187# r_dly_store_ring[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X4628 VGND clknet_0_w_dly_sig1_n_ana_[8] a_18773_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4629 VPWR net30 a_9585_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4630 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4631 net55 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4632 VPWR w_dly_sig1_n_ana_[5] a_14278_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4633 a_11863_6835# r_dly_store_ring[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4635 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4636 a_19635_13481# a_19499_13321# a_19215_13335# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4639 VPWR a_16210_6575# clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X4640 a_16486_7119# w_dly_sig1_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X4642 VPWR clknet_0_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4644 net75 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4645 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4646 dbg_dly_sig[13] a_22988_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4647 a_11337_6895# net31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4648 net38 w_dly_sig2_n_ana_[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4649 a_16749_9813# clknet_0_w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4651 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4652 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4653 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4654 VGND w_strt_pulse_n dbg_start_pulse VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4656 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4657 net18 w_dly_sig2_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4658 VGND clknet_1_0__leaf_i_stop a_17139_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4663 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4664 a_10337_10633# net50 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4665 VGND w_dly_stop a_14278_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4666 VPWR w_dly_stop_ana_[2] a_9871_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4670 VPWR w_dly_sig1_ana_[1] a_14809_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4671 VGND a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4672 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4674 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4675 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4676 VPWR a_13955_10357# dbg_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4677 a_18773_9269# w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4678 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4681 VGND a_19047_13335# r_ring_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4682 VPWR w_dly_sig2_n_ana_[4] net30 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4685 a_19047_13335# a_19215_13335# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4686 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4687 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4689 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4690 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4692 w_dly_sig2_n_ana_[9] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4694 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4695 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4696 r_ring_ctr[1] a_17714_12812# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X4697 VGND w_dly_sig2_n_ana_[10] net54 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4698 VGND a_10473_9460# w_dly_stop_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4701 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4703 dbg_ring_ctr[0] a_13955_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4704 a_24294_8573# a_23855_8207# a_24209_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4705 VPWR a_17682_12015# clknet_0_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4706 net4 clknet_2_2__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4708 VGND clknet_0_w_ring_ctr_clk a_14909_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4710 a_14917_10927# net77 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4711 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4712 VPWR clknet_0_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4713 VGND a_19154_7663# clknet_0_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4714 VGND r_dly_store_ring[6] a_16127_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X4717 VPWR w_strt_pulse_n w_dly_sig2_n_ana_[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4718 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4719 w_dly_sig1_n_ana_[4] net7 a_10141_9071# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4720 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4721 clknet_2_0__leaf_w_dly_stop a_11689_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4723 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4724 a_15002_5309# a_14729_4943# a_14917_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4725 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4726 clknet_0_w_dly_stop a_14278_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4731 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4732 VGND a_19216_6005# dbg_dly_sig[10] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4733 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4734 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[5] net37 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4735 VPWR w_dly_sig1_ana_[1] w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4737 a_15170_10901# a_15002_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4738 VGND clknet_0_w_dly_sig1_n_ana_[2] a_16210_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4740 VPWR a_22879_10749# a_23047_10651# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4741 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4742 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4743 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4744 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4745 VPWR clknet_2_3__leaf_w_dly_stop net17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4746 VPWR clknet_1_1__leaf_i_stop a_17967_6581# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4747 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4748 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[3] net28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4749 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[10] net56 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4750 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4752 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4753 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4754 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4756 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4758 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4759 clknet_0_w_ring_ctr_clk a_17682_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4760 VGND a_23119_10927# o_result_ctr[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4761 net60 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4762 VGND a_11863_9011# o_result_ring[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4765 a_12622_10357# a_12415_10357# a_12798_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4766 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4767 a_13875_8359# a_13971_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4769 clknet_2_3__leaf_w_dly_stop a_20626_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4771 dbg_dly_sig[8] a_17284_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4772 a_12551_10383# a_12415_10357# a_12131_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4773 w_dly_sig2_n_ana_[2] clknet_2_0__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4776 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4778 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4779 a_24420_8207# a_24021_8207# a_24294_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4781 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4784 VGND _02_ a_20053_13481# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4785 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4786 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4787 VPWR a_17314_7663# clknet_0_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4789 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4791 VGND a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4792 net65 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4796 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4797 VGND a_15116_13103# _05_ VGND sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X4798 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4799 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4800 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4801 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4802 a_17244_13481# a_16845_13109# a_17118_13103# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4803 VGND net58 w_dly_sig2_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4804 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4805 VPWR w_dly_sig2_n_ana_[13] net66 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4806 clknet_0_w_ring_ctr_clk a_17682_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4807 VPWR r_dly_store_ring[2] a_16403_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4808 a_19216_6005# net52 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X4809 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[1] net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4810 a_17025_8725# i_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4811 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4813 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4814 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4815 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4817 VPWR a_19860_7093# dbg_dly_sig[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4818 a_18773_8181# clknet_0_w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4820 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4821 VGND w_dly_sig1_n_ana_[12] a_20613_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4823 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X4825 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4826 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4827 net50 w_dly_sig2_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4828 dbg_dly_sig[0] a_11672_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X4829 a_15128_4943# a_14729_4943# a_15002_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4831 a_14250_9407# a_14082_9661# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4836 VGND a_18574_6549# a_18532_6953# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4837 w_dly_sig2_n_ana_[10] net50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4838 VPWR a_14278_7663# clknet_2_2__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4841 VGND clknet_0_w_dly_sig1_n_ana_[5] a_15014_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4842 VGND clknet_2_2__leaf_w_dly_stop net5 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4843 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4847 a_23202_9839# clknet_0_w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4848 VGND a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4850 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4851 clknet_0_i_stop a_17025_8725# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4852 VGND a_15427_5309# a_15595_5211# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4855 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4857 net51 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4858 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4859 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4861 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4862 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4863 VPWR w_dly_sig1_n_ana_[4] a_12438_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4864 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4866 a_19216_6005# net52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4867 a_14646_7119# clknet_0_w_dly_sig1_n_ana_[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4868 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[14] net72 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4869 a_21362_7663# w_dly_sig1_n_ana_[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4871 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4872 VPWR a_11863_9011# o_result_ring[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4873 VGND a_18929_13647# dbg_ring_ctr[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4874 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4875 VPWR a_23989_11471# dbg_ring_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4876 a_23005_10383# a_22015_10383# a_22879_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4877 o_result_ring[12] a_22443_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4879 a_17746_8319# a_17578_8573# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4881 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4883 VPWR clknet_0_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4884 a_17746_8319# a_17578_8573# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4885 VGND clknet_2_3__leaf_w_dly_stop net14 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4886 VPWR a_16127_5487# o_result_ring[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4887 VGND a_17286_12695# a_17224_12559# VGND sky130_fd_pr__nfet_01v8 ad=0.149 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X4889 VGND a_15170_5055# a_15128_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4891 net42 w_dly_sig2_n_ana_[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4892 VGND a_21575_10651# a_21533_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4895 w_dly_sig1_n_ana_[7] net4 a_16581_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4896 a_18574_6549# a_18406_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4897 VGND clknet_0_w_dly_sig1_n_ana_[15] a_14081_11445# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4898 VGND clknet_0_w_dly_sig1_n_ana_[13] a_21362_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4899 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4900 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4903 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4904 VPWR a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4905 VPWR a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4907 VPWR _08_ a_21281_12117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.0744 ps=0.815 w=0.42 l=0.15
X4908 a_15553_11305# a_14563_10933# a_15427_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4909 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4911 w_dly_sig1_n_ana_[15] net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4912 VPWR a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4914 dbg_ring_ctr[2] a_23989_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4918 a_20046_11989# a_19878_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4919 VPWR a_20626_8207# clknet_2_3__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4921 a_23202_7663# clknet_0_w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4922 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4924 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4925 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4926 r_dly_store_ring[15] a_18171_9563# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4927 VGND clknet_2_0__leaf_w_dly_stop net8 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4930 VPWR clknet_0_w_dly_sig1_n_ana_[13] a_16749_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4931 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4933 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4936 r_dly_store_ctr[0] a_17711_13077# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4937 a_12350_6031# a_12035_6183# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4938 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4939 clknet_0_w_dly_sig1_n_ana_[2] a_14278_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4940 r_dly_store_ctr[0] a_17711_13077# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4941 clknet_1_1__leaf_w_ring_ctr_clk a_20626_12559# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4942 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4943 VGND w_dly_sig1_n_ana_[7] a_17314_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4947 a_14542_4399# a_14269_4405# a_14457_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4948 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4949 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[9] net53 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4950 VGND a_16679_5495# dbg_dly_sig[7] VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4951 VGND w_dly_stop a_14278_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4952 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4955 VPWR clknet_0_w_dly_stop a_20626_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4958 a_21891_6835# r_dly_store_ring[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X4959 net31 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4960 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4961 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4964 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4966 r_dly_store_ctr[1] a_20471_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4968 r_dly_store_ctr[1] a_20471_11989# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4969 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4971 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4972 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4974 VPWR w_dly_sig2_n_ana_[0] w_dly_sig2_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4975 VPWR a_23119_8759# _87_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4977 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4979 r_ring_ctr[2] a_19047_13335# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4980 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4982 a_9849_7093# clknet_0_w_dly_sig1_n_ana_[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4984 a_14988_12233# clknet_1_0__leaf_w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4985 VPWR a_18773_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4986 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4987 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4988 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] a_11689_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4989 VGND a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4990 VGND w_dly_sig1_n_ana_[8] a_19154_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4991 VGND a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4992 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4993 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4994 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4996 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4997 VGND a_14909_12533# clknet_1_0__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X4998 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[1] net20 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4999 VGND clknet_0_w_dly_sig1_n_ana_[10] a_23570_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5001 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5003 VGND clknet_0_w_ring_ctr_clk a_14909_12533# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5004 a_16198_6397# a_15925_6031# a_16113_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5005 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5006 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5007 VPWR a_17284_6005# dbg_dly_sig[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5008 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5011 a_23989_11471# r_ring_ctr[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5012 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X5013 VGND a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5016 VPWR a_14350_11989# r_ring_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X5017 VPWR a_15014_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5019 a_20387_12015# a_19605_12021# a_20303_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5020 w_dly_sig2_n_ana_[0] w_strt_pulse_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5022 VGND a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5026 VPWR a_19430_11471# clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5027 a_11689_7093# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5029 clknet_2_0__leaf_w_dly_stop a_11689_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5030 o_result_ring[6] a_16127_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5031 VPWR a_13713_6005# clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5033 VGND w_dly_sig2_n_ana_[15] net74 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5034 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5035 VGND w_dly_sig1_n_ana_[0] w_dly_sig1_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5036 VPWR a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5037 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5039 VPWR a_21891_6835# o_result_ring[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X5040 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5041 VGND i_stop a_17025_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5042 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X5043 r_dly_store_ring[15] a_18171_9563# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5044 net8 clknet_2_0__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5049 VGND a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5050 a_18003_9661# a_17305_9295# a_17746_9407# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5051 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5052 VGND a_11672_7637# dbg_dly_sig[5] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5053 VPWR a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5055 VPWR clknet_1_0__leaf_i_stop a_14563_10933# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5057 w_ring_ctr_clk a_13551_12559# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5060 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5061 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X5062 VPWR net51 w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5065 a_16565_11445# w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5066 VPWR a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5067 VPWR a_18112_6005# dbg_dly_sig[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5068 a_20337_7093# w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5069 a_15851_11721# r_ring_ctr[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5070 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5073 a_12131_10357# a_12422_10657# a_12373_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5074 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5075 VPWR w_dly_sig1_ana_[1] a_14011_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5077 a_20626_8207# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5078 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] a_18773_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5079 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5080 a_14278_6575# w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5081 VPWR a_23356_8181# dbg_dly_sig[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5082 w_dly_sig1_n_ana_[13] net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5084 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5085 VGND w_dly_sig1_n_ana_[6] a_16486_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5090 VGND w_dly_sig2_n_ana_[12] net62 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5091 VPWR a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5092 VPWR a_14710_4373# a_14637_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5095 VPWR a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5096 VPWR a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5098 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5099 w_strt_pulse_n a_14103_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5101 VGND a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5102 VGND w_dly_stop_ana_[2] a_9871_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5103 clknet_1_1__leaf_i_stop a_21362_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5104 a_17033_13103# r_ring_ctr[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5105 VPWR a_11045_10901# clknet_2_1__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5106 VGND w_dly_sig1_n_ana_[10] a_21362_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5107 dbg_delay_stop clknet_2_0__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5108 VGND a_17314_5487# clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5110 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5111 a_18831_6575# a_17967_6581# a_18574_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5112 a_20613_9269# w_dly_sig1_n_ana_[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5113 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5115 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5117 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5118 net33 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5120 VGND net75 w_dly_sig1_n_ana_[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5122 VPWR a_18773_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5123 VGND a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5126 VGND a_11689_7093# clknet_2_0__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5127 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] a_13713_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5130 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5132 a_17314_5487# clknet_0_w_dly_sig1_n_ana_[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5133 VGND r_dly_store_ring[7] a_18703_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X5134 VPWR r_ring_ctr[1] a_18337_13103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5135 VGND clknet_0_w_dly_sig1_n_ana_[5] a_15014_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5136 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5137 VPWR a_16366_6143# a_16293_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5139 VPWR net57 a_23089_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5140 a_19430_11471# clknet_0_w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5141 a_23202_9839# clknet_0_w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X5142 VGND a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5143 VPWR clknet_0_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5144 a_17493_8207# net45 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5147 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5148 a_23570_8751# clknet_0_w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X5150 VGND a_22383_9295# o_result_ring[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5153 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5154 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5155 VPWR w_dly_strt_ana_[1] a_11711_11471# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5156 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[11] net59 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5157 VGND a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5158 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5159 VPWR a_11689_7093# clknet_2_0__leaf_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5160 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[7] net44 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5164 clknet_0_w_dly_sig1_n_ana_[10] a_21362_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5166 a_15511_5309# a_14729_4943# a_15427_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5168 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5170 a_12438_7663# w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5171 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5172 VGND a_11304_9269# dbg_dly_sig[2] VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5174 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[4] net32 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5175 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5177 net72 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5178 VPWR net78 a_21281_12117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5179 dbg_ring_ctr[2] a_23989_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5180 a_12350_10383# a_12035_10535# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5181 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5182 a_17025_8725# i_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5183 a_9589_8207# net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5184 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5185 VPWR a_21362_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5186 VGND clknet_1_1__leaf_i_stop a_19439_12021# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5187 VGND a_14081_11445# clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5188 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5189 a_16293_6397# a_15759_6031# a_16198_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5192 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5195 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5199 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5200 VGND a_20626_8207# clknet_2_3__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5201 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5203 VPWR a_18999_6549# a_18915_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5207 VPWR a_23989_11471# dbg_ring_ctr[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5209 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] a_16749_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5211 VPWR a_16565_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5212 VPWR r_ring_ctr[0] a_13955_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5216 a_19706_13380# a_19506_13225# a_19855_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5217 clknet_0_w_dly_sig1_n_ana_[13] a_19430_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5218 clknet_1_0__leaf_w_ring_ctr_clk a_14909_12533# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5219 clknet_0_w_dly_sig1_n_ana_[7] a_17314_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5222 VGND a_23202_7663# clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5223 dbg_dly_sig[7] a_16679_5495# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X5227 clknet_0_w_dly_sig1_n_ana_[1] a_15382_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5228 a_22155_7271# a_22251_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5229 o_result_ctr[1] a_21831_12015# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5230 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5232 _85_.X a_18296_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5233 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5234 net5 clknet_2_2__leaf_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5236 VPWR a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5237 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] a_15014_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5238 VGND a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5239 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X5240 a_18129_8207# a_17139_8207# a_18003_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5243 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] a_11689_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X5244 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] a_15185_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5246 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5247 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] a_18589_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5249 VPWR clknet_1_0__leaf_i_stop a_9595_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5250 dbg_dly_sig[11] a_19584_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5252 clknet_0_w_dly_sig1_n_ana_[15] a_16565_11445# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5254 w_dly_sig1_n_ana_[14] net11 a_19433_5807# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5256 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] a_18878_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5257 VPWR clknet_0_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5259 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] a_20626_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5260 a_20613_9269# w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5261 VPWR r_dly_store_ring[3] a_16127_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5262 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5263 VPWR a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5264 VPWR a_20613_9269# clknet_0_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5265 VPWR a_21362_8751# clknet_1_1__leaf_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5267 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[7] net43 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5268 net80 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5271 net76 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5272 r_ring_ctr[0] a_14350_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X5273 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5274 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[1] net21 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5275 clknet_0_i_stop a_17025_8725# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5279 VGND clknet_0_w_dly_sig1_n_ana_[2] a_16210_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5281 a_17033_12559# _01_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5282 _87_.X a_23119_8759# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5284 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5285 r_dly_store_ring[6] a_15135_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5286 VGND a_14646_7119# clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5288 _46_.X a_13144_11989# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5289 a_14081_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5290 a_24241_9661# a_23903_9447# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5292 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[2] net23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5295 a_18773_10357# clknet_0_w_dly_sig1_n_ana_[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5296 VGND a_17025_8725# clknet_0_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5298 VGND a_21270_11471# clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5299 o_result_ring[5] a_11863_6835# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5300 VPWR a_19982_6031# clknet_0_w_dly_sig1_n_ana_[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5301 VGND a_14278_6575# clknet_0_w_dly_sig1_n_ana_[5] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5302 VPWR r_ring_ctr[0] _08_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5303 w_dly_sig1_ana_[1] w_dly_sig1_n_ana_[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5304 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5305 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[13] net67 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5308 clknet_0_w_dly_sig1_n_ana_[4] a_12438_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5309 VGND w_dly_sig2_ana_[1] w_dly_sig2_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5310 a_22181_10383# a_22015_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5311 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[15] net77 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5312 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[14] net73 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5313 VGND a_21362_8751# clknet_1_1__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5316 VGND clknet_0_w_dly_sig1_n_ana_[3] a_14646_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5318 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[8] net48 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5319 VGND clknet_1_0__leaf_w_dly_sig1_n_ana_[5] net36 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5320 a_16749_9813# clknet_0_w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5321 VPWR a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5323 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5324 clknet_2_1__leaf_w_dly_stop a_11045_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X5325 VPWR a_9849_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5326 VPWR a_22443_8181# o_result_ring[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X5327 a_20154_6575# a_19881_6581# a_20069_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5328 VPWR a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5333 VPWR r_ring_ctr[0] a_15851_11721# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5334 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] a_19430_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5335 VPWR a_17714_12812# a_17627_12925# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0913 ps=0.855 w=0.42 l=0.15
X5338 a_15170_10901# a_15002_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5340 a_14729_4943# a_14563_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5342 w_dly_sig1_n_ana_[9] net47 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5345 net70 w_dly_sig2_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5346 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] a_9849_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5347 dbg_dly_sig[6] a_13696_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5348 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5349 clknet_0_w_dly_sig1_n_ana_[11] a_20337_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5351 VPWR a_18795_10927# o_result_ctr[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5353 a_15097_5309# a_14563_4943# a_15002_5309# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5355 a_17578_9661# a_17139_9295# a_17493_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5356 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5357 VPWR net24 a_13643_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X5359 VGND a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5361 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] a_23202_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5362 VPWR clknet_0_w_dly_sig1_n_ana_[11] a_23202_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5364 VGND a_9849_7093# clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5365 a_11304_9269# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5370 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] a_17038_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5371 VPWR a_19430_10927# clknet_0_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5372 VGND net28 a_11987_7671# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5373 VGND net80 a_15201_13469# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5374 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] a_14081_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5375 a_14909_12533# clknet_0_w_ring_ctr_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5376 VPWR a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5377 VGND a_20626_4943# clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5378 net81 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5379 a_18966_11721# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X5380 VPWR clknet_0_w_dly_sig1_n_ana_[9] a_21362_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5381 net63 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5382 dbg_dly_sig[10] a_19216_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5383 clknet_0_w_dly_sig1_n_ana_[12] a_20613_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5384 VPWR a_13059_11187# o_result_ring[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X5387 VGND clknet_1_1__leaf_w_dly_sig1_n_ana_[13] net69 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5388 a_18053_4943# net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5390 a_15051_4399# a_14269_4405# a_14967_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5391 VGND a_12425_8725# clknet_1_0__leaf_i_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5392 clknet_2_3__leaf_w_dly_stop a_20626_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5393 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5394 VPWR a_15382_8207# clknet_0_w_dly_sig1_n_ana_[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5396 VPWR a_16749_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5398 a_17543_12925# a_16845_12559# a_17286_12695# VGND sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X5399 w_dly_sig2_n_ana_[5] clknet_2_1__leaf_w_dly_stop VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5400 VPWR a_16486_7119# clknet_0_w_dly_sig1_n_ana_[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5402 w_dly_strt_ana_[3] a_12263_12015# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5403 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5406 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5410 VGND a_20337_7093# clknet_0_w_dly_sig1_n_ana_[11] VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X5411 VGND a_18786_12559# clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5412 VPWR a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5413 VPWR clknet_0_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5414 a_9769_10633# clknet_2_1__leaf_w_dly_stop w_dly_sig2_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5415 clknet_0_w_dly_sig1_n_ana_[14] a_18773_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5417 VPWR a_14081_5461# clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5419 dbg_dly_sig[5] a_11672_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5421 VPWR w_dly_sig2_n_ana_[8] net46 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5422 VGND a_21362_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5423 net73 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5424 clknet_0_w_dly_sig1_n_ana_[9] a_19982_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5425 clknet_0_w_dly_sig1_n_ana_[5] a_14278_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X5426 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] a_14081_11445# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5427 VPWR a_23570_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5429 VPWR a_18773_10357# clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5430 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5431 VPWR w_dly_sig1_n_ana_[4] a_12438_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5434 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] a_16854_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5439 a_17704_9295# a_17305_9295# a_17578_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5440 dbg_ring_ctr[0] a_13955_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5441 VPWR a_18589_9813# clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5442 VPWR a_17025_8725# clknet_0_i_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5443 a_23356_8181# net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5445 o_result_ring[12] a_22443_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5446 VGND a_18171_8475# a_18129_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5447 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5450 clknet_1_1__leaf_i_stop a_21362_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5451 VPWR clknet_0_w_dly_stop a_11689_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5452 VPWR a_16127_5487# o_result_ring[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5453 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] a_16210_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5455 VGND a_14278_9839# clknet_0_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5456 VPWR clknet_0_i_stop a_21362_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5458 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5459 net67 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5460 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[7] net45 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5461 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5463 VGND a_21362_7663# clknet_0_w_dly_sig1_n_ana_[10] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5465 VGND a_12438_7663# clknet_0_w_dly_sig1_n_ana_[3] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5466 VGND clknet_1_1__leaf_i_stop a_17967_6581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5467 a_19878_12015# a_19605_12021# a_19793_12015# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5470 VPWR a_20322_6549# a_20249_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5471 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] a_21362_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5473 VPWR a_20626_12559# clknet_1_1__leaf_w_ring_ctr_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5474 VPWR a_14278_9839# clknet_0_w_dly_stop VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5475 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] a_18773_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5476 a_23202_7663# clknet_0_w_dly_sig1_n_ana_[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5477 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] a_14646_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5478 VGND a_16854_10383# clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5479 a_13696_5461# net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5481 VPWR clknet_1_0__leaf_w_dly_sig1_n_ana_[12] net64 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5482 net52 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5483 VGND clknet_2_2__leaf_w_dly_stop net2 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5484 VGND w_dly_sig1_n_ana_[11] a_20337_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5487 VGND a_18878_8751# clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5489 VPWR a_19584_6005# dbg_dly_sig[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5490 clknet_0_w_dly_sig1_n_ana_[8] a_19154_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5493 a_19430_10927# w_dly_sig1_n_ana_[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5494 VPWR a_23202_9839# clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5495 a_13955_10357# r_ring_ctr[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5496 VGND a_17746_9407# a_17704_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5497 VGND a_14278_7663# clknet_2_2__leaf_w_dly_stop VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5500 VPWR clknet_0_w_dly_stop a_20626_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5502 VGND a_18773_4917# clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5504 a_12622_10357# a_12422_10657# a_12771_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5505 VPWR clknet_1_0__leaf_i_stop a_14103_4405# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5506 VGND a_14710_4373# a_14668_4777# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5507 VGND a_16623_6397# a_16791_6299# VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5508 a_19949_13812# _09_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5509 a_17286_13077# a_17118_13103# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5510 VGND clknet_2_2__leaf_w_dly_stop net7 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5511 clknet_0_w_dly_sig1_n_ana_[6] a_16486_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5512 o_result_ring[5] a_11863_6835# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5515 a_15014_10383# clknet_0_w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5516 a_12425_9813# clknet_0_w_dly_sig1_n_ana_[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5518 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] a_9849_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5520 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] a_17314_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X5521 clknet_0_w_dly_sig1_n_ana_[3] a_12438_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5523 a_21270_11471# clknet_0_w_dly_sig1_n_ana_[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5524 a_18878_8751# clknet_0_w_dly_sig1_n_ana_[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5525 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] a_23570_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5527 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] a_21270_11471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X5530 a_21362_7663# w_dly_sig1_n_ana_[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5531 net29 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5534 VPWR clknet_0_w_dly_sig1_n_ana_[15] a_18786_12559# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5535 VGND a_12438_6575# clknet_0_w_dly_sig1_n_ana_[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5536 a_16845_13109# a_16679_13109# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5537 a_11689_9269# clknet_0_w_dly_sig1_n_ana_[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5539 VPWR a_11689_9269# clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5540 VPWR a_14278_8751# clknet_0_w_dly_sig1_n_ana_[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5541 VPWR a_17038_10927# clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5543 a_20709_10383# a_20543_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5544 a_17578_8573# a_17305_8207# a_17493_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5546 a_11689_7093# clknet_0_w_dly_stop VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5547 VPWR clknet_1_1__leaf_w_dly_sig1_n_ana_[12] net65 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5548 clknet_2_2__leaf_w_dly_stop a_14278_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5551 VPWR clknet_0_w_dly_sig1_n_ana_[7] a_17314_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5555 a_14081_11445# clknet_0_w_dly_sig1_n_ana_[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5556 a_15185_9269# clknet_0_w_dly_sig1_n_ana_[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5557 VGND i_stop a_17025_8725# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5558 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] a_23202_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5559 _01_ r_ring_ctr[0] a_15938_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X5560 w_dly_sig1_n_ana_[14] net67 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5561 a_14081_5461# clknet_0_w_dly_sig1_n_ana_[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5562 VPWR w_dly_sig1_n_ana_[1] a_15382_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5564 VGND w_dly_strt_ana_[1] a_11711_11471# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5565 VGND a_15185_9269# clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5566 o_result_ring[14] a_22383_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5567 VGND a_11689_8181# clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
C0 dbg_dly_sig[7] VGND 2.99f
C1 o_result_ring[6] VGND 3.32f
C2 dbg_dly_sig[6] VGND 2.69f
C3 dbg_dly_sig[11] VGND 3.4f
C4 dbg_dly_sig[10] VGND 4.22f
C5 dbg_dly_sig[9] VGND 2.94f
C6 dbg_dly_sig[8] VGND 3.12f
C7 o_result_ring[11] VGND 5.41f
C8 o_result_ring[10] VGND 5.2f
C9 o_result_ring[5] VGND 3.84f
C10 dbg_dly_sig[14] VGND 7.42f
C11 o_result_ring[9] VGND 3.79f
C12 o_result_ring[7] VGND 4.18f
C13 dbg_dly_sig[1] VGND 5.44f
C14 dbg_dly_sig[3] VGND 4.44f
C15 dbg_dly_sig[15] VGND 5.27f
C16 o_result_ring[3] VGND 3.75f
C17 dbg_dly_sig[4] VGND 3.57f
C18 dbg_dly_sig[5] VGND 3.68f
C19 dbg_dly_sig[12] VGND 4.25f
C20 dbg_dly_sig[13] VGND 4.72f
C21 o_result_ring[12] VGND 5.05f
C22 o_result_ring[8] VGND 4.87f
C23 o_result_ring[2] VGND 4.48f
C24 o_result_ring[4] VGND 4.41f
C25 i_stop VGND 6.06f
C26 o_result_ring[13] VGND 4.83f
C27 o_result_ring[14] VGND 5.65f
C28 dbg_dly_sig[2] VGND 4.4f
C29 dbg_delay_stop VGND 9.73f
C30 o_result_ring[15] VGND 5.59f
C31 o_result_ring[0] VGND 4.55f
C32 dbg_ring_ctr[0] VGND 5.17f
C33 dbg_dly_sig[0] VGND 5.45f
C34 o_result_ctr[2] VGND 4.45f
C35 o_result_ctr[0] VGND 4.52f
C36 o_result_ring[1] VGND 5.68f
C37 dbg_ring_ctr[2] VGND 5.62f
C38 o_result_ctr[1] VGND 4.63f
C39 dbg_start_pulse VGND 6.52f
C40 dbg_ring_ctr[1] VGND 3.21f
C41 i_start VGND 1f
C42 VPWR VGND 2.7p
C43 a_14457_4399# VGND 0.23f $ **FLOATING
C44 a_14967_4399# VGND 0.609f $ **FLOATING
C45 a_15135_4373# VGND 0.817f $ **FLOATING
C46 a_14542_4399# VGND 0.626f $ **FLOATING
C47 a_14710_4373# VGND 0.581f $ **FLOATING
C48 a_14269_4405# VGND 1.43f $ **FLOATING
C49 a_14103_4405# VGND 1.81f $ **FLOATING
C50 a_14917_4943# VGND 0.23f $ **FLOATING
C51 a_20626_4943# VGND 4.03f $ **FLOATING
C52 a_18773_4917# VGND 4.03f $ **FLOATING
C53 net3 VGND 0.729f $ **FLOATING
C54 net43 VGND 0.773f $ **FLOATING
C55 a_15427_5309# VGND 0.609f $ **FLOATING
C56 a_15595_5211# VGND 0.817f $ **FLOATING
C57 a_15002_5309# VGND 0.626f $ **FLOATING
C58 a_15170_5055# VGND 0.581f $ **FLOATING
C59 a_14729_4943# VGND 1.43f $ **FLOATING
C60 a_14563_4943# VGND 1.81f $ **FLOATING
C61 net37 VGND 0.959f $ **FLOATING
C62 net2 VGND 1.77f $ **FLOATING
C63 net47 VGND 1.74f $ **FLOATING
C64 clknet_1_0__leaf_w_dly_sig1_n_ana_[5] VGND 3.34f $ **FLOATING
C65 clknet_1_0__leaf_w_dly_sig1_n_ana_[8] VGND 4.87f $ **FLOATING
C66 net67 VGND 0.625f $ **FLOATING
C67 a_17314_5487# VGND 4.03f $ **FLOATING
C68 a_16679_5495# VGND 0.648f $ **FLOATING
C69 a_16127_5487# VGND 1.2f $ **FLOATING
C70 r_dly_store_ring[6] VGND 1.46f $ **FLOATING
C71 a_14081_5461# VGND 4.03f $ **FLOATING
C72 net36 VGND 0.965f $ **FLOATING
C73 a_13696_5461# VGND 0.648f $ **FLOATING
C74 clknet_1_0__leaf_w_dly_sig1_n_ana_[9] VGND 3.82f $ **FLOATING
C75 a_19982_6031# VGND 4.03f $ **FLOATING
C76 w_dly_sig1_n_ana_[9] VGND 2.33f $ **FLOATING
C77 a_19584_6005# VGND 0.648f $ **FLOATING
C78 net52 VGND 1.93f $ **FLOATING
C79 a_19216_6005# VGND 0.648f $ **FLOATING
C80 net48 VGND 1.07f $ **FLOATING
C81 net39 VGND 1.53f $ **FLOATING
C82 a_18112_6005# VGND 0.648f $ **FLOATING
C83 a_16113_6031# VGND 0.23f $ **FLOATING
C84 a_17284_6005# VGND 0.648f $ **FLOATING
C85 a_16623_6397# VGND 0.609f $ **FLOATING
C86 a_16791_6299# VGND 0.817f $ **FLOATING
C87 a_16198_6397# VGND 0.626f $ **FLOATING
C88 a_16366_6143# VGND 0.581f $ **FLOATING
C89 a_15925_6031# VGND 1.43f $ **FLOATING
C90 net41 VGND 1.26f $ **FLOATING
C91 a_15759_6031# VGND 1.81f $ **FLOATING
C92 net40 VGND 1.33f $ **FLOATING
C93 clknet_1_0__leaf_w_dly_sig1_n_ana_[6] VGND 4.37f $ **FLOATING
C94 a_13713_6005# VGND 4.03f $ **FLOATING
C95 a_12969_6031# VGND 0.23f $ **FLOATING
C96 net33 VGND 1.24f $ **FLOATING
C97 a_12551_6031# VGND 0.581f $ **FLOATING
C98 a_12622_6005# VGND 0.626f $ **FLOATING
C99 a_12415_6005# VGND 1.81f $ **FLOATING
C100 a_12422_6305# VGND 1.43f $ **FLOATING
C101 a_12131_6005# VGND 0.609f $ **FLOATING
C102 a_12035_6183# VGND 0.817f $ **FLOATING
C103 net51 VGND 1.05f $ **FLOATING
C104 a_20069_6575# VGND 0.23f $ **FLOATING
C105 net44 VGND 1.76f $ **FLOATING
C106 a_18321_6575# VGND 0.23f $ **FLOATING
C107 net55 VGND 1.13f $ **FLOATING
C108 net14 VGND 1.74f $ **FLOATING
C109 a_21891_6835# VGND 1.2f $ **FLOATING
C110 a_21279_6575# VGND 1.2f $ **FLOATING
C111 r_dly_store_ring[10] VGND 0.764f $ **FLOATING
C112 a_20579_6575# VGND 0.609f $ **FLOATING
C113 a_20747_6549# VGND 0.817f $ **FLOATING
C114 a_20154_6575# VGND 0.626f $ **FLOATING
C115 a_20322_6549# VGND 0.581f $ **FLOATING
C116 a_19881_6581# VGND 1.43f $ **FLOATING
C117 net53 VGND 1.91f $ **FLOATING
C118 a_19715_6581# VGND 1.81f $ **FLOATING
C119 clknet_1_0__leaf_w_dly_sig1_n_ana_[7] VGND 4.69f $ **FLOATING
C120 a_18831_6575# VGND 0.609f $ **FLOATING
C121 a_18999_6549# VGND 0.817f $ **FLOATING
C122 a_18406_6575# VGND 0.626f $ **FLOATING
C123 a_18574_6549# VGND 0.581f $ **FLOATING
C124 a_18133_6581# VGND 1.43f $ **FLOATING
C125 net49 VGND 1.68f $ **FLOATING
C126 a_17967_6581# VGND 1.81f $ **FLOATING
C127 a_16210_6575# VGND 4.03f $ **FLOATING
C128 a_14278_6575# VGND 4.03f $ **FLOATING
C129 w_dly_sig1_n_ana_[5] VGND 2.45f $ **FLOATING
C130 a_12438_6575# VGND 4.03f $ **FLOATING
C131 r_dly_store_ring[5] VGND 1.18f $ **FLOATING
C132 a_11863_6835# VGND 1.2f $ **FLOATING
C133 net6 VGND 1.93f $ **FLOATING
C134 net31 VGND 0.734f $ **FLOATING
C135 a_23089_7119# VGND 0.23f $ **FLOATING
C136 r_dly_store_ring[11] VGND 0.84f $ **FLOATING
C137 net57 VGND 1f $ **FLOATING
C138 a_22671_7119# VGND 0.581f $ **FLOATING
C139 a_22742_7093# VGND 0.626f $ **FLOATING
C140 a_22535_7093# VGND 1.81f $ **FLOATING
C141 a_22542_7393# VGND 1.43f $ **FLOATING
C142 a_22251_7093# VGND 0.609f $ **FLOATING
C143 a_22155_7271# VGND 0.817f $ **FLOATING
C144 w_dly_sig1_n_ana_[11] VGND 1.55f $ **FLOATING
C145 a_20337_7093# VGND 4.03f $ **FLOATING
C146 a_19860_7093# VGND 0.648f $ **FLOATING
C147 a_19255_7119# VGND 1.2f $ **FLOATING
C148 r_dly_store_ring[9] VGND 1.15f $ **FLOATING
C149 a_18703_7119# VGND 1.2f $ **FLOATING
C150 r_dly_store_ring[7] VGND 1.72f $ **FLOATING
C151 _85_.X VGND 0.226f $ **FLOATING
C152 a_18296_7093# VGND 0.648f $ **FLOATING
C153 a_16486_7119# VGND 4.03f $ **FLOATING
C154 a_14646_7119# VGND 4.03f $ **FLOATING
C155 a_14011_7119# VGND 1.2f $ **FLOATING
C156 a_13643_7119# VGND 0.648f $ **FLOATING
C157 clknet_1_0__leaf_w_dly_sig1_n_ana_[4] VGND 4.72f $ **FLOATING
C158 a_11689_7093# VGND 4.03f $ **FLOATING
C159 a_9849_7093# VGND 4.03f $ **FLOATING
C160 clknet_1_1__leaf_w_dly_sig1_n_ana_[11] VGND 4.73f $ **FLOATING
C161 net4 VGND 3.49f $ **FLOATING
C162 net25 VGND 3.38f $ **FLOATING
C163 w_dly_sig1_n_ana_[6] VGND 3.99f $ **FLOATING
C164 a_23202_7663# VGND 4.03f $ **FLOATING
C165 a_21362_7663# VGND 4.03f $ **FLOATING
C166 w_dly_sig1_n_ana_[10] VGND 2.22f $ **FLOATING
C167 a_19154_7663# VGND 4.03f $ **FLOATING
C168 w_dly_sig1_n_ana_[8] VGND 2.73f $ **FLOATING
C169 a_17314_7663# VGND 4.03f $ **FLOATING
C170 w_dly_sig1_n_ana_[7] VGND 2.56f $ **FLOATING
C171 a_16916_7637# VGND 0.648f $ **FLOATING
C172 a_16127_7663# VGND 1.2f $ **FLOATING
C173 r_dly_store_ring[3] VGND 1.94f $ **FLOATING
C174 a_14278_7663# VGND 4.03f $ **FLOATING
C175 a_12438_7663# VGND 4.03f $ **FLOATING
C176 a_11987_7671# VGND 0.648f $ **FLOATING
C177 net32 VGND 1.96f $ **FLOATING
C178 a_11672_7637# VGND 0.648f $ **FLOATING
C179 clknet_1_1__leaf_w_dly_sig1_n_ana_[2] VGND 5.63f $ **FLOATING
C180 net5 VGND 0.846f $ **FLOATING
C181 clknet_1_1__leaf_w_dly_sig1_n_ana_[3] VGND 5.19f $ **FLOATING
C182 net15 VGND 3.01f $ **FLOATING
C183 net56 VGND 4.04f $ **FLOATING
C184 a_24209_8207# VGND 0.23f $ **FLOATING
C185 a_24719_8573# VGND 0.609f $ **FLOATING
C186 a_24887_8475# VGND 0.817f $ **FLOATING
C187 a_24294_8573# VGND 0.626f $ **FLOATING
C188 a_24462_8319# VGND 0.581f $ **FLOATING
C189 a_24021_8207# VGND 1.43f $ **FLOATING
C190 net61 VGND 3.06f $ **FLOATING
C191 a_23855_8207# VGND 1.81f $ **FLOATING
C192 a_23356_8181# VGND 0.648f $ **FLOATING
C193 clknet_1_0__leaf_w_dly_sig1_n_ana_[10] VGND 6.65f $ **FLOATING
C194 a_17493_8207# VGND 0.23f $ **FLOATING
C195 a_22988_8181# VGND 0.648f $ **FLOATING
C196 r_dly_store_ring[12] VGND 1.73f $ **FLOATING
C197 a_22443_8181# VGND 1.2f $ **FLOATING
C198 a_20626_8207# VGND 4.03f $ **FLOATING
C199 a_18773_8181# VGND 4.03f $ **FLOATING
C200 a_18003_8573# VGND 0.609f $ **FLOATING
C201 a_18171_8475# VGND 0.817f $ **FLOATING
C202 a_17578_8573# VGND 0.626f $ **FLOATING
C203 a_17746_8319# VGND 0.581f $ **FLOATING
C204 a_17305_8207# VGND 1.43f $ **FLOATING
C205 net45 VGND 2.22f $ **FLOATING
C206 a_17139_8207# VGND 1.81f $ **FLOATING
C207 a_15382_8207# VGND 4.03f $ **FLOATING
C208 a_14809_8207# VGND 0.23f $ **FLOATING
C209 w_dly_sig1_n_ana_[3] VGND 2.68f $ **FLOATING
C210 net28 VGND 2.02f $ **FLOATING
C211 a_14391_8207# VGND 0.581f $ **FLOATING
C212 a_14462_8181# VGND 0.626f $ **FLOATING
C213 a_14255_8181# VGND 1.81f $ **FLOATING
C214 a_14262_8481# VGND 1.43f $ **FLOATING
C215 a_13971_8181# VGND 0.609f $ **FLOATING
C216 a_13875_8359# VGND 0.817f $ **FLOATING
C217 a_11689_8181# VGND 4.03f $ **FLOATING
C218 clknet_0_w_dly_sig1_n_ana_[3] VGND 5.7f $ **FLOATING
C219 a_9849_8181# VGND 4.03f $ **FLOATING
C220 net23 VGND 1.41f $ **FLOATING
C221 clknet_1_1__leaf_w_dly_sig1_n_ana_[10] VGND 4.12f $ **FLOATING
C222 _87_.X VGND 0.226f $ **FLOATING
C223 clknet_1_1__leaf_w_dly_sig1_n_ana_[6] VGND 4.63f $ **FLOATING
C224 clknet_0_w_dly_sig1_n_ana_[2] VGND 6.29f $ **FLOATING
C225 net35 VGND 1.32f $ **FLOATING
C226 net8 VGND 1.25f $ **FLOATING
C227 w_dly_sig1_n_ana_[4] VGND 3.21f $ **FLOATING
C228 a_23570_8751# VGND 4.03f $ **FLOATING
C229 clknet_0_w_dly_sig1_n_ana_[10] VGND 5.82f $ **FLOATING
C230 a_23119_8759# VGND 0.648f $ **FLOATING
C231 net17 VGND 3.39f $ **FLOATING
C232 a_21362_8751# VGND 4.03f $ **FLOATING
C233 a_20635_8751# VGND 1.2f $ **FLOATING
C234 r_dly_store_ring[8] VGND 1.8f $ **FLOATING
C235 a_18878_8751# VGND 4.03f $ **FLOATING
C236 clknet_0_w_dly_sig1_n_ana_[6] VGND 6.73f $ **FLOATING
C237 a_17025_8725# VGND 4.03f $ **FLOATING
C238 a_16403_8751# VGND 1.2f $ **FLOATING
C239 a_14278_8751# VGND 4.03f $ **FLOATING
C240 w_dly_sig1_n_ana_[2] VGND 2.47f $ **FLOATING
C241 clknet_0_i_stop VGND 7.01f $ **FLOATING
C242 a_12425_8725# VGND 4.03f $ **FLOATING
C243 a_11863_9011# VGND 1.2f $ **FLOATING
C244 net9 VGND 0.62f $ **FLOATING
C245 clknet_2_2__leaf_w_dly_stop VGND 13.5f $ **FLOATING
C246 net7 VGND 0.62f $ **FLOATING
C247 net27 VGND 1.06f $ **FLOATING
C248 net63 VGND 4.68f $ **FLOATING
C249 net12 VGND 4.66f $ **FLOATING
C250 a_24837_9295# VGND 0.23f $ **FLOATING
C251 net11 VGND 4.32f $ **FLOATING
C252 a_17493_9295# VGND 0.23f $ **FLOATING
C253 net65 VGND 1.12f $ **FLOATING
C254 a_24419_9295# VGND 0.581f $ **FLOATING
C255 a_24490_9269# VGND 0.626f $ **FLOATING
C256 a_24283_9269# VGND 1.81f $ **FLOATING
C257 a_24290_9569# VGND 1.43f $ **FLOATING
C258 a_23999_9269# VGND 0.609f $ **FLOATING
C259 a_23903_9447# VGND 0.817f $ **FLOATING
C260 r_dly_store_ring[13] VGND 1.04f $ **FLOATING
C261 a_22995_9269# VGND 1.2f $ **FLOATING
C262 a_22383_9295# VGND 1.2f $ **FLOATING
C263 w_dly_sig1_n_ana_[12] VGND 2.72f $ **FLOATING
C264 a_20613_9269# VGND 4.03f $ **FLOATING
C265 w_dly_sig1_n_ana_[14] VGND 3.19f $ **FLOATING
C266 a_18773_9269# VGND 4.03f $ **FLOATING
C267 a_18003_9661# VGND 0.609f $ **FLOATING
C268 a_18171_9563# VGND 0.817f $ **FLOATING
C269 a_17578_9661# VGND 0.626f $ **FLOATING
C270 a_17746_9407# VGND 0.581f $ **FLOATING
C271 a_17305_9295# VGND 1.43f $ **FLOATING
C272 net73 VGND 1.51f $ **FLOATING
C273 a_17139_9295# VGND 1.81f $ **FLOATING
C274 r_dly_store_ring[2] VGND 1.44f $ **FLOATING
C275 a_13997_9295# VGND 0.23f $ **FLOATING
C276 a_15185_9269# VGND 4.03f $ **FLOATING
C277 a_14507_9661# VGND 0.609f $ **FLOATING
C278 a_14675_9563# VGND 0.817f $ **FLOATING
C279 a_14082_9661# VGND 0.626f $ **FLOATING
C280 a_14250_9407# VGND 0.581f $ **FLOATING
C281 a_13809_9295# VGND 1.43f $ **FLOATING
C282 net21 VGND 1.25f $ **FLOATING
C283 a_13643_9295# VGND 1.81f $ **FLOATING
C284 clknet_1_1__leaf_w_dly_sig1_n_ana_[4] VGND 3.78f $ **FLOATING
C285 clknet_0_w_dly_sig1_n_ana_[4] VGND 5.97f $ **FLOATING
C286 a_11689_9269# VGND 4.03f $ **FLOATING
C287 net19 VGND 0.928f $ **FLOATING
C288 a_11304_9269# VGND 0.648f $ **FLOATING
C289 w_dly_stop_ana_[1] VGND 1.36f $ **FLOATING
C290 a_10473_9460# VGND 0.524f $ **FLOATING
C291 a_9871_9295# VGND 0.524f $ **FLOATING
C292 w_dly_stop_ana_[2] VGND 1.04f $ **FLOATING
C293 a_9595_9295# VGND 0.524f $ **FLOATING
C294 net60 VGND 2f $ **FLOATING
C295 clknet_1_1__leaf_w_dly_sig1_n_ana_[12] VGND 3.3f $ **FLOATING
C296 clknet_1_1__leaf_w_dly_sig1_n_ana_[9] VGND 3.88f $ **FLOATING
C297 _86_.X VGND 0.226f $ **FLOATING
C298 net20 VGND 1f $ **FLOATING
C299 net24 VGND 2.75f $ **FLOATING
C300 w_dly_sig1_n_ana_[1] VGND 3.92f $ **FLOATING
C301 a_23202_9839# VGND 4.03f $ **FLOATING
C302 a_21362_9839# VGND 4.03f $ **FLOATING
C303 clknet_0_w_dly_sig1_n_ana_[9] VGND 6.23f $ **FLOATING
C304 a_20359_9839# VGND 1.2f $ **FLOATING
C305 r_dly_store_ring[15] VGND 1.81f $ **FLOATING
C306 clknet_0_w_dly_sig1_n_ana_[12] VGND 5.52f $ **FLOATING
C307 a_18589_9813# VGND 4.03f $ **FLOATING
C308 a_16749_9813# VGND 4.03f $ **FLOATING
C309 a_16127_9839# VGND 1.2f $ **FLOATING
C310 a_14278_9839# VGND 4.03f $ **FLOATING
C311 w_dly_stop VGND 3.52f $ **FLOATING
C312 a_12425_9813# VGND 4.03f $ **FLOATING
C313 a_12040_9813# VGND 0.648f $ **FLOATING
C314 clknet_1_0__leaf_w_dly_sig1_n_ana_[1] VGND 3.94f $ **FLOATING
C315 clknet_1_0__leaf_w_dly_sig1_n_ana_[2] VGND 4.44f $ **FLOATING
C316 net10 VGND 0.996f $ **FLOATING
C317 clknet_1_0__leaf_w_dly_sig1_n_ana_[3] VGND 4.13f $ **FLOATING
C318 net59 VGND 1.65f $ **FLOATING
C319 net64 VGND 2.04f $ **FLOATING
C320 a_22369_10383# VGND 0.23f $ **FLOATING
C321 clknet_1_0__leaf_w_dly_sig1_n_ana_[12] VGND 6.47f $ **FLOATING
C322 a_22879_10749# VGND 0.609f $ **FLOATING
C323 a_23047_10651# VGND 0.817f $ **FLOATING
C324 a_22454_10749# VGND 0.626f $ **FLOATING
C325 a_22622_10495# VGND 0.581f $ **FLOATING
C326 a_22181_10383# VGND 1.43f $ **FLOATING
C327 a_22015_10383# VGND 1.81f $ **FLOATING
C328 r_dly_store_ring[14] VGND 1.45f $ **FLOATING
C329 a_20897_10383# VGND 0.23f $ **FLOATING
C330 a_21407_10749# VGND 0.609f $ **FLOATING
C331 a_21575_10651# VGND 0.817f $ **FLOATING
C332 a_20982_10749# VGND 0.626f $ **FLOATING
C333 a_21150_10495# VGND 0.581f $ **FLOATING
C334 a_20709_10383# VGND 1.43f $ **FLOATING
C335 net69 VGND 2.1f $ **FLOATING
C336 a_20543_10383# VGND 1.81f $ **FLOATING
C337 clknet_1_1__leaf_w_dly_sig1_n_ana_[8] VGND 4.86f $ **FLOATING
C338 clknet_1_1__leaf_w_dly_sig1_n_ana_[1] VGND 5.29f $ **FLOATING
C339 clknet_1_1__leaf_w_dly_sig1_n_ana_[5] VGND 5.42f $ **FLOATING
C340 clknet_0_w_dly_sig1_n_ana_[8] VGND 6.12f $ **FLOATING
C341 a_18773_10357# VGND 4.03f $ **FLOATING
C342 a_16854_10383# VGND 4.03f $ **FLOATING
C343 clknet_0_w_dly_sig1_n_ana_[1] VGND 5.99f $ **FLOATING
C344 a_15014_10383# VGND 4.03f $ **FLOATING
C345 clknet_0_w_dly_sig1_n_ana_[5] VGND 6.17f $ **FLOATING
C346 a_13955_10357# VGND 2.1f $ **FLOATING
C347 a_12969_10383# VGND 0.23f $ **FLOATING
C348 r_dly_store_ring[4] VGND 1.46f $ **FLOATING
C349 net29 VGND 2.23f $ **FLOATING
C350 a_12551_10383# VGND 0.581f $ **FLOATING
C351 a_12622_10357# VGND 0.626f $ **FLOATING
C352 a_12415_10357# VGND 1.81f $ **FLOATING
C353 a_12422_10657# VGND 1.43f $ **FLOATING
C354 a_12131_10357# VGND 0.609f $ **FLOATING
C355 a_12035_10535# VGND 0.817f $ **FLOATING
C356 net18 VGND 0.96f $ **FLOATING
C357 net22 VGND 1.13f $ **FLOATING
C358 net26 VGND 1.08f $ **FLOATING
C359 net38 VGND 0.921f $ **FLOATING
C360 a_11672_10357# VGND 0.648f $ **FLOATING
C361 clknet_2_0__leaf_w_dly_stop VGND 10.4f $ **FLOATING
C362 w_dly_sig2_n_ana_[1] VGND 0.847f $ **FLOATING
C363 w_dly_sig2_n_ana_[2] VGND 1.02f $ **FLOATING
C364 w_dly_sig2_n_ana_[3] VGND 1.13f $ **FLOATING
C365 net50 VGND 0.632f $ **FLOATING
C366 w_dly_sig2_n_ana_[9] VGND 1.03f $ **FLOATING
C367 w_dly_sig2_n_ana_[6] VGND 0.972f $ **FLOATING
C368 net13 VGND 2.11f $ **FLOATING
C369 clknet_1_1__leaf_w_dly_sig1_n_ana_[13] VGND 3.22f $ **FLOATING
C370 clknet_1_1__leaf_w_dly_sig1_n_ana_[7] VGND 4.55f $ **FLOATING
C371 r_dly_store_ring[0] VGND 1.15f $ **FLOATING
C372 a_14917_10927# VGND 0.23f $ **FLOATING
C373 net30 VGND 1.46f $ **FLOATING
C374 net42 VGND 1.12f $ **FLOATING
C375 net34 VGND 1.38f $ **FLOATING
C376 clknet_2_3__leaf_w_dly_stop VGND 12.3f $ **FLOATING
C377 a_23119_10927# VGND 1.2f $ **FLOATING
C378 r_dly_store_ctr[2] VGND 0.932f $ **FLOATING
C379 a_21362_10927# VGND 4.03f $ **FLOATING
C380 clknet_0_w_dly_sig1_n_ana_[13] VGND 5.56f $ **FLOATING
C381 a_19430_10927# VGND 4.03f $ **FLOATING
C382 w_dly_sig1_n_ana_[13] VGND 3.47f $ **FLOATING
C383 a_18795_10927# VGND 1.2f $ **FLOATING
C384 a_17038_10927# VGND 4.03f $ **FLOATING
C385 clknet_0_w_dly_sig1_n_ana_[7] VGND 7.14f $ **FLOATING
C386 a_15427_10927# VGND 0.609f $ **FLOATING
C387 a_15595_10901# VGND 0.817f $ **FLOATING
C388 a_15002_10927# VGND 0.626f $ **FLOATING
C389 a_15170_10901# VGND 0.581f $ **FLOATING
C390 a_14729_10933# VGND 1.43f $ **FLOATING
C391 net77 VGND 1.48f $ **FLOATING
C392 a_14563_10933# VGND 1.81f $ **FLOATING
C393 a_14103_10927# VGND 0.698f $ **FLOATING
C394 r_dly_store_ring[1] VGND 1.98f $ **FLOATING
C395 a_13059_11187# VGND 1.2f $ **FLOATING
C396 clknet_0_w_dly_stop VGND 11.7f $ **FLOATING
C397 a_11045_10901# VGND 4.03f $ **FLOATING
C398 w_dly_sig2_n_ana_[4] VGND 1.56f $ **FLOATING
C399 w_dly_sig2_n_ana_[7] VGND 1.91f $ **FLOATING
C400 w_dly_sig2_n_ana_[5] VGND 1.41f $ **FLOATING
C401 a_18703_11471# VGND 0.424f $ **FLOATING
C402 a_12539_11471# VGND 0.279f $ **FLOATING
C403 clknet_1_0__leaf_w_dly_sig1_n_ana_[11] VGND 4.64f $ **FLOATING
C404 clknet_1_1__leaf_w_dly_sig1_n_ana_[14] VGND 4.06f $ **FLOATING
C405 a_18966_11721# VGND 0.171f $ **FLOATING
C406 net72 VGND 2.68f $ **FLOATING
C407 a_15851_11721# VGND 0.436f $ **FLOATING
C408 a_13551_11721# VGND 0.388f $ **FLOATING
C409 net46 VGND 1.5f $ **FLOATING
C410 net54 VGND 0.999f $ **FLOATING
C411 a_23989_11471# VGND 1.33f $ **FLOATING
C412 a_21270_11471# VGND 4.03f $ **FLOATING
C413 clknet_0_w_dly_sig1_n_ana_[11] VGND 6.62f $ **FLOATING
C414 a_19430_11471# VGND 4.03f $ **FLOATING
C415 clknet_0_w_dly_sig1_n_ana_[14] VGND 5.96f $ **FLOATING
C416 clknet_1_0__leaf_w_dly_sig1_n_ana_[14] VGND 5.57f $ **FLOATING
C417 a_16565_11445# VGND 4.03f $ **FLOATING
C418 _06_ VGND 1.86f $ **FLOATING
C419 a_14081_11445# VGND 4.03f $ **FLOATING
C420 net75 VGND 1.71f $ **FLOATING
C421 a_13054_11445# VGND 0.642f $ **FLOATING
C422 w_strt_pulse_n VGND 3.83f $ **FLOATING
C423 net74 VGND 0.965f $ **FLOATING
C424 w_dly_sig2_n_ana_[15] VGND 0.964f $ **FLOATING
C425 a_11711_11471# VGND 0.524f $ **FLOATING
C426 clknet_2_1__leaf_w_dly_stop VGND 8.27f $ **FLOATING
C427 net62 VGND 0.632f $ **FLOATING
C428 w_dly_sig2_n_ana_[12] VGND 1.3f $ **FLOATING
C429 w_dly_sig2_n_ana_[8] VGND 1.53f $ **FLOATING
C430 w_dly_sig2_n_ana_[10] VGND 1.27f $ **FLOATING
C431 a_21831_12015# VGND 1.2f $ **FLOATING
C432 a_21281_12117# VGND 0.759f $ **FLOATING
C433 net68 VGND 3.01f $ **FLOATING
C434 r_dly_store_ctr[1] VGND 1.08f $ **FLOATING
C435 a_19793_12015# VGND 0.23f $ **FLOATING
C436 a_15562_12393# VGND 0.216f $ **FLOATING
C437 _03_ VGND 1.1f $ **FLOATING
C438 clknet_1_0__leaf_w_dly_sig1_n_ana_[13] VGND 7.43f $ **FLOATING
C439 a_20303_12015# VGND 0.609f $ **FLOATING
C440 a_20471_11989# VGND 0.817f $ **FLOATING
C441 a_19878_12015# VGND 0.626f $ **FLOATING
C442 a_20046_11989# VGND 0.581f $ **FLOATING
C443 a_19605_12021# VGND 1.43f $ **FLOATING
C444 a_19439_12021# VGND 1.81f $ **FLOATING
C445 clknet_1_1__leaf_i_stop VGND 15.9f $ **FLOATING
C446 a_17682_12015# VGND 4.03f $ **FLOATING
C447 a_15121_12393# VGND 0.587f $ **FLOATING
C448 a_15192_12292# VGND 0.627f $ **FLOATING
C449 a_14998_12137# VGND 1.39f $ **FLOATING
C450 a_14988_12233# VGND 1.77f $ **FLOATING
C451 a_14700_11989# VGND 0.599f $ **FLOATING
C452 a_14350_11989# VGND 1.41f $ **FLOATING
C453 a_13743_12131# VGND 0.485f $ **FLOATING
C454 a_13551_12375# VGND 0.478f $ **FLOATING
C455 _46_.X VGND 0.226f $ **FLOATING
C456 w_dly_sig1_ana_[1] VGND 5.83f $ **FLOATING
C457 w_dly_sig2_ana_[1] VGND 1.82f $ **FLOATING
C458 w_dly_strt_ana_[3] VGND 1.32f $ **FLOATING
C459 net70 VGND 1.04f $ **FLOATING
C460 net66 VGND 1.03f $ **FLOATING
C461 net58 VGND 1.47f $ **FLOATING
C462 a_13144_11989# VGND 0.648f $ **FLOATING
C463 w_dly_sig1_n_ana_[0] VGND 1.53f $ **FLOATING
C464 w_dly_sig2_n_ana_[0] VGND 1.21f $ **FLOATING
C465 a_12263_12015# VGND 0.524f $ **FLOATING
C466 w_dly_strt_ana_[2] VGND 1.17f $ **FLOATING
C467 w_dly_sig2_n_ana_[14] VGND 1.37f $ **FLOATING
C468 w_dly_sig2_n_ana_[13] VGND 1.28f $ **FLOATING
C469 w_dly_sig2_n_ana_[11] VGND 1.8f $ **FLOATING
C470 a_17033_12559# VGND 0.216f $ **FLOATING
C471 a_20626_12559# VGND 4.03f $ **FLOATING
C472 a_18786_12559# VGND 4.03f $ **FLOATING
C473 clknet_0_w_dly_sig1_n_ana_[15] VGND 5.69f $ **FLOATING
C474 a_17543_12925# VGND 0.599f $ **FLOATING
C475 a_17714_12812# VGND 1.41f $ **FLOATING
C476 a_17127_12925# VGND 0.627f $ **FLOATING
C477 a_17286_12695# VGND 0.587f $ **FLOATING
C478 a_16845_12559# VGND 1.39f $ **FLOATING
C479 _01_ VGND 1.53f $ **FLOATING
C480 a_16679_12559# VGND 1.77f $ **FLOATING
C481 clknet_1_0__leaf_w_ring_ctr_clk VGND 3.95f $ **FLOATING
C482 net76 VGND 2.69f $ **FLOATING
C483 clknet_0_w_ring_ctr_clk VGND 5.86f $ **FLOATING
C484 a_14909_12533# VGND 4.03f $ **FLOATING
C485 _88_.X VGND 0.226f $ **FLOATING
C486 net81 VGND 1.34f $ **FLOATING
C487 w_ring_ctr_clk VGND 3.04f $ **FLOATING
C488 w_dly_strt_ana_[1] VGND 1.69f $ **FLOATING
C489 a_14156_12533# VGND 0.648f $ **FLOATING
C490 a_13551_12559# VGND 0.524f $ **FLOATING
C491 _04_ VGND 1.29f $ **FLOATING
C492 a_13233_12724# VGND 0.524f $ **FLOATING
C493 a_20053_13481# VGND 0.23f $ **FLOATING
C494 a_18337_13103# VGND 0.253f $ **FLOATING
C495 _07_ VGND 2.4f $ **FLOATING
C496 r_dly_store_ctr[0] VGND 1.79f $ **FLOATING
C497 a_17033_13103# VGND 0.23f $ **FLOATING
C498 _00_ VGND 1.14f $ **FLOATING
C499 clknet_1_1__leaf_w_ring_ctr_clk VGND 3.34f $ **FLOATING
C500 a_19635_13481# VGND 0.581f $ **FLOATING
C501 a_19706_13380# VGND 0.626f $ **FLOATING
C502 a_19506_13225# VGND 1.43f $ **FLOATING
C503 a_19499_13321# VGND 1.81f $ **FLOATING
C504 a_19215_13335# VGND 0.609f $ **FLOATING
C505 a_19047_13335# VGND 0.97f $ **FLOATING
C506 a_18506_13423# VGND 0.55f $ **FLOATING
C507 a_17543_13103# VGND 0.609f $ **FLOATING
C508 a_17711_13077# VGND 0.817f $ **FLOATING
C509 a_17118_13103# VGND 0.626f $ **FLOATING
C510 a_17286_13077# VGND 0.581f $ **FLOATING
C511 a_16845_13109# VGND 1.43f $ **FLOATING
C512 a_16679_13109# VGND 1.81f $ **FLOATING
C513 clknet_1_0__leaf_i_stop VGND 17.7f $ **FLOATING
C514 a_15575_13103# VGND 0.524f $ **FLOATING
C515 _05_ VGND 0.715f $ **FLOATING
C516 a_15116_13103# VGND 0.672f $ **FLOATING
C517 a_14931_13103# VGND 0.604f $ **FLOATING
C518 _02_ VGND 1.03f $ **FLOATING
C519 net78 VGND 2.02f $ **FLOATING
C520 _08_ VGND 2.97f $ **FLOATING
C521 w_dly_sig1_n_ana_[15] VGND 2.16f $ **FLOATING
C522 net79 VGND 2.27f $ **FLOATING
C523 net80 VGND 0.996f $ **FLOATING
C524 _09_ VGND 1.96f $ **FLOATING
C525 a_19949_13812# VGND 0.524f $ **FLOATING
C526 a_18929_13647# VGND 1.33f $ **FLOATING
C527 r_ring_ctr[2] VGND 5.68f $ **FLOATING
C528 r_ring_ctr[1] VGND 6.76f $ **FLOATING
C529 r_ring_ctr[0] VGND 8.67f $ **FLOATING
C530 net71 VGND 4.87f $ **FLOATING
C531 net16 VGND 3.49f $ **FLOATING
C532 clknet_1_1__leaf_w_dly_sig1_n_ana_[15] VGND 4.93f $ **FLOATING
C533 clknet_1_0__leaf_w_dly_sig1_n_ana_[15] VGND 7.73f $ **FLOATING
C534 net1 VGND 4.96f $ **FLOATING
C535 a_13693_18762# VGND 0.524f $ **FLOATING
.ends
