* PEX produced on Fri Mar 29 11:56:26 PM CET 2024 using /foss/tools/osic-multitool/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tt_um_hpretl_tt06_tdc_v2.ext - technology: sky130A

.subckt tt_um_hpretl_tt06_tdc_v2 clk ena rst_n ui_in[3] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[6] uo_out[0] uo_out[3] uo_out[5] uo_out[6] uo_out[7] ui_in[0] ui_in[2] uio_out[1]
+ ui_in[4] uio_out[0] uo_out[1] uio_oe[5] uio_out[6] uio_oe[3] uio_out[5] uio_oe[2]
+ uio_out[7] uio_oe[7] uio_out[4] uio_oe[4] uio_out[3] uio_oe[0] uio_oe[1] uio_out[2]
+ uo_out[4] uo_out[2] ui_in[1] VPWR VGND
X0 VPWR a_19751_15279 a_19919_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1 VGND a_14894_19199 a_14852_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2 VPWR _052_ a_26575_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND a_9004_20149 net21 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR tdc1.r_ring_ctr0 a_28529_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_18723_19605 a_18639_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7 VGND net33 a_21463_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8 tdc1.r_dly_store_ring13 a_30591_18267 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR a_19899_18543 net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_29887_18775 a_30178_18665 a_30129_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X15 a_15511_20719 a_14729_20725 a_15427_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 a_25593_20719 net42 tdc1.w_ring_int_norsz1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X17 _026_ _170_ a_26689_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_22917_19637 a_22751_19637 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_24113_10383 a_23947_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VGND a_3851_13621 _002_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_26141_14735 tdc1.r_ring_ctr5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VPWR a_17208_20149 uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 a_7423_13103 a_6725_13109 a_7166_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X25 VGND a_3571_19252 tdc0.w_dly_stop3 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X27 a_28997_16367 net17 tdc1.w_ring_norsz28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 a_2413_16911 a_1223_16911 a_2304_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X30 a_7710_10749 a_6633_10383 a_7548_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X31 a_3946_15935 a_3778_16189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X32 a_11580_11293 _009_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X35 a_24571_10749 _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X36 VGND a_27403_17973 net24 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X37 a_22178_17277 a_21739_16911 a_22093_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X39 a_27135_15797 net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X41 VPWR net29 a_10975_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X42 tdc1.w_ring_buf31 a_26983_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X43 tdc1.r_ring_ctr7 a_25571_12319 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X44 VPWR tdc0.w_dly_stop5 a_7111_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X45 a_17596_20425 _089_ a_17208_20149 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X46 a_14857_17753 _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X47 VGND a_16825_15797 _077_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X48 uo_out[6] a_13344_20693 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X49 a_25502_15556 a_25295_15497 a_25678_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
R0 VPWR tt_um_hpretl_tt06_tdc_v2_85.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X52 a_22067_13335 a_22351_13321 a_22286_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
R1 uio_oe[7] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X53 VGND _060_ a_17181_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X55 VPWR _099_ a_17044_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X57 VPWR a_12375_13915 a_12291_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X59 net16 a_17567_10099 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X60 VPWR tdc0.w_ring_norsz8 a_11435_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X61 VGND _145_ _148_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X62 a_25431_15657 a_25295_15497 a_25011_15511 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X66 VGND a_16991_14191 a_17159_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X69 a_24571_10749 a_23947_10383 a_24463_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X71 a_17961_11471 a_16771_11471 a_17852_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X73 a_24385_18249 _067_ a_24131_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 a_21307_15101 a_20525_14735 a_21223_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 VPWR tdc1.w_ring_int_norsz5 a_19237_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X76 a_16821_20502 tdc0.r_dly_store_ring1 a_16607_20502 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X77 a_21633_12015 tdc1.r_ring_ctr11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X79 a_14799_11445 net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X81 a_29089_18543 net42 tdc1.w_ring_int_norsz14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X82 VGND a_9723_12925 a_9891_12827 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X83 VPWR tdc0.r_ring_ctr11 a_4154_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X84 a_20832_16911 a_20433_16911 a_20706_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X85 a_4111_17277 a_3247_16911 a_3854_17023 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X86 VGND a_30534_16341 a_30492_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X87 a_8178_14165 a_8010_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X88 a_25321_11247 _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X89 a_30250_12015 a_29173_12021 a_30088_12393 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X90 VPWR a_7201_10625 a_7091_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X91 a_22351_13321 net33 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X92 a_13861_17161 _116_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X93 a_11582_11989 a_11414_12015 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X94 a_24294_15101 a_23855_14735 a_24209_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X95 tdc0.w_ring_buf13 a_6927_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X97 a_19951_11159 _184_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X98 tdc1.w_ring_buf21 a_19071_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X100 VGND a_9374_15935 a_9332_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X101 a_9631_16189 a_8767_15823 a_9374_15935 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X102 a_5445_19631 net19 tdc0.w_ring_norsz15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X105 a_10129_17161 tdc0.w_ring_norsz3 a_10045_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X106 tdc0.w_ring_buf10 a_9135_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X107 VGND tdc0.w_ring_norsz29 tdc0.w_ring_norsz13 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X108 a_16367_12559 a_16017_12559 a_16272_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X109 a_20533_19337 net71 tdc1.w_ring_int_norsz24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X110 tdc0.w_ring_int_norsz9 net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X111 a_17853_13647 a_16863_13647 a_17727_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X112 a_10325_18249 tdc0.w_ring_norsz4 a_10241_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X113 a_23891_20719 a_23193_20725 a_23634_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X114 _003_ a_863_13897 a_1113_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X116 a_12805_17161 tdc0.r_dly_store_ring28 a_12723_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X117 a_18114_13077 a_17946_13103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X118 a_14166_20719 _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X121 a_13603_11445 tdc0.r_ring_ctr1 a_14001_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X123 a_27717_11713 a_27499_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X124 a_26721_12381 a_26686_12147 a_26483_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X125 _001_ a_1099_12744 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X126 a_24915_15511 a_25011_15511 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X129 VPWR a_22495_11739 a_22411_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X130 a_26895_17429 _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X132 a_20445_18543 tdc1.w_ring_norsz9 a_20361_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X133 a_4909_19631 net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X134 VPWR tdc0.w_ring_norsz12 a_7479_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X136 VGND a_27346_17687 _123_ VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X138 VGND tdc0.w_ring_norsz14 tdc0.w_ring_norsz30 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X139 a_22178_17277 a_21905_16911 a_22093_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X140 net35 a_23907_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X141 VPWR net20 _045_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X142 VPWR _188_ a_18417_12809 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X143 tdc0.w_ring_int_norsz1 tdc0.w_ring_norsz0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X144 VGND net46 tdc0.w_ring_int_norsz17 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X145 a_16831_9813 tdc1.r_ring_ctr12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X146 VPWR a_13323_11159 _145_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X147 VGND _198_ _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X149 a_25093_13647 a_25049_13889 a_24927_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X150 tdc0.w_ring_buf12 a_7479_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X151 VGND a_8775_10633 _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X152 a_16692_18921 a_16293_18549 a_16566_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X154 a_8565_16911 a_8399_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X155 VGND tdc1.w_ring_buf31 a_27689_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X156 VPWR a_11915_18267 a_11831_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X157 VGND net21 tdc0.w_ring_norsz3 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X158 a_7097_20175 tdc0.w_ring_buf14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X160 a_30272_13647 a_29191_13647 a_29925_13889 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X161 VGND _198_ _049_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X162 VPWR _076_ a_14166_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X164 _191_ a_13551_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X166 a_11582_17023 a_11414_17277 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X167 VGND _079_ a_13161_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X168 a_18877_17161 _083_ a_18731_17063 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X169 a_29173_12021 a_29007_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X170 a_15731_16483 _073_ a_15659_16483 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X171 a_13814_20719 _134_ a_13344_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X172 a_17673_13109 a_17507_13109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X175 a_6917_17161 net58 tdc0.w_ring_int_norsz29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X176 VPWR _076_ a_16821_20502 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X180 a_12864_20719 _128_ a_12762_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.18 ps=1.36 w=1 l=0.15
X182 VGND tdc0.r_ring_ctr15 a_1047_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X183 a_10229_13897 net54 tdc0.w_ring_int_norsz25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X184 VGND net18 tdc1.w_ring_norsz31 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X185 tdc1.r_dly_store_ctr14 a_18539_13077 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X186 VPWR a_15595_11989 a_15511_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X188 a_15519_14013 a_14821_13647 a_15262_13759 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X190 tdc1.r_dly_store_ctr14 a_18539_13077 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X191 VGND a_14032_16911 uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X193 _119_ a_12723_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X194 tdc0.r_dly_store_ring0 a_16607_15003 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X196 a_15904_11445 net30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X197 VGND _185_ a_18249_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X198 a_2743_12711 tdc0.r_ring_ctr8 a_2977_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X199 VPWR net8 a_13643_9845 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X200 a_5993_13647 tdc0.r_ring_ctr10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X203 _175_ a_24591_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X204 tdc1.w_ring_int_norsz27 tdc1.w_ring_norsz26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R2 net64 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X205 VPWR a_11490_18111 a_11417_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X207 VGND a_18723_19605 a_18681_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X208 tdc0.w_ring_norsz25 net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X209 a_21886_18517 a_21718_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X210 _027_ _174_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X211 a_5694_17023 a_5526_17277 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X212 VGND net41 tdc1.w_ring_int_norsz10 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X213 a_23029_14735 _083_ a_22595_14887 VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X214 a_8730_15253 a_8562_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X216 tdc0.w_ring_int_norsz18 tdc0.w_ring_norsz17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X217 VPWR a_9063_13077 a_8979_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X218 VPWR a_9631_20719 a_9799_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X219 a_6998_13103 a_6559_13109 a_6913_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X221 VGND a_27251_13077 a_27182_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X224 tdc1.r_dly_store_ring26 a_25163_16091 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X225 tdc1.r_dly_store_ring22 a_17987_17429 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X226 a_27403_14709 a_27687_14709 a_27622_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X228 VGND a_15715_17674 tdc1.w_ring_buf4 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X229 VGND a_27095_13345 a_27056_13219 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X233 tdc1.r_dly_store_ring22 a_17987_17429 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X234 a_25558_12015 a_24481_12021 a_25396_12393 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X235 a_19609_14191 tdc1.w_ring_buf24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
R3 tdc0.g_ring319.stg01_48.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X236 a_8838_17277 a_8399_16911 a_8753_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X237 VGND net14 tdc1.w_ring_norsz6 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X239 VGND a_25932_12533 net9 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X240 VPWR a_30959_16341 a_30875_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X241 a_16017_12559 a_15851_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X242 a_11057_17455 net21 tdc0.w_ring_norsz2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X243 VGND a_29883_21428 net1 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X244 VPWR a_9799_20693 a_9715_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X245 VGND net7 a_1315_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X248 a_18455_13103 a_17673_13109 a_18371_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 uo_out[7] a_14172_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X250 VPWR a_16607_15003 a_16523_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X251 _069_ a_14623_16627 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X252 VGND net36 a_24131_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X253 VGND a_14123_11989 a_14081_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X254 a_29913_17999 tdc1.w_ring_buf13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X255 VPWR a_2212_14569 a_2387_14495 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X256 a_23063_14013 a_22199_13647 a_22806_13759 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X257 a_21445_18549 a_21279_18549 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X258 _144_ tdc0.r_ring_ctr1 a_13634_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X259 VPWR a_5087_11471 _197_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X261 VGND a_23358_19605 a_23316_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X262 VGND tdc1.w_ring_norsz16 a_25787_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X263 a_19876_10383 a_18961_10383 a_19529_10625 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X264 VGND net27 a_3247_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X265 a_27149_11471 a_26983_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X266 a_14172_20149 _138_ a_14994_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X267 tdc1.r_dly_store_ring21 a_22311_18517 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X268 a_11672_10205 _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X270 a_12448_20719 tdc0.r_dly_store_ring6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.135 ps=1.27 w=1 l=0.15
X271 tdc1.r_dly_store_ctr7 a_24887_15003 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X272 a_30263_12319 a_30088_12393 a_30442_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X273 a_27156_17999 tdc1.r_dly_store_ring13 a_26581_18145 VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X274 a_14821_13647 a_14655_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X275 a_14642_20175 _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X276 tdc1.r_dly_store_ring21 a_22311_18517 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X277 VGND a_6319_15101 a_6487_15003 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X279 a_24681_20425 _084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X280 a_9577_10383 a_9411_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X281 VPWR tdc1.w_ring_int_norsz28 a_29081_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X283 a_30534_14165 a_30366_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X285 VGND net28 a_8767_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X287 VPWR net30 a_15299_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X289 VPWR net16 _063_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X290 VPWR _054_ a_27304_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X291 a_15427_20719 a_14729_20725 a_15170_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X292 a_22898_19199 a_22730_19453 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X294 VGND _198_ _053_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X296 a_7350_20287 a_7182_20541 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X297 a_5257_19087 tdc0.w_ring_buf15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X299 VPWR tdc1.r_ring_ctr3 a_28823_14557 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X300 a_6813_14569 a_5823_14197 a_6687_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X301 a_27403_14709 a_27694_15009 a_27645_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X302 a_19494_15253 a_19326_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X304 a_15904_11445 net30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X305 tdc1.w_dly_stop1 a_15299_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X306 _101_ a_13091_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X307 a_2304_16911 a_1389_16911 a_1957_17153 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X309 a_25225_20719 net64 tdc1.w_ring_int_norsz17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X310 a_12805_18543 net3 a_12723_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X311 a_7001_12559 a_6835_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X312 VPWR a_16182_14847 a_16109_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X313 VGND net36 a_29927_14197 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X314 tdc0.w_ring_int_norsz0 tdc0.w_ring_norsz31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X315 tdc0.w_ring_buf8 a_15483_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X316 VGND net7 a_1131_13109 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X318 VPWR _070_ a_15731_16483 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X319 VGND _089_ a_14642_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X320 net8 a_9503_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X322 VGND ui_in[5] a_25879_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X323 VPWR a_21791_20327 _090_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X324 a_25016_11721 _175_ a_24551_11623 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X325 a_10869_12559 tdc0.r_ring_ctr4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X326 VGND _133_ a_18703_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X328 VPWR a_20051_10357 a_20038_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 a_10593_15823 tdc0.w_ring_buf3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X330 VGND net76 tdc1.w_ring_int_norsz29 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X331 a_16187_19891 _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X332 a_20119_14191 a_19421_14197 a_19862_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X333 a_14729_13103 a_14195_13109 a_14634_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X334 VPWR tdc1.w_ring_norsz0 a_25593_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X335 VPWR a_12851_12925 a_13019_12827 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X337 VGND a_5602_15935 a_5560_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X338 a_5859_16189 a_4995_15823 a_5602_15935 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X341 _121_ a_26747_18863 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X345 a_8838_17277 a_8565_16911 a_8753_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X346 VPWR net28 a_6559_19637 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X347 VGND tdc1.w_dly_stop4 a_16587_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X348 tdc0.r_dly_store_ring1 a_15595_20693 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X349 a_28977_15657 a_28423_15497 a_28630_15556 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X351 a_29969_13647 a_29925_13889 a_29803_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X352 a_10492_10383 a_9411_10383 a_10145_10625 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X353 a_17852_11471 a_16937_11471 a_17505_11713 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X356 VPWR a_7423_19631 a_7591_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X357 a_17213_14985 tdc0.r_dly_store_ring8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X358 VPWR a_28415_21237 net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X359 a_4420_14735 a_3505_14735 a_4073_14977 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X360 VGND a_7423_19631 a_7591_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X361 net28 a_9279_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X362 VGND a_22311_18517 a_22269_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X363 VGND a_25551_17545 a_25381_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X364 a_13161_17775 tdc0.r_dly_store_ctr7 a_12815_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X365 _074_ _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X368 VPWR a_11582_15253 a_11509_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X370 a_19326_15279 a_18887_15285 a_19241_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X372 tdc1.r_dly_store_ctr13 a_19735_11989 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X373 VPWR net37 a_29559_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X374 VPWR tdc0.w_ring_norsz28 a_7571_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X375 VPWR net6 a_24822_19133 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X376 tdc1.w_ring_buf30 a_29743_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X377 a_27806_16911 a_27491_17063 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X379 a_1739_16911 a_1389_16911 a_1644_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X381 a_9723_12925 a_9025_12559 a_9466_12671 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X383 VGND a_24059_20693 a_24017_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X384 a_20249_12559 a_20083_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X385 tdc0.r_dly_store_ctr14 a_4371_16091 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X386 a_30216_17833 a_29817_17461 a_30090_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X387 VGND net6 a_24822_19133 VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X388 VPWR net27 a_6743_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X389 tdc1.r_dly_store_ctr9 a_22495_11739 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X390 a_29803_13647 a_29357_13647 a_29707_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X392 VGND net17 tdc1.w_ring_norsz29 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X394 tdc0.w_ring_int_norsz26 tdc0.w_ring_norsz25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X395 a_11329_16911 tdc0.w_ring_buf18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X396 a_11782_14013 a_11509_13647 a_11697_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X397 a_4130_16341 a_3962_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X398 VPWR a_23542_10901 a_23469_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X400 a_13603_11445 tdc0.r_ring_ctr3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X402 a_6078_14013 a_5805_13647 a_5993_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X403 _065_ a_27259_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X406 VPWR _185_ a_17417_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X407 a_19311_10383 a_18961_10383 a_19216_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X408 _155_ a_5271_12128 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X410 a_20707_12925 a_20083_12559 a_20599_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X411 a_21905_21263 a_21739_21263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X412 VGND a_22898_19199 a_22856_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X413 a_20533_19631 net15 tdc1.w_ring_norsz19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X414 VPWR a_17107_20937 a_17114_20841 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X416 a_13173_14191 tdc0.r_dly_store_ctr11 a_13091_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X417 VGND net26 a_3339_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X419 a_21647_16367 _083_ a_21729_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X420 VPWR a_10287_20938 tdc0.w_ring_buf22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X421 a_4073_10901 a_3855_11305 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X422 a_17861_13103 tdc1.r_ring_ctr14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X423 VPWR a_9839_17715 net39 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X424 VGND tdc0.w_ring_norsz30 a_6651_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X425 VGND a_9063_13077 a_9021_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X426 a_28529_12015 tdc1.r_ring_ctr1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X427 a_20448_15823 tdc1.r_dly_store_ring5 a_20258_16073 VGND sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X428 a_15027_15823 _102_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
X429 VPWR a_12207_14013 a_12375_13915 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X430 VGND a_27342_15797 a_27271_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X431 a_5510_19199 a_5342_19453 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X433 VGND a_19951_11159 _018_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X434 a_14886_9839 a_13809_9845 a_14724_10217 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X436 a_10287_20938 tdc0.w_ring_norsz22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X437 net15 a_19899_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X438 a_2953_12015 tdc0.r_ring_ctr9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X439 a_15427_20719 a_14563_20725 a_15170_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X440 a_14377_9813 a_14159_10217 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X441 a_26689_14511 tdc1.r_ring_ctr4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X443 a_17133_19631 tdc1.w_ring_norsz23 a_17049_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X444 tdc1.w_ring_norsz30 net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X445 uo_out[1] a_17208_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 a_15170_19605 a_15002_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X447 VGND _148_ _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X448 VGND tdc0.w_ring_norsz11 tdc0.w_ring_int_norsz12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X449 a_17903_16599 tdc1.r_dly_store_ring20 a_18049_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X451 VGND _190_ a_13551_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X452 a_9006_17023 a_8838_17277 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X453 a_15097_20719 a_14563_20725 a_15002_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X454 a_26851_19863 a_27135_19849 a_27070_19997 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X455 a_24681_10625 a_24463_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X456 VPWR tdc1.w_ring_buf7 a_17661_21097 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X457 VGND a_15719_21237 net32 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X459 VGND a_24546_20327 _142_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X461 a_21445_12021 a_21279_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X462 VPWR net16 _060_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X463 a_28714_20719 a_28467_21097 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X464 a_2905_12559 _156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X465 a_17208_20149 _091_ a_17596_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X466 VGND _053_ a_25093_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X467 VPWR _198_ _051_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X469 VPWR tdc0.w_ring_norsz19 a_10515_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X470 a_4387_16367 a_3689_16373 a_4130_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X471 VGND a_13344_20693 uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X473 a_22227_12015 a_21445_12021 a_22143_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 a_21902_11837 a_21629_11471 a_21817_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X476 VPWR net28 a_7571_14197 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X477 net17 a_27772_16341 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X478 a_29818_16189 a_29571_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X479 VPWR a_8343_17455 a_8511_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X481 a_30281_16367 tdc1.w_ring_buf28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X484 VPWR a_8435_14191 a_8603_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X485 a_9121_20719 tdc0.w_ring_buf6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X486 a_17804_15279 _084_ a_17638_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X487 VGND net19 _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 a_11237_17999 tdc0.w_ring_buf20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X490 a_6430_14165 a_6262_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X491 a_25011_15511 a_25302_15401 a_25253_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X492 VGND a_8343_17455 a_8511_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X493 VPWR tdc0.w_ring_norsz28 a_6917_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X494 VGND a_1368_17429 net7 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
R4 VPWR tdc1.stg01_79.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X496 a_7189_12559 tdc0.r_ring_ctr7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X497 a_15002_20719 a_14563_20725 a_14917_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X498 a_7013_11305 a_5823_10933 a_6904_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X499 a_11767_10217 a_11251_9845 a_11672_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X502 VPWR a_10145_10625 a_10035_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X505 a_24451_18864 _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X507 VPWR a_20287_14165 a_20203_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X508 VGND a_28078_16885 a_28007_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X509 VGND a_19131_21237 a_19138_21537 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X510 VGND net23 tdc0.w_ring_norsz10 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X513 a_19337_17455 net14 tdc1.w_ring_norsz20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X514 VGND _097_ a_23996_16599 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X515 a_17302_14013 a_16863_13647 a_17217_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X516 a_28621_20425 tdc1.w_ring_norsz31 a_28537_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 a_14075_19747 _136_ a_14003_19747 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X521 VPWR tdc0.w_ring_norsz6 a_8675_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X522 a_22820_10383 a_21905_10383 a_22473_10625 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X523 a_1865_14165 a_1647_14569 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X526 VPWR _112_ a_13861_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X527 a_15002_12015 a_14729_12021 a_14917_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X528 VPWR a_30591_18267 a_30507_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X530 a_6771_14191 a_5989_14197 a_6687_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X531 a_23055_15975 tdc1.r_dly_store_ring12 a_23201_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X532 VGND a_24275_16885 _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X533 a_1831_15823 a_1481_15823 a_1736_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X535 a_16481_14191 tdc0.w_ring_buf8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X536 a_8638_13077 a_8470_13103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X537 a_12333_13647 a_11343_13647 a_12207_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X538 a_13625_12015 a_13091_12021 a_13530_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X539 a_11965_16911 a_10975_16911 a_11839_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X540 a_26581_18145 _121_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X541 a_25111_20327 tdc1.r_dly_store_ring15 a_25285_20203 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X542 VPWR _092_ a_15271_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X543 a_20717_13897 tdc1.r_dly_store_ring24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X544 _093_ a_13551_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X545 a_22160_10383 _017_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X546 a_8343_17455 a_7479_17461 a_8086_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X547 VPWR a_6557_10901 a_6447_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X548 VPWR a_14415_18365 a_14583_18267 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X549 VGND a_17559_11159 _020_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X550 a_13330_13077 a_13162_13103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X551 a_19066_21263 a_18751_21415 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X553 a_8435_14191 a_7571_14197 a_8178_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
R5 uio_out[1] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X554 a_18731_17063 tdc1.r_dly_store_ring30 a_18877_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X555 a_12977_12559 a_11987_12559 a_12851_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X556 a_8470_13103 a_8197_13109 a_8385_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X557 a_25229_16687 _066_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X558 a_28538_20996 a_28331_20937 a_28714_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X559 VGND net21 tdc0.w_ring_norsz5 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X560 a_10110_11471 _037_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X561 a_23381_20719 tdc1.w_ring_buf18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X562 VGND a_15451_20149 _075_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X563 net10 a_26615_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X564 a_26226_15101 a_25787_14735 a_26141_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X565 a_7423_13103 a_6559_13109 a_7166_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X566 VPWR tdc0.w_ring_norsz27 a_7295_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X567 a_14821_13647 a_14655_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X568 tdc0.w_ring_norsz30 tdc0.w_ring_int_norsz30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X569 tdc0.w_ring_norsz0 net19 a_5173_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X570 a_13162_13103 a_12889_13109 a_13077_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X571 VGND net11 a_15483_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X572 a_20131_20340 tdc1.w_ring_norsz2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X574 a_24485_15823 tdc1.w_ring_buf26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X575 _050_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X576 net19 a_4404_19061 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X577 a_28467_21097 a_28331_20937 a_28047_20951 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X579 a_29887_18775 a_30171_18761 a_30106_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X581 a_11763_11445 _146_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X582 VGND a_19402_16341 a_19360_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X584 a_7093_13103 a_6559_13109 a_6998_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X585 a_4595_11231 _040_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X586 _118_ a_12079_16073 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X588 a_3854_17023 a_3686_17277 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X590 VGND tdc0.w_ring_int_norsz28 tdc0.w_ring_norsz28 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X591 a_24363_14423 a_24459_14423 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X592 a_10597_14191 net39 tdc0.w_ring_int_norsz10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X593 VGND _198_ _048_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X595 a_16481_18543 tdc0.w_ring_buf30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X597 VGND net9 a_29007_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X598 a_20817_12801 a_20599_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X600 a_13729_14735 tdc0.r_dly_store_ring16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X601 VGND _065_ _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X602 a_23084_16367 _104_ a_22741_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X603 a_13344_20693 _134_ a_13814_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X604 a_29393_20541 a_29055_20327 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X605 VPWR net33 a_17507_13109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X607 a_7001_12559 a_6835_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X608 a_13809_9845 a_13643_9845 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X609 tdc1.w_ring_norsz27 net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X611 VGND a_24455_17687 _081_ VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X612 tdc0.w_ring_int_norsz13 net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X614 a_9945_15101 a_9411_14735 a_9850_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X615 a_1047_16367 _165_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X616 VGND a_30683_17429 a_30641_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X617 VPWR a_18371_13103 a_18539_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
R6 uio_oe[1] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X618 tdc0.w_ring_norsz16 net19 a_4621_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X621 a_20433_16911 a_20267_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X622 VGND tdc0.w_ring_norsz28 a_7571_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X623 _198_ a_28915_10927 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X625 a_14549_13103 tdc0.w_ring_buf25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X626 tdc1.r_dly_store_ring3 a_22771_17179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X627 VPWR _076_ a_16353_20502 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X628 a_30171_18761 net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X629 VGND net42 tdc1.w_ring_int_norsz13 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X630 a_28173_11471 a_26983_11471 a_28064_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X631 VPWR a_16439_15101 a_16607_15003 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X632 a_9025_10383 tdc0.r_ring_ctr4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X633 a_27772_16341 net18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X634 a_12901_15823 tdc0.r_dly_store_ring21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X635 VPWR tdc1.w_ring_norsz16 a_25225_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X636 VPWR a_19211_19850 tdc1.w_ring_buf6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X637 VPWR tdc1.w_ring_norsz3 a_20349_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X638 _043_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X639 a_7442_12671 a_7274_12925 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X640 VPWR a_4585_17674 tdc0.w_ring_buf0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R7 VPWR tt_um_hpretl_tt06_tdc_v2_94.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X642 VPWR a_13698_11989 a_13625_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X643 VPWR a_9723_12925 a_9891_12827 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X644 a_30791_15279 a_29927_15285 a_30534_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X646 a_3855_11305 a_3339_10933 a_3760_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X647 a_29185_18249 tdc1.w_ring_norsz29 a_29101_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X648 a_11697_19631 tdc0.w_ring_buf23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X650 a_27951_20951 a_28047_20951 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X651 tdc0.w_ring_buf11 a_7847_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X652 a_26111_20938 tdc1.w_ring_norsz16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X653 VPWR net33 a_18703_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
R8 VGND net58 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X654 VGND a_22495_11739 a_22453_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X655 a_30461_15279 a_29927_15285 a_30366_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X656 a_17468_15797 net25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X658 a_2396_15823 a_1315_15823 a_2049_16065 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X659 tdc0.w_ring_buf26 a_9227_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X660 VPWR a_17819_17455 a_17987_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X661 a_21489_10205 _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X664 VGND a_22346_21375 a_22304_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X666 _627_.X a_29467_15287 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X667 VPWR tdc0.r_ring_ctr12 a_2227_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.162 ps=1.33 w=1 l=0.15
X668 VGND a_17819_17455 a_17987_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X669 VPWR tdc0.w_ring_int_norsz14 a_6817_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X671 a_9213_12559 tdc0.r_ring_ctr6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X672 VPWR net16 a_19899_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X673 VGND a_24363_14423 tdc1.r_dly_store_ctr4 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X674 a_24294_15101 a_24021_14735 a_24209_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X675 _034_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X676 tdc1.w_ring_buf31 a_26983_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X677 VPWR a_7166_13077 a_7093_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R9 tdc0.g_ring320.stg01_49.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X678 _012_ _153_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X679 a_11747_15101 a_11049_14735 a_11490_14847 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X681 VPWR a_7350_20287 a_7277_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X682 a_19065_20175 _075_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X683 a_2387_14495 _044_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X684 VGND a_4443_18543 net20 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R10 net46 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X685 VGND _101_ a_14379_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X686 a_20249_12559 a_20083_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X687 VGND net27 a_6743_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X688 a_3963_10927 _040_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X691 tdc1.r_dly_store_ctr12 a_17895_13915 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X692 a_30005_17455 tdc1.w_ring_buf30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X693 VGND a_16991_18543 a_17159_18517 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X694 VPWR a_17852_11471 a_18027_11445 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X695 a_19329_16367 a_18795_16373 a_19234_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X697 a_18681_20009 a_17691_19637 a_18555_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X698 a_17861_12559 tdc1.r_ring_ctr13 a_17773_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X699 a_15929_14735 net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X701 VGND tdc0.w_ring_norsz8 a_11435_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X703 VPWR a_24719_15101 a_24887_15003 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X704 a_6888_10383 _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X705 VGND net29 a_12723_13109 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X707 VPWR _072_ a_12889_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X708 VGND a_22806_13759 a_22764_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X709 a_25221_19605 net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X710 tdc0.r_dly_store_ctr13 a_6027_16091 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X711 VGND _137_ a_13921_19747 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X712 a_20165_19631 net15 tdc1.w_ring_norsz3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X714 a_27709_20425 net42 tdc1.w_ring_int_norsz16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X715 a_24397_19951 _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X716 VPWR _197_ _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X719 VGND _079_ a_19141_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X720 VGND tdc0.w_ring_int_norsz6 tdc0.w_ring_norsz6 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X721 VPWR tdc1.r_ring_ctr0 a_28823_14557 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X722 VGND a_7111_17999 net23 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X725 VPWR tdc1.r_dly_store_ctr1 a_22469_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X726 tdc0.w_ring_norsz12 tdc0.w_ring_norsz28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R11 tdc1.g_ring328.stg01_75.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X729 VPWR net31 a_10883_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X731 VPWR _065_ a_24275_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X732 _115_ a_12723_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X733 VPWR a_9155_15253 a_9071_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X735 VPWR net26 a_6835_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X736 VGND a_19494_15253 a_19452_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X737 VPWR tdc0.r_dly_store_ctr6 a_12993_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X738 VPWR a_2396_15823 a_2571_15797 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X739 tdc1.w_ring_norsz14 net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X740 VGND tdc0.w_ring_norsz3 tdc0.w_ring_int_norsz4 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X741 tdc1.r_dly_store_ctr5 a_26819_15003 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X742 a_3693_15823 tdc0.r_ring_ctr14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X743 _134_ a_18703_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X746 a_9033_19337 net51 tdc0.w_ring_int_norsz22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X748 VPWR a_30534_15253 a_30461_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X749 a_9453_11471 a_9409_11713 a_9287_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X750 a_14729_12021 a_14563_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X751 VGND _197_ _036_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X752 a_15235_19453 a_14453_19087 a_15151_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X753 a_30791_14191 a_29927_14197 a_30534_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X754 a_26920_10927 a_26483_10901 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X755 VGND net28 a_8123_15285 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X757 VPWR a_19862_14165 a_19789_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X758 a_14729_19637 a_14563_19637 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X759 net34 a_23264_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X760 a_14511_21590 a_14329_21590 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X761 a_30461_14191 a_29927_14197 a_30366_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X762 net31 a_16180_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X764 a_7815_11623 _147_ a_7989_11499 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X765 a_24738_15935 a_24570_16189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X766 VGND a_26426_17687 _104_ VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.165 ps=1.82 w=0.65 l=0.15
X767 VGND a_7423_16189 a_7591_16091 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X768 VPWR a_23907_21237 net35 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X770 a_3505_10933 a_3339_10933 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X771 a_6904_11305 a_5989_10933 a_6557_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X772 a_10405_15823 a_10239_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X774 a_24819_17776 _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X777 tdc0.w_ring_norsz17 tdc0.w_ring_int_norsz17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X779 a_22527_20327 tdc1.r_dly_store_ring17 a_22653_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X780 VGND a_12467_19355 a_12425_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X782 a_2977_12559 tdc0.r_ring_ctr9 a_2905_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X783 a_1551_15253 _162_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X784 a_16140_14735 a_15741_14735 a_16014_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X785 VPWR tdc0.w_ring_int_norsz12 a_7737_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X786 a_2374_13103 a_1297_13109 a_2212_13481 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X787 VGND a_15151_19453 a_15319_19355 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X788 VGND _139_ a_24546_20327 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X790 a_17044_17161 _089_ a_16656_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X793 VGND a_10018_14847 a_9976_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X794 VGND tdc0.w_ring_norsz27 a_7295_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X795 a_25381_17429 net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X796 a_28993_14557 tdc1.r_ring_ctr0 a_28905_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X797 a_2049_16065 a_1831_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X798 a_2861_12335 tdc0.r_ring_ctr9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X799 VPWR tdc0.w_dly_stop3 a_3247_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X800 tdc1.w_ring_norsz11 net17 a_27529_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X802 a_18027_11445 a_17852_11471 a_18206_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X803 a_29099_14557 tdc1.r_ring_ctr2 a_28993_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X804 VGND net23 tdc0.w_ring_norsz26 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X805 tdc1.r_ring_ctr1 a_30263_12319 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X806 a_17044_17161 _099_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X808 VGND a_19211_19850 tdc1.w_ring_buf6 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X809 a_30180_12559 a_29265_12559 a_29833_12801 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X810 a_19349_20175 _089_ a_18939_20327 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X812 uo_out[3] a_15196_16073 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X813 a_14399_11169 net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X814 a_20175_16073 _080_ a_20258_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X815 VPWR a_16175_20938 tdc0.w_ring_buf1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X816 VPWR a_5510_19199 a_5437_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X817 a_10145_10625 a_9927_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X819 a_28423_15497 net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X820 tdc0.r_dly_store_ring28 a_9431_17179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X821 VPWR a_6796_17973 net22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X822 _144_ tdc0.r_ring_ctr2 a_13551_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X823 VPWR tdc0.w_ring_norsz21 a_8767_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X824 VGND _115_ a_13461_17571 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X825 VGND net27 a_4903_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X826 _038_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X827 VGND _159_ a_4069_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X828 tdc1.r_ring_ctr10 a_22995_10357 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X829 a_13445_12015 tdc0.r_ring_ctr3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X830 VPWR _102_ a_15282_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X834 VPWR a_1551_15253 _165_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X835 VGND net31 a_14563_20725 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X836 VGND net39 tdc0.w_ring_int_norsz3 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X837 a_19311_10383 a_18795_10383 a_19216_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X838 VGND tdc1.r_ring_ctr15 a_19355_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X840 a_23101_17461 a_22935_17461 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X841 VPWR a_11893_10901 a_11783_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X843 a_25571_13621 a_25396_13647 a_25750_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X844 _184_ _179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X845 a_9103_12247 tdc0.r_ring_ctr4 a_9277_12353 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X847 VGND net27 a_8399_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X849 VGND tdc1.w_ring_int_norsz16 tdc1.w_ring_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X850 a_19421_15279 a_18887_15285 a_19326_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X851 a_18324_15823 tdc1.r_dly_store_ctr12 a_18021_15797 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X852 a_21729_16367 tdc1.r_dly_store_ring19 a_21647_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X853 VPWR net4 a_26754_19133 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X854 a_16658_15279 a_16481_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X855 VGND a_12875_20327 _128_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X856 a_30447_13621 a_30272_13647 a_30626_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X857 a_7550_18543 a_7111_18549 a_7465_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X859 a_7308_20175 a_6909_20175 a_7182_20541 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X860 _138_ a_13921_19747 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X861 a_29615_12559 a_29099_12559 a_29520_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X862 a_21905_16911 a_21739_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X863 VPWR a_30534_14165 a_30461_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X864 a_2387_14495 a_2212_14569 a_2566_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X866 a_21131_17277 a_20267_16911 a_20874_17023 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X867 VPWR _132_ a_13814_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X868 VPWR _170_ a_23947_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X870 VGND net4 a_26754_19133 VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X873 a_10678_16189 a_10239_15823 a_10593_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X874 VPWR net5 a_25221_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X876 VPWR tdc1.w_ring_buf14 a_29989_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X877 a_17049_19631 tdc1.w_ring_int_norsz7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X879 VGND a_12507_10143 tdc0.r_ring_ctr0 VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X881 a_18049_16367 _083_ a_17903_16599 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X882 VPWR tdc1.w_ring_int_norsz17 a_24757_21513 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X883 VGND tdc1.r_ring_ctr5 _174_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X884 VPWR net26 a_5823_14197 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X886 a_9873_18249 tdc0.w_ring_int_norsz4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X887 a_21103_10633 _181_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X888 a_22653_18249 tdc1.w_ring_norsz26 a_22569_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X889 VGND a_26439_14191 _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X890 tdc0.r_ring_ctr0 a_12507_10143 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X891 VPWR a_19919_15253 a_19835_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X895 net32 a_15719_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R12 VGND net70 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X897 a_12333_20009 a_11343_19637 a_12207_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X899 tdc0.w_ring_norsz29 net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X901 a_5791_12533 _160_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.28 ps=1.62 w=0.42 l=0.15
X902 _060_ net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X903 tdc0.r_ring_ctr12 a_2387_14495 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X904 VPWR a_24467_16599 _096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X906 VGND a_25163_16091 a_25121_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X908 a_13603_11445 tdc0.r_ring_ctr0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X911 a_28064_11471 a_27149_11471 a_27717_11713 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X912 a_17567_10099 tdc1.w_dly_stop5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X913 a_27127_16885 tdc1.w_dly_stop5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X914 a_16272_12559 _021_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X915 VPWR tdc0.w_ring_norsz9 a_10597_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X916 a_2705_12335 _157_ a_2623_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X917 a_17128_15823 tdc0.r_dly_store_ring9 a_16825_15797 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X918 a_16968_16745 a_16569_16373 a_16842_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X919 a_6457_19337 net60 tdc0.w_ring_int_norsz31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X920 VPWR a_7815_11623 _150_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X921 VGND net33 a_18887_15285 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X922 VGND a_12391_21629 a_12559_21531 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X923 a_24736_12381 _029_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
R13 tdc1.g_ring319.stg01_66.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X925 VGND tdc0.w_ring_norsz26 a_9227_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X926 a_3855_14735 a_3505_14735 a_3760_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X927 a_17638_15599 _084_ a_17804_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X928 a_13993_16073 tdc0.r_dly_store_ring11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X929 _047_ net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X931 tdc1.r_dly_store_ctr10 a_23967_10901 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X932 net7 a_1368_17429 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X933 VGND net30 a_15299_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X934 tdc0.r_dly_store_ctr10 a_6671_13915 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X935 a_3852_13469 _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X936 a_29435_15797 net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X937 a_30197_12393 a_29007_12021 a_30088_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X940 tdc1.w_dly_stop1 a_15299_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X941 a_7549_13481 a_6559_13109 a_7423_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X942 VGND tdc0.w_ring_norsz24 a_11159_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X943 VGND tdc1.w_ring_norsz5 tdc1.w_ring_int_norsz6 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X944 a_2656_18517 net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X945 VPWR a_19494_15253 a_19421_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X947 a_12723_15823 _083_ a_12901_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X948 a_24459_14423 a_24750_14313 a_24701_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X950 VPWR net34 a_21279_19637 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X951 VPWR a_27003_12257 a_26964_12131 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X952 a_11057_20719 net40 tdc0.w_ring_int_norsz8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X953 a_17468_15797 net25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X954 VPWR tdc1.w_ring_int_norsz1 a_24849_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X957 a_6246_13759 a_6078_14013 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X958 a_17661_21097 a_17107_20937 a_17314_20996 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X959 a_6687_14191 a_5823_14197 a_6430_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X960 a_22093_16911 tdc1.w_ring_buf3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X961 a_9279_21237 net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X962 VPWR a_22143_19631 a_22311_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X963 a_22160_10383 _017_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X964 tdc1.r_dly_store_ring13 a_30591_18267 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X965 a_29791_20175 a_29571_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X966 a_17638_15599 _191_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X967 VGND a_17659_10357 a_17593_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X970 a_13861_17161 _117_ a_14032_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X971 VGND tdc0.w_ring_norsz7 tdc0.w_ring_norsz23 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X972 VGND a_22143_19631 a_22311_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X973 VGND a_24551_11623 _029_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X975 VGND _135_ a_13921_19747 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X976 a_6357_14191 a_5823_14197 a_6262_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X977 a_10678_16189 a_10405_15823 a_10593_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X978 a_22487_13481 a_22358_13225 a_22067_13335 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X979 VGND a_15451_20149 _075_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X980 a_19149_16367 tdc1.w_ring_buf5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X981 a_15543_16885 net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X984 a_28445_19631 net42 tdc1.w_ring_int_norsz15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X985 _087_ a_25221_19605 a_25251_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X986 a_8912_21237 net28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X987 VPWR a_4555_16341 a_4471_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X988 VPWR net20 _046_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X989 VGND tdc0.w_dly_stop3 a_3247_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X991 a_7124_13481 a_6725_13109 a_6998_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X992 a_5468_19087 a_5069_19087 a_5342_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X993 net41 a_26031_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X995 VGND _031_ a_27722_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X997 a_14917_12015 tdc0.r_ring_ctr1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X998 a_16727_20951 a_16823_20951 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X999 VGND a_3854_17023 a_3812_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1001 a_8435_14191 a_7737_14197 a_8178_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1003 a_29519_14165 _169_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1004 a_24939_14013 a_24315_13647 a_24831_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1006 VGND a_15170_19605 a_15128_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1007 VGND tdc0.w_ring_norsz21 a_8767_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1008 a_22937_18249 tdc1.w_ring_int_norsz26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1010 a_29989_15823 a_29435_15797 a_29642_15797 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1011 tdc0.w_ring_norsz28 tdc0.w_ring_norsz12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1012 a_10035_10749 a_9411_10383 a_9927_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1013 VPWR a_24363_14423 tdc1.r_dly_store_ctr4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1014 VGND net27 a_3523_16373 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1016 _113_ a_13583_16705 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1017 VGND a_9839_17715 net39 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1018 tdc1.w_ring_buf30 a_29743_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1020 uo_out[0] a_17804_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1021 a_29571_15823 a_29442_16097 a_29151_15797 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1022 a_3781_17277 a_3247_16911 a_3686_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1023 VPWR a_7442_12671 a_7369_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1024 VPWR tdc0.w_ring_norsz4 a_12355_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1027 tdc1.r_ring_ctr5 a_25571_13621 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1028 _014_ a_2703_10927 a_2953_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1029 a_11789_19087 tdc0.w_ring_buf5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1030 a_16607_20175 a_16353_20502 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1031 _186_ tdc1.r_ring_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1032 VPWR _197_ _036_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1033 tdc1.r_dly_store_ring20 a_17435_16341 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1034 VGND net26 a_6835_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1035 VGND _032_ a_12029_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1037 a_22143_19631 a_21279_19637 a_21886_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1040 a_14001_11471 tdc0.r_ring_ctr0 a_13895_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X1041 a_27871_16885 net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1043 a_4420_14735 a_3339_14735 a_4073_14977 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1044 a_15170_11989 a_15002_12015 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1045 a_29428_12381 _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1046 a_19338_21237 a_19138_21537 a_19487_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1048 a_10402_20541 a_10129_20175 a_10317_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1049 a_3852_12381 _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1050 VGND net35 a_20267_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1051 a_11322_18365 a_10883_17999 a_11237_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1052 VGND _158_ a_1099_12744 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1053 a_24017_21097 a_23027_20725 a_23891_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1054 a_21273_12559 a_20083_12559 a_21164_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1056 a_25623_11247 _180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X1057 tdc0.w_ring_buf3 a_10147_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
R14 VPWR tt_um_hpretl_tt06_tdc_v2_90.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1059 a_27019_18863 tdc1.r_dly_store_ring21 a_26919_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1060 a_3483_14423 _164_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X1062 VGND a_17924_17063 _112_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X1063 VGND _074_ a_27156_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1065 VGND tdc1.w_ring_buf15 a_28885_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1066 a_22741_14985 _083_ a_22595_14887 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X1067 a_3703_15279 _162_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1069 VPWR tdc1.r_ring_ctr11 a_20254_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1070 VPWR a_7591_19605 a_7507_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1071 a_8730_15253 a_8562_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1072 VPWR net26 a_5639_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1073 a_21718_19631 a_21279_19637 a_21633_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1074 a_4241_18543 net44 a_4157_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1075 _005_ _166_ a_1137_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1076 a_25011_15511 a_25295_15497 a_25230_15645 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1078 _173_ a_24347_13441 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1079 a_6447_10927 a_5823_10933 a_6339_11305 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1080 a_1368_17429 tdc0.w_ring_buf0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1081 VGND a_4371_16091 a_4329_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1083 a_30180_12559 a_29099_12559 a_29833_12801 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1084 a_8562_15279 a_8289_15285 a_8477_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1085 a_29725_17999 a_29559_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1086 VPWR _162_ a_2227_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1087 VPWR tdc1.w_ring_int_norsz12 a_29173_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1089 VPWR a_12007_11989 a_11923_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1090 a_23281_19087 a_22291_19087 a_23155_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1091 a_1909_14557 a_1865_14165 a_1743_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1093 a_5271_12128 _149_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1094 a_3947_12393 a_3597_12021 a_3852_12381 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1095 a_20707_12925 _063_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1099 a_14583_21590 tdc1.r_dly_store_ring7 a_14511_21590 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1100 a_17351_16367 a_16569_16373 a_17267_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1102 _042_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1103 _116_ a_13461_17571 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1106 a_6601_11293 a_6557_10901 a_6435_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1107 VPWR net9 a_15851_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1108 VPWR _064_ a_24455_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X1109 a_8912_21237 net28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1110 VPWR _152_ a_7745_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1111 a_6817_18543 tdc0.w_ring_norsz30 a_6733_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R15 VPWR tt_um_hpretl_tt06_tdc_v2_82.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1113 VPWR tdc0.r_dly_store_ring22 a_12875_20327 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1114 VGND tdc0.w_ring_int_norsz31 tdc0.w_ring_norsz31 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1115 tdc0.w_ring_norsz22 net21 a_8853_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1116 VPWR a_26483_11989 tdc1.r_ring_ctr6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1118 _108_ a_22293_15395 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1119 a_19310_11989 a_19142_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1120 tdc1.w_ring_norsz21 net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1121 a_17107_20937 net34 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1124 VPWR _154_ a_5271_12128 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1125 a_29520_12559 _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1126 VPWR a_3854_17023 a_3781_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1127 VPWR a_4420_14735 a_4595_14709 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1128 a_27342_15797 a_27135_15797 a_27518_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1129 a_14583_21263 a_14329_21590 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X1130 a_14003_19747 _137_ a_13921_19747 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1131 a_29427_20693 net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1132 net12 a_5455_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1134 VGND net48 tdc0.w_ring_int_norsz19 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1135 a_19142_12015 a_18869_12021 a_19057_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1136 a_18027_11445 _061_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1139 tdc1.w_ring_norsz8 tdc1.w_ring_int_norsz8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1140 VGND tdc0.w_ring_norsz19 a_10515_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1141 a_22309_13103 a_21971_13335 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1142 a_12341_12559 tdc0.r_ring_ctr0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1143 a_27271_15823 a_27135_15797 a_26851_15797 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X1144 a_23105_19631 tdc1.w_ring_buf23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1145 _169_ a_28823_14557 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1147 a_8987_15279 a_8289_15285 a_8730_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1148 a_27793_18909 _064_ a_27693_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X1149 a_19241_15279 net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1150 tdc0.r_dly_store_ring22 a_10995_20443 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1151 VPWR net6 a_25221_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1152 a_17126_16911 _100_ a_16656_16885 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1153 VPWR net8 a_11251_9845 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1154 VGND a_5859_16189 a_6027_16091 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1157 VPWR a_14802_13077 a_14729_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1158 a_6272_12559 _149_ a_6166_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X1159 net21 a_9004_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1160 VPWR a_16587_10927 tdc1.w_dly_stop5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1161 a_16932_12559 a_15851_12559 a_16585_12801 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1162 a_23855_15279 _071_ a_23937_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1163 VPWR a_13755_13077 a_13671_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1164 tdc0.w_ring_norsz6 tdc0.w_ring_norsz22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1165 net23 a_7111_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X1166 VGND a_30423_18365 a_30591_18267 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1167 _157_ _156_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1168 a_14379_14735 _083_ a_14557_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1169 _055_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1170 VGND net35 a_22751_19637 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1171 a_28599_15797 net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1172 VGND tdc0.w_ring_norsz6 a_8675_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1173 a_22346_17023 a_22178_17277 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1174 a_15899_16911 a_15679_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1176 VGND a_24087_18775 _129_ VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1178 VGND tdc1.w_dly_stop5 a_29467_15287 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1179 a_5441_16911 tdc0.w_ring_buf17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1181 VPWR a_11950_19605 a_11877_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1182 a_8753_16911 tdc0.w_ring_buf28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1183 a_23239_19453 a_22457_19087 a_23155_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1185 VPWR a_26651_15101 a_26819_15003 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1186 a_17857_19637 a_17691_19637 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1187 a_29989_20175 a_29442_20449 a_29642_20149 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X1189 net24 a_27403_17973 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1190 a_18881_14735 tdc1.r_dly_store_ctr14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X1191 _036_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1193 VPWR a_4073_14977 a_3963_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1194 tdc1.r_ring_ctr14 a_17107_12533 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1195 a_23289_17455 tdc1.w_ring_buf25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1198 a_22733_14013 a_22199_13647 a_22638_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1199 a_21934_20221 _089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X1200 a_17691_12559 tdc1.r_ring_ctr14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1201 VGND a_5875_13077 _160_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1202 VGND _050_ a_29969_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1203 a_4512_12393 a_3431_12021 a_4165_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1204 VGND _068_ a_13621_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X1205 a_22982_10749 a_21905_10383 a_22820_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1206 a_30791_14191 a_30093_14197 a_30534_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1208 tdc0.r_dly_store_ring4 a_14583_18267 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1209 a_24743_14409 net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1210 VPWR tdc0.r_ring_ctr8 a_5875_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1211 a_20131_20340 tdc1.w_ring_norsz2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1216 VGND a_5791_12533 _162_ VGND sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.107 ps=0.98 w=0.65 l=0.15
X1217 VGND a_23155_19453 a_23323_19355 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1218 a_4043_12393 a_3597_12021 a_3947_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1219 a_13257_12021 a_13091_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1220 a_17903_17455 a_17121_17461 a_17819_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1221 a_30088_12393 a_29173_12021 a_29741_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1223 _141_ a_23855_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1224 VPWR a_16656_16885 uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1225 _100_ a_16055_19414 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X1226 a_12529_14511 tdc0.r_dly_store_ctr8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1227 VPWR _075_ a_17213_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1228 VPWR tdc0.w_ring_norsz23 a_11067_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1230 VGND a_28630_15556 a_28559_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1231 a_12000_19087 a_11601_19087 a_11874_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1233 VPWR a_14428_17687 _117_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1234 _137_ a_13183_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X1236 a_17727_14013 a_17029_13647 a_17470_13759 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1237 VGND tdc0.r_ring_ctr9 a_2705_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X1238 a_28455_13647 tdc1.r_ring_ctr0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1239 VPWR tdc1.r_dly_store_ring13 a_27012_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X1240 a_27529_16367 tdc1.w_ring_norsz27 a_27445_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1241 VPWR _069_ a_21729_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1242 a_20966_14847 a_20798_15101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1243 VPWR _095_ a_17044_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1244 a_29791_20938 tdc1.w_ring_norsz15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1245 VPWR a_21339_12533 a_21326_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1246 VGND a_14399_11169 a_14360_11043 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1247 a_20981_13647 tdc1.r_dly_store_ring24 a_20635_13897 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
R16 VPWR tdc0.stg01_61.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1248 VPWR a_24887_15003 a_24803_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1251 a_22160_20175 _082_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1252 a_15196_16073 _103_ a_15110_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1253 VGND a_25103_16599 _098_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1254 a_1644_16911 _006_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1255 a_16861_9839 _185_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R17 net53 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1256 VPWR a_28423_15497 a_28430_15401 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1257 a_13633_15599 tdc0.r_dly_store_ring10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1258 net22 a_6796_17973 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1260 a_10045_17161 net21 tdc0.w_ring_norsz19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1263 a_10241_18249 tdc0.w_ring_int_norsz20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1264 tdc1.r_dly_store_ctr2 a_30959_15253 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1265 a_10275_15101 a_9411_14735 a_10018_14847 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1266 a_19421_14197 a_19255_14197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1267 tdc0.r_ring_ctr11 a_4687_13407 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1269 a_14064_10205 _007_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1270 a_3947_12393 a_3431_12021 a_3852_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1271 tdc1.r_dly_store_ctr2 a_30959_15253 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1272 a_15128_21097 a_14729_20725 a_15002_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1273 a_11985_9813 a_11767_10217 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1274 a_21718_12015 a_21279_12021 a_21633_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1275 VGND a_16607_15003 a_16565_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1276 a_1113_13897 tdc0.r_ring_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1277 a_9277_12353 tdc0.r_ring_ctr5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X1278 a_1939_16189 _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1279 VGND _065_ a_26431_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X1280 a_4154_13897 _159_ a_3851_13621 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X1282 VPWR a_22806_13759 a_22733_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1283 _016_ tdc1.r_ring_ctr0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1284 a_9839_17715 net43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1287 a_13799_11471 tdc0.r_ring_ctr3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X1288 _045_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1289 VPWR a_11747_15101 a_11915_15003 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1290 a_1551_15253 tdc0.r_ring_ctr13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X1291 VGND a_4585_17674 tdc0.w_ring_buf0 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1292 tdc0.w_ring_int_norsz17 tdc0.w_ring_norsz16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1293 VGND tdc1.r_ring_ctr12 a_17049_10159 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1294 a_16828_20175 tdc1.r_dly_store_ring1 a_16607_20502 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1295 VPWR a_9756_11471 a_9931_11445 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1296 VPWR a_16585_12801 a_16475_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1297 tdc1.r_ring_ctr11 a_20051_10357 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1299 VPWR tdc1.r_ring_ctr1 a_28977_15657 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1300 a_8289_15285 a_8123_15285 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1301 VGND _167_ _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1302 a_18877_16911 _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X1303 tdc0.w_ring_buf11 a_7847_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1304 a_14166_20719 _131_ a_13344_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1305 a_14300_16911 _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X1307 a_24757_21513 tdc1.w_ring_norsz1 a_24673_21513 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1309 a_22569_18249 tdc1.w_ring_int_norsz10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1311 a_3760_14735 _004_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1313 _102_ a_14379_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
R18 VPWR tt_um_hpretl_tt06_tdc_v2_93.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1314 VPWR net43 a_9963_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1315 a_9849_12559 a_8859_12559 a_9723_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1316 a_11697_13647 tdc0.w_ring_buf24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1317 _010_ _147_ a_9025_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X1318 VPWR _054_ a_26483_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1322 VPWR tdc1.r_ring_ctr9 a_21327_10071 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1323 tdc1.r_dly_store_ring8 a_21391_15003 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1325 a_21164_12559 a_20249_12559 a_20817_12801 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1327 a_21445_18549 a_21279_18549 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1328 a_25190_10749 a_24113_10383 a_25028_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1329 uo_out[4] a_14032_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X1330 a_23542_17429 a_23374_17455 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1331 a_3962_16367 a_3689_16373 a_3877_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1332 tdc1.r_dly_store_ctr10 a_23967_10901 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1334 VGND tdc0.w_ring_int_norsz3 tdc0.w_ring_norsz3 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1335 _076_ a_13735_21263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1336 a_29101_19337 tdc1.w_ring_int_norsz14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1338 VPWR a_21337_14165 _196_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X1339 a_24696_15823 a_24297_15823 a_24570_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1340 VGND a_23996_16599 _099_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X1341 VGND net35 a_23211_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1342 VGND a_7775_20443 a_7733_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1343 VPWR a_16658_15279 a_16764_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X1344 VGND _197_ _035_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1347 VPWR a_4165_11989 a_4055_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1348 VPWR a_23799_10927 a_23967_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1349 VGND a_13755_13077 a_13713_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1350 a_23193_20725 a_23027_20725 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1351 VGND net26 a_5639_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1352 tdc0.r_dly_store_ring21 a_9799_16091 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1353 a_11783_10927 a_11159_10933 a_11675_11305 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1354 VGND a_29435_15797 a_29442_16097 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1355 VGND net10 a_23947_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1356 a_11863_10217 a_11417_9845 a_11767_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1357 _006_ _165_ a_1297_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X1360 VGND tdc1.w_ring_int_norsz31 tdc1.w_ring_norsz31 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1361 a_13897_18863 tdc0.r_dly_store_ring13 a_13459_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1363 a_30093_14197 a_29927_14197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1364 VGND a_14032_16911 uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X1367 a_9424_12559 a_9025_12559 a_9298_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1368 tdc0.w_ring_buf31 a_6007_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1370 VPWR a_10018_14847 a_9945_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1371 a_23907_21237 net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X1372 VPWR a_28047_21237 net43 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1373 a_16941_15279 a_16764_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1374 VGND a_15750_16885 a_15679_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1376 VGND a_19899_18543 net15 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1377 tdc1.r_dly_store_ctr3 a_30959_14165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1378 VPWR _197_ _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1379 VGND a_27135_15797 a_27142_16097 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1380 VPWR _135_ a_14075_19747 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1381 _197_ a_5087_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1382 a_14804_21263 tdc1.r_dly_store_ring7 a_14583_21590 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1383 a_24849_20719 tdc1.w_ring_norsz17 a_24765_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1387 VGND net9 a_15851_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1389 a_8197_13109 a_8031_13109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1391 a_5791_12533 _149_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X1392 VPWR a_15262_13759 a_15189_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1393 VGND _192_ a_17638_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1396 tdc1.w_ring_int_norsz23 tdc1.w_ring_norsz22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1398 tdc0.w_ring_norsz23 tdc0.w_ring_int_norsz23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1399 VPWR tdc1.r_ring_ctr6 a_23363_12711 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1400 a_10145_10625 a_9927_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1401 VGND net14 tdc1.w_ring_norsz23 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1402 _005_ _165_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1403 a_13921_19747 _136_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1404 VPWR _177_ a_22711_12533 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1406 VGND a_7079_11231 a_7013_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1407 VGND _064_ a_24631_16891 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.118 ps=1.4 w=0.42 l=0.15
X1408 a_11582_11989 a_11414_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1409 VPWR tdc1.r_ring_ctr0 a_28241_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1410 VGND a_9155_15253 a_9113_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1411 a_6687_14191 a_5989_14197 a_6430_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1412 VGND a_15543_16885 a_15550_17185 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1413 VGND tdc0.w_ring_norsz23 a_11067_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1414 a_10705_18543 tdc0.w_ring_norsz23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1415 VGND _039_ a_6601_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1416 VGND tdc1.w_ring_norsz3 tdc1.w_ring_int_norsz4 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1417 a_13323_11159 tdc0.r_ring_ctr2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X1418 VGND _176_ _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1419 net41 a_26031_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1420 tdc0.w_ring_norsz7 net22 a_10049_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1421 a_6913_15823 tdc0.w_ring_buf29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1422 tdc1.w_ring_norsz12 tdc1.w_ring_norsz28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1423 VGND a_18298_19605 a_18256_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1424 a_11049_17999 a_10883_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1425 a_30492_16745 a_30093_16373 a_30366_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1426 a_25103_16599 tdc1.r_dly_store_ctr2 a_25229_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1427 _161_ _156_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1428 VGND tdc1.w_ring_int_norsz6 tdc1.w_ring_norsz6 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1429 VPWR a_23211_12015 _179_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1430 a_11463_12925 a_10681_12559 a_11379_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1431 VPWR tdc1.w_dly_stop3 a_16311_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1432 tdc1.w_ring_buf8 a_20083_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1433 a_17720_15279 _191_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X1434 VPWR a_12007_17179 a_11923_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1435 a_28043_15511 a_28139_15511 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1436 VGND a_16727_20951 tdc1.r_dly_store_ring7 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1437 uo_out[7] a_14172_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1438 tdc1.r_dly_store_ring19 a_21299_17179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1439 a_12989_16687 tdc0.r_dly_store_ring17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1444 VPWR a_17804_15279 uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1445 a_14280_15599 _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1447 a_16919_10383 a_16569_10383 a_16824_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1448 VPWR a_17267_16367 a_17435_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1449 a_5875_13077 tdc0.r_ring_ctr11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X1450 VGND _142_ a_14994_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1451 tdc0.r_dly_store_ring3 a_11271_16091 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1452 a_14197_15279 tdc0.r_dly_store_ring18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1454 _073_ a_12907_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1456 a_9021_13481 a_8031_13109 a_8895_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1457 a_28823_14557 tdc1.r_ring_ctr1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1458 VGND a_17267_16367 a_17435_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1459 a_14760_13481 a_14361_13109 a_14634_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1460 a_6633_10383 a_6467_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1461 a_7669_14985 tdc0.w_ring_norsz26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1464 a_13713_13481 a_12723_13109 a_13587_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1465 a_30442_12381 _049_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1466 _030_ a_23403_9839 a_23653_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1467 a_1552_13469 _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1468 a_28139_15511 a_28423_15497 a_28358_15645 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1469 VGND net29 a_10239_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1470 a_16535_20502 a_16353_20502 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1471 VGND a_5935_19355 a_5893_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1473 VPWR a_24915_15511 tdc1.r_dly_store_ring16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1474 _032_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1476 VPWR a_6119_17179 a_6035_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1477 VPWR a_26667_21237 net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1478 a_14372_18543 _126_ a_14195_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1479 VGND a_15595_20693 a_15553_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1480 VPWR a_22247_20938 tdc1.w_ring_buf17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R19 net54 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1482 a_12805_18543 net24 a_12889_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1483 VPWR a_4595_11231 tdc0.r_ring_ctr8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1484 a_4157_18543 net19 tdc0.w_ring_norsz16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1486 a_22247_20938 tdc1.w_ring_norsz17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1487 a_11540_15657 a_11141_15285 a_11414_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1488 VGND a_9431_17179 a_9389_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1489 VGND a_21327_10071 _181_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1490 a_18703_14735 _080_ a_18881_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1491 a_14159_10217 a_13643_9845 a_14064_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1492 VPWR a_17468_15797 _079_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1493 a_3951_11305 a_3505_10933 a_3855_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1494 a_30307_18921 a_30178_18665 a_29887_18775 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1495 VPWR a_19402_16341 a_19329_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1496 VGND a_9103_12247 _149_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1497 VPWR a_13019_12827 a_12935_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1498 VGND a_23063_14013 a_23231_13915 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1499 a_3904_15823 a_3505_15823 a_3778_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1500 net3 a_28415_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1501 a_30554_18543 a_30307_18921 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1504 tdc0.r_ring_ctr10 a_2387_13407 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1505 VPWR net9 a_16403_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1507 tdc0.w_ring_norsz8 tdc0.w_ring_norsz24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1508 a_17213_14985 tdc0.r_dly_store_ring0 a_17129_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1509 VGND _067_ a_25643_18775 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.118 ps=1.4 w=0.42 l=0.15
X1510 a_17267_16367 a_16403_16373 a_17010_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1512 a_5069_19087 a_4903_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1513 a_6204_13647 a_5805_13647 a_6078_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1514 a_8933_20725 a_8767_20725 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1516 a_12875_20327 _083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X1517 tdc0.w_ring_norsz31 net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1518 a_11329_12015 tdc0.r_ring_ctr5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1520 a_8010_14191 a_7737_14197 a_7925_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1521 VGND a_27259_19087 _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1523 a_25126_14191 a_24879_14569 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1524 VPWR tdc1.w_ring_norsz12 a_28271_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1525 a_5602_15935 a_5434_16189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1527 a_25099_14557 a_24879_14569 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X1528 tdc1.w_ring_buf19 a_19991_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1529 _159_ a_3431_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1530 VPWR _183_ _184_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1531 VPWR a_4512_13481 a_4687_13407 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1532 VPWR net36 a_29927_15285 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1533 a_18939_20327 tdc1.r_dly_store_ring14 a_19065_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1534 a_9121_15823 tdc0.w_ring_buf21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1535 a_26297_20340 tdc1.w_ring_norsz0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1536 VGND a_27159_11989 a_27090_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1537 a_26031_16885 net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X1539 VPWR net7 a_1131_14197 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1540 VGND net28 a_7571_14197 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1541 a_17208_20149 _078_ a_18030_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1542 a_21666_14191 _194_ a_21586_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X1543 tdc0.w_ring_int_norsz19 tdc0.w_ring_norsz18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1544 a_27621_18909 a_27351_18543 a_27517_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1545 VPWR a_22143_12015 a_22311_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1546 tdc0.w_ring_norsz21 tdc0.w_ring_int_norsz21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1547 VGND a_12867_15511 _130_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1548 a_3689_16373 a_3523_16373 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1549 VGND net34 a_21739_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1550 a_13349_19631 tdc0.r_dly_store_ring31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1551 VGND a_22143_12015 a_22311_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1552 tdc1.w_ring_int_norsz10 tdc1.w_ring_norsz9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1553 a_26851_15797 a_27142_16097 a_27093_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1554 a_28721_19631 net78 tdc1.w_ring_int_norsz31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1555 VPWR tdc1.r_dly_store_ring18 a_24397_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X1558 VGND _185_ a_17967_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1559 VPWR a_1957_17153 a_1847_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1561 VPWR tdc1.r_ring_ctr1 a_28361_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R20 VPWR tdc1.g_ring316.stg01_63.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1562 a_11141_16911 a_10975_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1563 a_16656_16885 _095_ a_17478_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1564 VGND a_3483_14423 _004_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1565 VGND tdc1.w_ring_int_norsz29 tdc1.w_ring_norsz29 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1568 tdc0.r_dly_store_ctr11 a_6855_14165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1569 a_24209_14735 tdc1.r_ring_ctr7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1570 VGND tdc0.w_ring_norsz8 tdc0.w_ring_norsz24 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1572 a_22143_18543 a_21445_18549 a_21886_18517 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1574 VGND a_11763_11445 _147_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1575 VPWR net10 a_29191_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1577 a_19057_12015 tdc1.r_ring_ctr13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1579 VGND a_19338_21237 a_19267_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1580 a_30378_18820 a_30171_18761 a_30554_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1583 a_23925_17833 a_22935_17461 a_23799_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1586 VGND a_24950_14468 a_24879_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1587 a_19609_14191 tdc1.w_ring_buf24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1588 VPWR a_10995_20443 a_10911_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1589 a_7465_18543 tdc0.w_ring_buf13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1592 a_22143_12015 a_21279_12021 a_21886_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1594 a_17967_12559 tdc1.r_ring_ctr14 a_17861_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1595 a_24087_18775 tdc0.r_dly_store_ring30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.141 ps=1.33 w=0.42 l=0.15
X1596 a_5253_16911 a_5087_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1598 a_24950_14468 a_24743_14409 a_25126_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X1600 a_27397_12381 _054_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X1603 VGND a_4279_17179 a_4237_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1605 VGND tdc0.w_ring_int_norsz19 tdc0.w_ring_norsz19 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1606 VGND a_21886_11989 a_21844_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1607 VPWR a_7723_10357 a_7710_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1608 VPWR a_24743_14409 a_24750_14313 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1609 a_26961_12381 a_26483_11989 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X1610 a_21331_10901 tdc1.r_ring_ctr8 a_21729_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X1611 a_28425_16911 a_27871_16885 a_28078_16885 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1612 VGND _177_ a_22353_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1613 VPWR tdc0.r_ring_ctr10 a_1129_12809 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1614 _008_ _145_ a_14017_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1615 VPWR net35 a_23211_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1618 VPWR tdc0.w_ring_norsz5 a_9309_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1619 a_14361_13109 a_14195_13109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1620 a_17819_17455 a_16955_17461 a_17562_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1624 a_22375_15395 _107_ a_22293_15395 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1625 uo_out[2] a_16656_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1626 a_19153_18249 net14 tdc1.w_ring_norsz5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1627 a_19573_10383 a_19529_10625 a_19407_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
R21 uio_out[6] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1628 tdc0.r_dly_store_ring25 a_15227_13077 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1629 tdc1.w_ring_buf8 a_20083_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1630 a_17489_17455 a_16955_17461 a_17394_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1631 a_11839_17277 a_11141_16911 a_11582_17023 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1633 a_23996_16599 _096_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X1634 _153_ tdc0.r_ring_ctr6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1635 tdc0.r_dly_store_ring25 a_15227_13077 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1637 a_11414_17277 a_10975_16911 a_11329_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1638 VPWR a_25971_18551 _067_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1639 VGND a_4555_16341 a_4513_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1640 a_13861_17161 _112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1641 VGND a_12007_11989 a_11965_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1642 VGND tdc1.r_ring_ctr3 a_29099_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1643 VGND a_27003_11169 a_26964_11043 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1644 VPWR a_6059_11989 _156_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1645 a_21326_12925 a_20249_12559 a_21164_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1647 a_16991_18543 a_16127_18549 a_16734_18517 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1648 VGND _085_ a_22160_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1650 a_26321_15101 a_25787_14735 a_26226_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1651 a_29877_12559 a_29833_12801 a_29711_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1652 a_12426_12925 a_11987_12559 a_12341_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1654 tdc0.r_dly_store_ring8 a_17159_14165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1656 VPWR a_19951_11159 _018_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X1659 VGND tdc1.r_dly_store_ring22 a_19165_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1660 a_24131_18249 _067_ a_24385_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1661 VGND _043_ a_4209_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1663 a_16661_18543 a_16127_18549 a_16566_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1664 VPWR _031_ a_27722_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1665 VPWR a_22771_21531 a_22687_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1666 VPWR a_25381_17429 _086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X1668 a_26394_14847 a_26226_15101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1669 VGND tdc0.w_ring_norsz28 tdc0.w_ring_int_norsz29 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1670 tdc0.r_dly_store_ring23 a_12375_19605 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1671 VPWR a_30791_15279 a_30959_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1673 VPWR a_19735_11989 a_19651_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1674 _187_ a_17586_12335 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1676 a_4195_17277 a_3413_16911 a_4111_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1677 _074_ a_26754_19133 a_27017_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X1679 tdc0.w_ring_buf3 a_10147_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1680 _180_ tdc1.r_ring_ctr8 a_25321_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1681 a_18225_19337 tdc1.w_ring_norsz6 a_18141_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1682 a_24559_10383 a_24113_10383 a_24463_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1683 VPWR a_30263_12319 a_30250_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1685 a_22653_20425 _083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X1687 a_1755_14191 _044_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1688 VPWR a_26819_15003 a_26735_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1689 VPWR tdc1.r_dly_store_ctr0 a_22741_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X1690 a_5526_17277 a_5087_16911 a_5441_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1691 uo_out[6] a_13344_20693 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1694 a_10570_20287 a_10402_20541 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1695 a_17049_10159 _185_ _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.25 ps=1.42 w=0.65 l=0.15
X1696 a_29711_12559 a_29265_12559 a_29615_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1697 VGND a_10827_20541 a_10995_20443 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1698 a_24920_11471 a_24694_11517 a_24551_11623 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1699 a_15143_13103 a_14361_13109 a_15059_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1700 a_22304_16911 a_21905_16911 a_22178_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1701 tdc1.w_ring_int_norsz30 net77 a_28829_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1702 tdc0.w_ring_norsz20 net21 a_10325_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1703 _024_ _168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1704 VPWR a_27815_17429 a_27346_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1705 VPWR a_14583_18267 a_14499_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1707 a_12723_17161 _069_ a_12805_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1708 tdc0.w_ring_int_norsz24 net53 a_10705_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1709 _193_ a_20635_13897 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1710 a_24845_14735 a_23855_14735 a_24719_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1711 VGND tdc1.w_ring_norsz10 tdc1.w_ring_norsz26 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1713 a_18239_16073 _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1714 a_21718_18543 a_21445_18549 a_21633_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1715 a_24915_15511 a_25011_15511 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1716 a_25287_18517 net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.146 ps=1.34 w=0.42 l=0.15
X1717 VPWR a_4443_18543 net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1718 VPWR a_15904_11445 _624_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1719 a_26483_11989 a_26686_12147 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X1720 a_24481_12021 a_24315_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1721 tdc0.w_ring_int_norsz16 net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1722 a_11601_19087 a_11435_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1723 a_22595_14887 tdc1.r_dly_store_ring16 a_22741_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1724 tdc1.w_ring_buf26 a_23671_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1725 tdc0.w_ring_norsz30 net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1726 VPWR a_13344_20693 uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X1727 tdc0.r_ring_ctr0 a_12507_10143 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1729 VPWR a_27127_16885 net18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1730 a_12291_19631 a_11509_19637 a_12207_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1731 _163_ tdc0.r_ring_ctr13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1732 a_26805_20425 tdc1.w_ring_norsz15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1733 a_7205_17455 tdc0.w_ring_int_norsz13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1734 a_15170_19605 a_15002_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1736 a_7423_16189 a_6725_15823 a_7166_15935 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1739 VGND a_23799_10927 a_23967_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1740 _019_ a_16831_9813 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1741 tdc0.w_ring_norsz3 tdc0.w_ring_norsz19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1743 VGND tdc1.w_ring_norsz12 a_28271_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1744 VGND tdc0.r_ring_ctr4 a_8775_10633 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1745 VPWR a_23155_19453 a_23323_19355 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1746 tdc1.w_ring_buf19 a_19991_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1747 VPWR a_26394_14847 a_26321_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1749 a_15151_19453 a_14453_19087 a_14894_19199 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1750 VGND a_20874_17023 a_20832_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1751 VPWR _075_ a_13993_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1752 tdc1.w_dly_stop3 a_15759_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1753 VPWR a_16734_18517 a_16661_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1754 tdc0.w_ring_buf16 a_5087_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1755 VGND net34 a_23027_20725 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1756 a_12042_19199 a_11874_19453 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1757 a_15009_13647 tdc0.w_ring_buf9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1758 a_1297_16687 tdc0.r_ring_ctr15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1759 a_26919_18863 a_26627_18543 a_26833_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1760 a_24420_14735 a_24021_14735 a_24294_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R22 uio_oe[5] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1761 a_14377_9813 a_14159_10217 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1762 a_26830_18249 _123_ a_26581_18145 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X1764 tdc0.r_ring_ctr1 a_14899_10143 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X1765 a_29523_12393 a_29173_12021 a_29428_12381 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1766 VGND a_11122_12671 a_11080_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1767 a_17043_16073 _075_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1769 a_25049_11989 a_24831_12393 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1770 a_10593_15823 tdc0.w_ring_buf3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1771 uo_out[4] a_14032_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1772 VGND _041_ a_4209_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1773 a_16175_20938 net12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1775 VGND a_4111_17277 a_4279_17179 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1776 net43 a_28047_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1778 a_16475_12925 a_15851_12559 a_16367_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1779 _080_ a_19860_15797 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1780 _072_ a_24635_17973 a_24385_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1781 VGND a_23783_19605 a_23741_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1782 net15 a_19899_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X1783 VPWR a_30791_14191 a_30959_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1784 a_16523_15101 a_15741_14735 a_16439_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1785 a_22469_15823 _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X1786 VPWR net3 a_13735_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1787 VPWR a_3485_15253 _164_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1789 a_4165_13077 a_3947_13481 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1790 a_8850_11247 _147_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
R23 tt_um_hpretl_tt06_tdc_v2_88.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1791 a_18555_19631 a_17857_19637 a_18298_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1793 VGND net74 tdc1.w_ring_int_norsz27 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1795 a_2703_10927 _156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1796 VGND _130_ a_12618_21039 VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.101 ps=0.96 w=0.65 l=0.15
X1797 VGND _071_ a_13253_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1798 VPWR tdc1.r_dly_store_ring29 a_27517_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
R24 VPWR tdc0.g_ring325.stg01_54.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1799 VPWR a_11915_15003 a_11831_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1800 tdc1.w_ring_buf18 a_21647_20719 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1801 VGND tdc0.w_ring_norsz22 tdc0.w_ring_int_norsz23 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1802 VGND a_23542_10901 a_23500_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X1803 VPWR a_25571_13621 a_25558_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1804 VPWR a_17727_14013 a_17895_13915 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1805 a_22653_20425 _075_ a_22855_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1807 a_28538_20996 a_28338_20841 a_28687_21085 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1808 VGND _069_ a_13897_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1810 VGND a_23403_9839 _030_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X1811 a_27095_13345 net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1812 tdc1.w_ring_int_norsz4 net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1813 a_10049_19337 tdc0.w_ring_norsz23 a_9965_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1814 VPWR a_9647_15253 net26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1816 VGND net17 tdc1.w_ring_norsz12 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1817 VPWR a_30515_17455 a_30683_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1818 VPWR a_23259_18164 tdc1.w_ring_buf25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1820 VPWR a_30447_13621 a_30434_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1822 VPWR a_21391_15003 a_21307_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1823 _179_ a_23211_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1824 tdc1.w_ring_norsz6 tdc1.w_ring_norsz22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1825 a_11379_12925 a_10515_12559 a_11122_12671 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1826 VGND a_30515_17455 a_30683_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1827 a_24459_14423 a_24743_14409 a_24678_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1828 a_17777_11247 _184_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1829 a_4055_12015 a_3431_12021 a_3947_12393 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1830 VGND a_14172_20149 uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1832 _131_ a_12618_21039 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.275 ps=1.5 w=0.65 l=0.15
X1834 _122_ a_27517_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X1835 a_24297_15823 a_24131_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1836 a_11782_14013 a_11343_13647 a_11697_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1837 a_9832_10383 _010_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1838 a_23147_14013 a_22365_13647 a_23063_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1840 a_24455_17687 _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X1841 VGND a_23967_17429 a_23925_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1842 a_11049_12925 a_10515_12559 a_10954_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1843 a_27693_18909 _065_ a_27621_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X1844 a_16919_10383 a_16403_10383 a_16824_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1845 VGND a_16155_15975 _070_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1846 tdc1.r_ring_ctr8 a_25203_10357 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X1847 a_11923_15279 a_11141_15285 a_11839_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1848 a_6725_15823 a_6559_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1850 a_11329_16911 tdc0.w_ring_buf18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1852 a_21527_11293 _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X1853 a_24451_18864 _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1855 VPWR tdc1.w_ring_norsz30 a_28721_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1856 a_9374_20693 a_9206_20719 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1858 a_16607_20502 tdc0.r_dly_store_ring1 a_16607_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1860 a_15659_16483 _077_ a_15577_16483 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1862 VPWR a_11490_14847 a_11417_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X1864 VGND net7 a_6467_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1867 VGND net10 a_29191_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1868 VPWR net29 a_14563_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1869 a_28423_15497 net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1870 VGND net18 tdc1.w_ring_norsz0 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1871 VPWR tdc1.w_ring_int_norsz3 a_20249_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1872 a_14724_10217 a_13643_9845 a_14377_9813 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1873 VPWR a_7079_11231 a_7066_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1874 VPWR a_22995_10357 a_22982_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1875 a_12391_21629 a_11693_21263 a_12134_21375 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1877 a_18049_16367 _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1878 VGND a_30378_18820 a_30307_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X1879 VGND net32 a_14563_19637 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1880 a_23883_10927 a_23101_10933 a_23799_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1881 VPWR a_26031_16885 net41 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1884 VPWR tdc0.w_ring_norsz10 a_9135_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1885 a_25229_16367 _068_ a_25431_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1886 net5 a_26667_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1887 a_7166_19605 a_6998_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1888 a_14894_19199 a_14726_19453 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1891 a_23101_17461 a_22935_17461 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1894 a_24681_10625 a_24463_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1895 a_17217_13647 tdc1.r_ring_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1896 a_20175_16073 _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X1897 a_30515_17455 a_29651_17461 a_30258_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X1898 a_12889_18543 tdc0.r_dly_store_ring12 a_12805_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1900 tdc1.w_ring_int_norsz2 tdc1.w_ring_norsz1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1901 a_16481_14191 tdc0.w_ring_buf8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1902 VGND net61 tdc0.w_ring_int_norsz0 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1904 a_5985_15823 a_4995_15823 a_5859_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1905 a_1297_13109 a_1131_13109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1906 VPWR a_9503_12015 net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1909 _079_ a_17468_15797 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1910 a_6796_17973 net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1911 VPWR tdc1.r_ring_ctr11 a_20819_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1912 a_8964_16911 a_8565_16911 a_8838_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1913 a_30185_17455 a_29651_17461 a_30090_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1915 VPWR a_25839_16341 net25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1916 _053_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1919 a_29707_13647 a_29357_13647 a_29612_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1920 a_5353_12381 _147_ a_5271_12128 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1921 a_16585_12801 a_16367_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1922 VGND net22 tdc0.w_ring_norsz8 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1923 a_5875_13077 tdc0.r_ring_ctr9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X1924 VPWR a_22135_14423 _107_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1925 a_17129_14985 _076_ a_17047_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1926 VPWR tdc1.w_ring_norsz21 a_19071_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1927 a_27469_12381 a_27090_12015 a_27397_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1928 net14 a_18243_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1930 a_21095_11471 tdc1.r_ring_ctr10 a_20989_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1931 VGND net26 a_5823_14197 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1932 VPWR net27 a_8767_20725 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1934 VGND tdc1.w_ring_norsz25 tdc1.w_ring_norsz9 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1936 a_25571_12319 _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1937 VGND tdc1.w_dly_stop5 a_28915_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1939 a_26141_14735 tdc1.r_ring_ctr5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1940 VGND a_27951_20951 tdc1.r_dly_store_ring15 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1942 a_6998_16189 a_6559_15823 a_6913_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1943 VGND a_30791_16367 a_30959_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1944 tdc0.w_ring_norsz17 net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1945 a_19131_21237 net34 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1948 a_22447_15395 _106_ a_22375_15395 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1949 a_27346_17687 tdc1.r_dly_store_ctr5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X1950 a_4687_13407 _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1951 _017_ a_21103_10633 a_21353_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1952 VGND _059_ a_19573_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1953 a_6018_11517 _156_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X1954 VPWR _197_ _032_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1956 VGND a_22595_14887 _195_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1957 a_30281_15279 tdc1.r_ring_ctr2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1958 tdc0.r_dly_store_ring1 a_15595_20693 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1959 uo_out[5] a_14372_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.172 ps=1.83 w=0.65 l=0.15
X1965 VGND tdc0.w_ring_int_norsz26 tdc0.w_ring_norsz26 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1966 VPWR _198_ _057_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1967 tdc1.w_ring_norsz16 net62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1968 a_25678_15279 a_25431_15657 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1971 a_10846_15935 a_10678_16189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X1973 a_10018_14847 a_9850_15101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X1974 tdc0.w_ring_norsz1 tdc0.w_ring_int_norsz1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1975 VGND _051_ a_29877_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1976 a_3855_11305 a_3505_10933 a_3760_11293 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1977 a_29055_15975 a_29151_15797 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1978 a_18206_11471 _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1979 a_18225_19631 a_17691_19637 a_18130_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X1980 VPWR _161_ a_3786_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1981 VPWR a_28599_15797 net36 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1982 VPWR net31 a_10975_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1983 VGND tdc1.r_ring_ctr2 a_28609_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1984 VGND a_6671_13915 a_6629_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1986 a_17478_16911 _099_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X1987 a_6909_20175 a_6743_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1988 a_24368_10383 _030_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1989 VGND _047_ a_2001_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1990 tdc0.w_ring_buf31 a_6007_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1992 VGND net55 tdc0.w_ring_int_norsz26 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1993 a_12529_14191 tdc0.r_dly_store_ring24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1997 VPWR _170_ a_22199_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1998 VGND tdc1.r_dly_store_ring10 a_24685_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1999 a_25839_16341 _066_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2000 uo_out[1] a_17208_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2002 a_19693_12393 a_18703_12021 a_19567_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2003 tdc0.r_ring_ctr0 a_12507_10143 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2004 VPWR tdc0.r_dly_store_ctr1 a_16301_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2006 tdc0.w_ring_norsz24 tdc0.w_ring_int_norsz24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2007 a_13530_12015 a_13091_12021 a_13445_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2008 a_26627_18543 _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X2009 VPWR a_30258_17429 a_30185_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2010 VGND net15 tdc1.w_ring_norsz18 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2012 _040_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2013 VPWR tdc0.r_ring_ctr4 a_9103_12247 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2014 a_17586_12335 tdc1.r_ring_ctr12 a_17500_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X2016 a_3505_15823 a_3339_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2018 a_13091_14191 _080_ a_13173_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2019 a_6244_11471 tdc0.r_ring_ctr7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2020 a_12134_21375 a_11966_21629 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2021 VPWR a_26581_18145 _124_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
X2022 tdc0.w_ring_buf5 a_10331_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2023 tdc1.r_ring_ctr3 a_30355_12533 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2025 a_8086_17429 a_7918_17455 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2027 _054_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2028 a_25750_13647 _053_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2029 tdc0.r_dly_store_ring24 a_12375_13915 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2030 VGND net16 a_19899_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2032 VGND _116_ a_13948_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2034 a_30626_13647 _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2037 VPWR a_11582_11989 a_11509_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2038 VPWR net27 a_5087_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2040 a_2566_14557 _044_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2041 VGND a_18027_11445 a_17961_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2042 tdc0.w_ring_norsz19 tdc0.w_ring_norsz3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2043 a_28731_13103 tdc1.r_ring_ctr1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X2044 a_13091_14191 _080_ a_13173_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2045 tdc0.w_ring_int_norsz2 net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2046 VPWR tdc1.w_ring_norsz31 a_26983_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2047 a_21353_10383 tdc1.r_ring_ctr10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2048 a_1129_12809 _158_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2049 a_19452_15657 a_19053_15285 a_19326_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2050 a_28779_15645 a_28559_15657 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2051 a_12805_16911 tdc0.r_dly_store_ring28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2052 VPWR a_28331_20937 a_28338_20841 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2054 a_13990_18365 a_13717_17999 a_13905_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2055 a_12815_17455 _071_ a_12897_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2056 VPWR net30 a_14195_13109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2057 a_6998_16189 a_6725_15823 a_6913_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2058 a_11950_13759 a_11782_14013 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2059 tdc1.w_ring_int_norsz16 net63 a_26805_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2061 a_22741_14985 _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2062 a_1847_17277 a_1223_16911 a_1739_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2063 a_13785_20203 _075_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2065 a_4055_13103 _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2066 VPWR a_15059_13103 a_15227_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2067 VGND tdc1.w_ring_buf12 a_29989_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2069 tdc1.w_ring_int_norsz6 net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2071 tdc0.w_ring_buf25 a_11067_13103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2072 a_7737_14197 a_7571_14197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2073 VGND a_27772_16341 net17 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2074 VGND a_15059_13103 a_15227_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2075 _067_ a_25971_18551 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2076 tdc0.r_dly_store_ring12 a_8511_17429 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2077 VPWR a_18298_19605 a_18225_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2078 a_8841_11471 a_8675_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2079 a_6725_13109 a_6559_13109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2080 _156_ a_6059_11989 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2081 a_1647_14569 a_1297_14197 a_1552_14557 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2082 VGND net56 tdc0.w_ring_int_norsz27 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2085 tdc0.r_dly_store_ring12 a_8511_17429 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2086 VPWR net31 a_11343_19637 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2087 a_27090_10927 a_26964_11043 a_26686_11059 VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2088 VGND tdc0.w_ring_norsz24 tdc0.w_ring_int_norsz25 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2089 a_26635_17775 tdc1.r_dly_store_ring11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
X2090 VGND a_30447_13621 a_30381_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2091 VGND tdc1.w_ring_buf27 a_27689_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2092 VPWR a_30423_18365 a_30591_18267 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2094 tdc0.r_dly_store_ctr8 a_7591_13077 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2096 a_1865_14165 a_1647_14569 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2097 VPWR a_22311_18517 a_22227_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2099 VPWR a_12207_19631 a_12375_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2100 a_4420_11305 a_3339_10933 a_4073_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2101 tdc0.r_dly_store_ctr8 a_7591_13077 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2102 a_7989_11499 _149_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2103 a_29833_12801 a_29615_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2105 tdc0.w_ring_int_norsz29 net58 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2106 VGND a_12207_19631 a_12375_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2107 a_4529_14735 a_3339_14735 a_4420_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2109 a_29619_12393 a_29173_12021 a_29523_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2110 VGND a_11271_16091 a_11229_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2111 a_28007_16911 a_27871_16885 a_27587_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2113 a_30917_14569 a_29927_14197 a_30791_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2114 a_30423_18365 a_29725_17999 a_30166_18111 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2115 a_23996_16599 _098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2116 VPWR tdc1.w_ring_int_norsz15 a_28621_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2117 _162_ a_5791_12533 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X2119 VGND net16 _059_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2121 a_29151_15797 a_29435_15797 a_29370_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X2122 VGND tdc1.w_ring_norsz21 a_19071_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2123 a_29641_16367 net42 tdc1.w_ring_int_norsz12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2125 VGND tdc0.w_ring_norsz10 a_9135_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2126 a_27012_13103 a_26575_13077 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
R25 VPWR tt_um_hpretl_tt06_tdc_v2_95.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2127 a_5993_13647 tdc0.r_ring_ctr10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2128 a_13895_11471 tdc0.r_ring_ctr2 a_13799_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X2129 a_3295_19252 net27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2130 a_13861_17161 _089_ a_14032_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2131 VPWR a_27307_14887 tdc1.r_dly_store_ctr0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2132 a_14726_19453 a_14453_19087 a_14641_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2133 a_20051_10357 a_19876_10383 a_20230_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2134 VGND _076_ a_16828_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X2135 a_15059_13103 a_14195_13109 a_14802_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2136 VPWR a_30378_18820 a_30307_18921 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2137 a_11417_18365 a_10883_17999 a_11322_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2138 VPWR net7 a_5823_10933 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2139 VPWR net5 a_25971_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2141 VPWR a_28064_11471 a_28239_11445 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2142 a_23466_20719 a_23027_20725 a_23381_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2145 tdc0.r_dly_store_ring4 a_14583_18267 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2146 VGND tdc1.r_ring_ctr6 a_22905_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X2148 a_11490_18111 a_11322_18365 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2149 VPWR a_12042_19199 a_11969_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2150 tdc0.w_ring_norsz5 tdc0.w_ring_norsz21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2152 a_11237_14735 tdc0.w_ring_buf26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2153 VPWR a_26615_13647 net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2155 a_29370_20175 a_29055_20327 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2156 VGND net10 a_24315_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2157 tdc0.w_ring_buf4 a_12355_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
R26 VGND net48 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2158 a_7507_13103 a_6725_13109 a_7423_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2159 a_30355_12533 a_30180_12559 a_30534_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2160 VPWR net29 a_11343_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2161 VGND net31 a_11435_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2162 a_5894_15101 a_5455_14735 a_5809_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2163 a_26297_20340 tdc1.w_ring_norsz0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2164 net18 a_27127_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2165 a_12207_19631 a_11343_19637 a_11950_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2166 a_4537_18249 tdc0.w_ring_int_norsz16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2167 a_7691_20541 a_6909_20175 a_7607_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2168 a_16585_12801 a_16367_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2170 VPWR net35 a_22935_17461 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2174 VPWR a_4420_11305 a_4595_11231 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2175 a_23155_19453 a_22457_19087 a_22898_19199 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2176 a_8775_10633 _147_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2179 VGND a_8603_14165 a_8561_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2180 a_9206_16189 a_8933_15823 a_9121_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2182 tdc1.w_ring_norsz20 tdc1.w_ring_norsz4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2183 VGND a_11582_15253 a_11540_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2184 VGND a_22771_17179 a_22729_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2185 _066_ a_24822_19133 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X2187 VGND tdc0.w_ring_norsz6 tdc0.w_ring_int_norsz7 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2188 a_17428_13647 a_17029_13647 a_17302_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2190 a_2505_15823 a_1315_15823 a_2396_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2191 a_11782_19631 a_11343_19637 a_11697_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2193 VGND tdc0.w_ring_norsz12 tdc0.w_ring_int_norsz13 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2194 a_2212_14569 a_1131_14197 a_1865_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2195 a_14541_17999 a_13551_17999 a_14415_18365 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2196 VPWR _076_ a_14797_21590 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X2197 a_19973_19337 tdc1.w_ring_norsz8 a_19889_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2198 tdc1.r_ring_ctr13 a_18027_11445 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2199 a_23653_9839 tdc1.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2200 VGND net37 a_29559_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2202 a_27617_20719 net79 tdc1.w_ring_int_norsz0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2203 VGND a_28915_10927 _198_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2204 VGND _075_ a_13897_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X2205 a_6725_19637 a_6559_19637 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2207 a_10601_10383 a_9411_10383 a_10492_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2208 VGND a_18539_13077 a_18497_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2209 VGND a_1047_16367 _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X2210 a_14017_10633 _144_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2211 a_15741_14735 a_15575_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2212 a_6365_18249 net59 tdc0.w_ring_int_norsz30 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
R27 VPWR tdc0.g_ring323.stg01_52.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2213 a_6733_18543 net19 tdc0.w_ring_norsz14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2214 _166_ tdc0.r_ring_ctr14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.176 ps=1.84 w=0.65 l=0.15
X2216 VGND _076_ a_14804_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X2218 a_8767_10927 tdc0.r_ring_ctr4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X2219 _168_ a_28455_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X2220 tdc0.w_ring_norsz18 tdc0.w_ring_int_norsz18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2222 tdc0.r_dly_store_ring18 a_12007_17179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2223 a_27161_16367 tdc1.w_ring_norsz11 a_27077_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2224 a_26910_18249 _122_ a_26830_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X2225 a_30875_15279 a_30093_15285 a_30791_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2227 VPWR _197_ _041_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2228 a_16109_15101 a_15575_14735 a_16014_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2229 tdc1.w_ring_norsz13 net17 a_29185_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2230 a_20254_10927 _182_ a_19951_11159 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X2231 a_6166_12559 _154_ a_6070_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X2232 a_26352_14735 a_25953_14735 a_26226_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2234 a_20441_20425 net41 tdc1.w_ring_int_norsz3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2235 a_18869_12021 a_18703_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2238 tdc0.w_ring_norsz1 net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2239 a_20169_11247 _184_ a_19951_11159 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2240 VPWR a_4073_10901 a_3963_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2241 VGND _178_ a_23211_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2242 VPWR a_12559_21531 a_12475_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2243 tdc0.w_ring_int_norsz23 net52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R28 net61 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2244 tdc1.r_ring_ctr2 a_30447_13621 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2245 a_25558_14013 a_24481_13647 a_25396_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2246 a_14278_18543 _119_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.265 ps=2.53 w=1 l=0.15
X2247 a_16182_14847 a_16014_15101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2248 VGND a_2743_12711 _158_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X2249 VPWR a_22615_16599 _105_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X2250 a_28239_11445 a_28064_11471 a_28418_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2252 tdc0.w_ring_buf25 a_11067_13103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2253 net26 a_9647_15253 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2254 a_24743_14409 net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2255 a_9832_10383 _010_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2256 a_7159_17076 tdc0.w_ring_norsz29 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
R29 VPWR tt_um_hpretl_tt06_tdc_v2_86.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2257 VPWR a_10827_20541 a_10995_20443 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2258 a_17484_10383 a_16403_10383 a_17137_10625 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2259 a_22929_10383 a_21739_10383 a_22820_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2260 a_4203_16189 a_3339_15823 a_3946_15935 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2261 a_24363_14423 a_24459_14423 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2262 VPWR a_29642_15797 a_29571_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2263 a_26426_17687 a_26785_17687 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2264 a_18045_19631 tdc1.w_ring_buf6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2265 a_16293_18549 a_16127_18549 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2266 VGND _186_ a_17777_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X2269 a_13809_9545 tdc0.r_ring_ctr1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2270 a_23741_20009 a_22751_19637 a_23615_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2271 tdc0.r_dly_store_ring17 a_6119_17179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2272 tdc0.r_dly_store_ring30 a_17159_18517 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2273 VPWR a_13955_12015 a_14123_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2274 a_6909_20175 a_6743_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2275 tdc0.r_dly_store_ring30 a_17159_18517 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2276 VGND a_13955_12015 a_14123_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2278 a_13735_14191 _080_ a_13817_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2279 a_12889_13109 a_12723_13109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2282 a_6244_11471 a_6018_11517 a_5875_11623 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2283 VPWR a_14724_10217 a_14899_10143 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2285 a_11965_12393 a_10975_12021 a_11839_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2286 a_11509_15279 a_10975_15285 a_11414_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2287 VGND _068_ a_24477_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
R30 VGND net50 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2288 a_20249_19631 tdc1.w_ring_norsz19 a_20165_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2289 VGND a_28423_15497 a_28430_15401 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2290 a_5851_19453 a_5069_19087 a_5767_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2291 a_7066_10927 a_5989_10933 a_6904_11305 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2292 _151_ tdc0.r_ring_ctr5 a_8767_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2294 VPWR tdc1.w_dly_stop4 a_16587_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2295 a_6888_10383 _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2296 a_29612_13647 _024_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2298 a_23799_10927 a_22935_10933 a_23542_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2299 VGND net14 tdc1.w_ring_norsz4 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2303 a_13323_11159 tdc0.r_ring_ctr1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2304 a_19421_14197 a_19255_14197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2305 VPWR net11 a_15483_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2306 a_24275_16885 a_24631_16891 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2307 a_13735_14191 _080_ a_13817_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2308 VPWR a_6607_11623 _152_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2309 a_23937_15279 tdc1.r_dly_store_ctr15 a_23855_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2310 a_15170_11989 a_15002_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2311 a_20504_12559 _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2312 a_15741_14735 a_15575_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2313 VPWR _067_ a_26785_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X2314 a_23469_10927 a_22935_10933 a_23374_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2316 VPWR tdc1.r_ring_ctr9 a_20819_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X2317 a_6913_13103 tdc0.r_ring_ctr8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2318 tdc0.r_dly_store_ring16 a_6487_15003 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2319 a_14255_10217 a_13809_9845 a_14159_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2320 a_10317_20175 tdc0.w_ring_buf22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2321 a_5621_17277 a_5087_16911 a_5526_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2322 a_20547_18249 _124_ a_20451_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2323 VGND a_15687_13915 a_15645_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
R31 tdc0.g_ring328.stg01_57.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2324 a_3760_11293 _014_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2325 a_30875_14191 a_30093_14197 a_30791_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2326 VPWR a_2656_18517 _626_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2327 net25 a_25839_16341 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2328 VPWR a_26895_17429 a_26426_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2329 VGND _065_ _072_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2330 a_7653_16367 net22 tdc0.w_ring_norsz12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2331 VPWR a_15451_20149 _075_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2332 a_26686_11059 a_26964_11043 a_26920_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2333 a_17075_18543 a_16293_18549 a_16991_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2334 _049_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2335 _010_ a_8775_10633 a_9025_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X2337 a_8289_15285 a_8123_15285 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2339 a_15478_16911 a_15163_17063 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2340 VGND a_23264_21237 net34 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2341 net2 a_29559_21263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2342 VPWR a_14372_18543 uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X2344 a_25651_15645 a_25431_15657 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2345 a_27445_16367 tdc1.w_ring_int_norsz11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2346 VGND a_22603_21629 a_22771_21531 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R32 VPWR tdc1.g_ring330.stg01_77.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2348 a_10401_14735 a_9411_14735 a_10275_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2349 a_23937_15279 tdc1.r_dly_store_ctr7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2350 VPWR a_16180_21237 net31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2351 VGND a_13698_11989 a_13656_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2352 a_16301_16073 net25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2353 a_9585_17455 net39 tdc0.w_ring_int_norsz4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2354 tdc1.w_ring_norsz9 tdc1.w_ring_int_norsz9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2355 a_12521_12925 a_11987_12559 a_12426_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2356 a_26686_11059 a_27003_11169 a_26961_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2357 a_13323_11159 tdc0.r_ring_ctr1 a_13557_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
R33 tdc0.g_ring329.stg01_58.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2358 _083_ a_16187_19891 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2360 a_29817_17461 a_29651_17461 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2363 VGND a_30959_14165 a_30917_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2365 VGND net6 a_25251_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X2366 a_28559_15657 a_28430_15401 a_28139_15511 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2367 VGND tdc0.w_ring_norsz1 tdc0.w_ring_norsz17 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2368 VGND a_17159_18517 a_17117_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2369 VPWR tdc1.w_ring_buf1 a_19685_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2372 VPWR a_11582_17023 a_11509_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2373 tdc1.w_ring_buf26 a_23671_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2374 a_21647_16367 _083_ a_21729_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2375 VPWR a_15170_19605 a_15097_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2376 VPWR tdc0.w_ring_norsz13 a_6927_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2377 VPWR a_2387_13407 a_2374_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2378 tdc0.r_dly_store_ring2 a_15319_19355 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2379 a_24546_20327 _140_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X2381 a_14064_10205 _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2382 a_9374_20693 a_9206_20719 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2383 VPWR tdc1.w_ring_norsz30 a_29743_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2384 tdc1.w_dly_stop4 a_16311_10927 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2386 tdc1.r_dly_store_ctr13 a_19735_11989 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2389 VPWR a_6487_15003 a_6403_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2390 VPWR net38 a_29099_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2391 a_22905_13481 a_22358_13225 a_22558_13380 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2392 _094_ a_13735_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2393 tdc0.w_ring_norsz26 tdc0.w_ring_norsz10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R34 VPWR tdc0.g_ring317.stg01_46.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2395 VGND net17 tdc1.w_ring_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2397 a_17586_12335 tdc1.r_ring_ctr13 a_17417_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X2398 a_26521_14191 _170_ a_26439_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2399 tdc1.w_ring_norsz26 net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2400 VGND a_29055_15975 tdc1.r_dly_store_ring12 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2401 net36 a_28599_15797 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2402 tdc1.w_ring_buf3 a_20911_17455 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2403 VGND a_16219_11471 _625_.X VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2404 a_17041_12559 a_15851_12559 a_16932_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2405 tdc0.w_ring_buf16 a_5087_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2406 a_11237_17999 tdc0.w_ring_buf20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2408 a_30093_14197 a_29927_14197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2409 VPWR _076_ a_15801_19414 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X2410 VGND _197_ _038_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2412 VPWR a_17470_13759 a_17397_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2413 a_4069_13647 tdc0.r_ring_ctr11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2414 VPWR tdc1.w_ring_norsz1 a_18887_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2415 a_24467_16599 tdc1.r_dly_store_ctr10 a_24641_16705 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2418 a_19517_11471 tdc1.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2420 VGND a_23891_20719 a_24059_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2421 a_7201_10625 a_6983_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2422 VPWR a_13611_20327 _127_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X2423 VGND a_12507_10143 tdc0.r_ring_ctr0 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2424 VPWR tdc0.r_ring_ctr12 _163_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2426 a_19605_13423 tdc1.r_ring_ctr15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2427 a_16937_16367 a_16403_16373 a_16842_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2429 _026_ a_26439_14191 a_26689_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X2430 VPWR a_5694_17023 a_5621_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2431 a_9103_12247 tdc0.r_ring_ctr5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X2432 a_8565_16911 a_8399_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2433 a_28381_15279 a_28043_15511 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2436 tdc0.w_ring_norsz29 tdc0.w_ring_int_norsz29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2437 a_22297_18249 tdc1.w_ring_norsz25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2439 VGND a_21223_15101 a_21391_15003 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2440 VGND net29 a_11343_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2442 a_13948_16911 _112_ a_14032_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2444 VPWR net16 _061_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2445 VGND a_7166_19605 a_7124_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2446 VPWR a_12594_12671 a_12521_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2447 a_11875_9839 _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2448 VGND a_17567_10099 net16 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2449 _106_ a_21647_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2452 a_27342_19908 a_27135_19849 a_27518_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X2454 a_23063_14013 a_22365_13647 a_22806_13759 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2455 VGND tdc1.r_dly_store_ring12 a_23489_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2457 a_4420_11305 a_3505_10933 a_4073_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2458 a_9957_18249 tdc0.w_ring_norsz20 a_9873_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2460 a_5989_14197 a_5823_14197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2461 VGND tdc1.w_ring_int_norsz18 tdc1.w_ring_norsz18 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2462 VGND tdc1.r_ring_ctr10 a_21103_10633 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2463 tdc1.w_ring_norsz10 net15 a_22653_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2465 VGND a_21886_18517 a_21844_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2466 a_2396_15823 a_1481_15823 a_2049_16065 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2467 a_27271_20009 a_27135_19849 a_26851_19863 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2468 VGND a_9631_16189 a_9799_16091 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2469 tdc1.w_ring_int_norsz5 net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2471 a_18051_12015 tdc1.r_ring_ctr14 _189_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.27 ps=2.54 w=1 l=0.15
X2472 a_12897_17455 tdc0.r_dly_store_ctr15 a_12815_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2473 a_7393_15279 tdc0.w_ring_norsz27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2474 a_15259_16885 a_15550_17185 a_15501_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2475 tdc1.w_ring_buf1 a_18887_20719 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
R35 net47 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2476 a_10953_20175 a_9963_20175 a_10827_20541 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2478 VPWR a_2387_14495 tdc0.r_ring_ctr12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2479 a_7159_17076 tdc0.w_ring_norsz29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2480 a_7166_19605 a_6998_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2482 _084_ net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2483 _140_ a_24131_19337 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2484 tdc0.w_ring_buf7 a_11251_20719 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2485 a_10492_10383 a_9577_10383 a_10145_10625 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2488 VPWR net32 a_16162_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X2489 VGND a_10275_15101 a_10443_15003 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2490 a_21886_19605 a_21718_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2491 VGND a_29099_19631 net37 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2492 a_9025_12559 a_8859_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2493 VPWR tdc1.w_ring_buf16 a_25849_15657 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2494 a_22269_18921 a_21279_18549 a_22143_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2495 VGND a_23634_20693 a_23592_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2496 a_14172_20149 _143_ a_14560_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2497 a_7783_12925 a_7001_12559 a_7699_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2498 VGND _069_ a_12793_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2499 tdc0.r_dly_store_ring7 a_12559_21531 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2500 VPWR net8 a_8675_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2502 tdc0.w_ring_int_norsz27 tdc0.w_ring_norsz26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2504 a_16734_14165 a_16566_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2505 _118_ a_12079_16073 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2506 tdc0.w_ring_int_norsz25 net54 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2507 a_17043_16073 _076_ a_16825_15797 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2509 VPWR a_8912_21237 net27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2510 VPWR a_12332_10217 a_12507_10143 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2511 VGND tdc1.r_dly_store_ctr11 a_22569_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2512 a_6921_17455 tdc0.w_ring_norsz13 a_6837_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2513 a_17287_11471 a_16937_11471 a_17192_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2515 VPWR tdc1.w_ring_norsz31 a_27617_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2517 VPWR net25 a_12805_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2518 tdc0.r_dly_store_ring29 a_7591_16091 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2519 a_7676_18921 a_7277_18549 a_7550_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2522 VGND a_7350_20287 a_7308_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2524 VPWR _167_ a_29457_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2526 VGND a_8638_13077 a_8596_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2527 VGND a_15595_19605 a_15553_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2528 VPWR tdc0.w_ring_norsz29 a_6365_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2530 a_20273_19337 tdc1.w_ring_norsz8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2531 _059_ net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2532 a_24879_14569 a_24743_14409 a_24459_14423 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2533 VGND net16 a_18243_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2534 a_10804_15823 a_10405_15823 a_10678_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2535 a_21445_19637 a_21279_19637 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2536 a_11789_19087 tdc0.w_ring_buf5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2537 a_27003_12257 net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2538 VGND a_13330_13077 a_13288_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2539 a_13253_16687 tdc0.r_dly_store_ctr9 a_12907_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2540 VGND net31 a_10883_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2541 a_18072_15279 _196_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X2542 VGND tdc1.w_ring_int_norsz24 tdc1.w_ring_norsz24 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2544 a_30289_12559 a_29099_12559 a_30180_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2545 a_8895_13103 a_8197_13109 a_8638_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2546 VGND net30 a_16481_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2547 VGND net67 tdc1.w_ring_int_norsz20 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2548 tdc1.r_dly_store_ring9 a_22311_19605 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2552 a_14032_16911 _117_ a_13861_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2553 a_13897_15599 tdc0.r_dly_store_ring26 a_13551_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2554 VGND a_21131_17277 a_21299_17179 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2555 a_13587_13103 a_12889_13109 a_13330_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2557 tdc0.w_ring_norsz23 net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2558 tdc1.r_dly_store_ring9 a_22311_19605 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2559 VGND tdc1.w_ring_int_norsz23 tdc1.w_ring_norsz23 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2562 VGND _062_ a_16629_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2564 a_28239_11445 _048_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2565 a_11122_12671 a_10954_12925 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2566 VPWR a_27679_21237 net42 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2567 a_30534_15253 a_30366_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2568 _188_ a_17691_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X2569 a_13097_10927 tdc0.r_ring_ctr3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2570 _178_ a_22199_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
R36 net63 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2572 a_21791_20327 a_21934_20221 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X2573 VGND a_4687_13407 a_4621_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2574 VGND _076_ a_16353_20502 VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X2575 VPWR a_20131_20340 tdc1.w_ring_buf2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2576 VPWR a_27159_11989 a_27090_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X2577 VGND a_6855_14165 a_6813_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2578 a_2001_16911 a_1957_17153 a_1835_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2579 VPWR _196_ a_18072_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2580 VGND net41 tdc1.w_ring_int_norsz8 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2582 a_11966_21629 a_11693_21263 a_11881_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2583 a_24087_18775 a_24451_18864 a_24409_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2585 VGND net72 tdc1.w_ring_int_norsz25 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2586 a_3963_15101 a_3339_14735 a_3855_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2587 a_7607_20541 a_6743_20175 a_7350_20287 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2588 a_12402_10927 a_11325_10933 a_12240_11305 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2589 VGND net36 a_29927_15285 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2591 VGND net7 a_1131_14197 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2593 tdc0.r_ring_ctr13 a_4595_14709 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2594 a_14421_10205 a_14377_9813 a_14255_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2595 a_7277_20541 a_6743_20175 a_7182_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2597 a_3689_16373 a_3523_16373 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2598 a_11141_12021 a_10975_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2599 VPWR a_17804_15279 uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2601 a_11672_10205 _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2602 _087_ a_25221_19605 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2603 a_17121_17461 a_16955_17461 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2604 tdc0.w_ring_int_norsz7 net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2607 VGND net3 a_13183_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2609 a_5441_16911 tdc0.w_ring_buf17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2611 a_23542_17429 a_23374_17455 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2612 a_19889_19337 net14 tdc1.w_ring_norsz24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2614 a_29553_19337 tdc1.w_ring_norsz14 a_29469_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2617 VPWR a_20817_12801 a_20707_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2618 a_29642_20149 a_29442_20449 a_29791_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2619 VPWR tdc1.r_ring_ctr9 a_25623_11247 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X2620 a_27951_20951 a_28047_20951 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2621 a_6557_10901 a_6339_11305 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2622 a_22070_11583 a_21902_11837 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2623 a_11985_9813 a_11767_10217 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2624 a_23374_17455 a_23101_17461 a_23289_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2625 a_7285_16367 net22 tdc0.w_ring_norsz28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2627 VGND net30 a_15575_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2628 VGND _071_ a_13669_16705 VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2629 a_17217_9839 tdc1.r_ring_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2630 a_12341_12559 tdc0.r_ring_ctr0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2631 a_22343_15975 tdc1.r_dly_store_ctr1 a_22469_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2632 _076_ a_13735_21263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2633 tdc0.w_ring_buf5 a_10331_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2634 VGND net19 tdc0.w_ring_norsz31 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2635 a_5805_13647 a_5639_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2636 a_22741_16367 _087_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X2637 a_13161_18863 tdc0.r_dly_store_ring20 a_12723_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2638 a_27077_16367 tdc1.w_ring_int_norsz27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2639 VPWR a_11839_17277 a_12007_17179 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2641 VPWR tdc0.w_ring_norsz11 a_7847_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2642 a_17463_21085 a_17243_21097 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X2643 VGND a_26111_20938 tdc1.w_ring_buf16 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2645 a_19770_11583 a_19602_11837 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X2647 _041_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2648 tdc0.w_ring_int_norsz5 net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2651 VPWR tdc0.w_ring_norsz26 a_9227_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2652 a_7549_15823 a_6559_15823 a_7423_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2653 VGND a_5510_19199 a_5468_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2654 a_7161_12353 tdc0.r_ring_ctr7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2656 a_18030_20175 _090_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2657 a_21339_12533 a_21164_12559 a_21518_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2659 a_6796_17973 net23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
R37 uio_out[3] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2661 VGND tdc1.w_ring_norsz31 a_26983_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2662 a_23190_19631 a_22751_19637 a_23105_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2664 VGND net20 _042_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2665 a_25849_15657 a_25295_15497 a_25502_15556 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2666 a_15277_19087 a_14287_19087 a_15151_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2668 a_16055_19414 tdc1.r_dly_store_ring2 a_15983_19414 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2669 VGND a_24743_14409 a_24750_14313 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2670 a_25431_15657 a_25302_15401 a_25011_15511 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2671 VPWR tdc0.w_ring_norsz24 a_11159_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2672 VPWR tdc0.w_ring_norsz3 a_9585_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2673 VPWR a_30088_12393 a_30263_12319 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2674 a_19789_14191 a_19255_14197 a_19694_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2675 VGND a_9006_17023 a_8964_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2676 a_9263_17277 a_8399_16911 a_9006_17023 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2678 VGND a_4687_12319 a_4621_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2679 VGND a_25287_18517 _068_ VGND sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2681 VPWR net31 a_16127_18549 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2682 VPWR a_20195_11739 a_20111_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2683 a_17485_14735 tdc0.r_dly_store_ring8 a_17047_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2684 a_23799_17455 a_23101_17461 a_23542_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2685 _083_ a_16187_19891 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2686 a_23374_17455 a_22935_17461 a_23289_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2687 a_11322_15101 a_10883_14735 a_11237_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2688 a_5921_17455 tdc0.w_ring_norsz17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2689 a_4404_19061 net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2692 VPWR a_5951_17277 a_6119_17179 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
R38 VGND net45 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2693 a_17773_12559 tdc1.r_ring_ctr12 a_17691_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X2694 VPWR a_16991_18543 a_17159_18517 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2695 a_19685_21263 a_19131_21237 a_19338_21237 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X2696 VGND tdc0.r_ring_ctr0 _000_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2697 VGND _090_ a_18030_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R39 tdc1.g_ring326.stg01_73.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2698 a_17015_10383 a_16569_10383 a_16919_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2700 a_11448_17999 a_11049_17999 a_11322_18365 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2701 _092_ a_14366_15599 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X2702 VPWR _198_ _054_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2703 VGND a_26581_18145 _124_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X2704 VGND a_26819_15003 a_26777_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2705 tdc0.w_ring_norsz4 net21 a_9957_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2706 a_21623_11293 tdc1.r_ring_ctr10 a_21527_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X2707 a_13817_14191 tdc0.r_dly_store_ctr10 a_13735_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2708 a_7124_15823 a_6725_15823 a_6998_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2709 a_6607_11623 tdc0.r_ring_ctr6 a_6841_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2711 VGND _089_ a_17126_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2713 a_17065_20719 a_16727_20951 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X2714 VGND _065_ a_27705_17687 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X2715 a_5767_19453 a_4903_19087 a_5510_19199 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2717 a_21844_20009 a_21445_19637 a_21718_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2721 a_5894_15101 a_5621_14735 a_5809_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X2722 VPWR tdc0.r_ring_ctr8 _157_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2723 VGND _099_ a_17478_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2724 _135_ a_13583_19115 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2726 a_12332_10217 a_11251_9845 a_11985_9813 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2727 VGND _198_ _055_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2728 a_5437_19453 a_4903_19087 a_5342_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2729 VPWR a_30355_12533 a_30342_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2731 VGND tdc0.w_ring_buf0 a_9503_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2733 _183_ a_20819_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X2735 VPWR net30 a_15575_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2736 VPWR _087_ a_20175_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X2737 VPWR a_9799_16091 a_9715_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2738 a_17924_17063 _111_ a_18155_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2741 a_24879_14569 a_24750_14313 a_24459_14423 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2743 a_3295_19252 net27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2744 a_6018_11517 _156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X2745 a_17659_10357 _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2746 VPWR a_6319_15101 a_6487_15003 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2747 VPWR _072_ a_13583_19115 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2749 tdc1.w_ring_int_norsz26 net73 a_22297_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2752 a_9125_19631 net21 tdc0.w_ring_norsz6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2757 _626_.X a_2656_18517 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2759 _072_ _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2761 a_14917_19631 tdc1.w_ring_buf2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2762 a_24213_19337 tdc1.r_dly_store_ring23 a_24131_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2764 tdc0.w_ring_norsz10 tdc0.w_ring_norsz26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2767 a_9631_20719 a_8933_20725 a_9374_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2768 VPWR a_6027_16091 a_5943_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2769 _083_ a_16187_19891 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2770 a_9631_16189 a_8933_15823 a_9374_15935 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2771 a_12594_12671 a_12426_12925 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2773 a_7833_17455 tdc0.w_ring_buf12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2774 a_15451_20149 net24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2777 tdc1.r_dly_store_ring24 a_20287_14165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2779 VGND tdc1.r_ring_ctr11 a_21095_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X2780 tdc0.w_ring_buf14 a_6283_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2782 a_9025_12559 a_8859_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2783 a_14623_16627 _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2784 tdc0.r_ring_ctr5 a_9931_11445 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2785 VPWR a_9006_17023 a_8933_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2786 a_21633_19631 tdc1.w_ring_buf9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2787 tdc0.r_ring_ctr4 a_10667_10357 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2789 a_12517_21263 a_11527_21263 a_12391_21629 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2790 tdc1.r_dly_store_ring10 a_23323_19355 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2793 a_28905_14557 tdc1.r_ring_ctr1 a_28823_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X2794 tdc0.w_ring_int_norsz28 net57 a_7393_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2796 a_9287_11471 a_8841_11471 a_9191_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2797 VPWR _105_ a_22447_15395 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2798 uo_out[2] a_16656_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2799 a_15196_16073 _108_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X2801 VPWR net7 a_3431_13109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2802 VGND a_25971_17999 _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2803 a_4621_12393 a_3431_12021 a_4512_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2804 a_13277_15599 _071_ a_12867_15511 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X2805 a_26778_13235 a_27056_13219 a_27012_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2806 a_25551_17545 _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.157 ps=1.17 w=0.42 l=0.15
X2808 a_23485_9839 _179_ a_23403_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2809 a_21912_14511 tdc1.r_dly_store_ring8 a_21337_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X2810 a_9647_15253 net28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2811 a_5694_17023 a_5526_17277 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2812 a_27012_18249 _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X2813 a_18141_19337 net14 tdc1.w_ring_norsz22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2814 a_24719_15101 a_24021_14735 a_24462_14847 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2815 VPWR a_2049_16065 a_1939_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2817 a_15750_16885 a_15550_17185 a_15899_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X2818 a_27307_14887 a_27403_14709 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2819 VPWR net16 _058_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2820 a_29615_12559 a_29265_12559 a_29520_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2821 VGND a_15262_13759 a_15220_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2822 VPWR a_23055_15975 _110_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X2823 _625_.X a_16219_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2824 a_16589_15823 _069_ a_16155_15975 VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2826 a_14265_15823 tdc0.r_dly_store_ring11 a_13827_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2827 net13 a_5087_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2829 a_10359_15101 a_9577_14735 a_10275_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2830 VGND a_14799_11445 net29 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2831 VGND a_4130_16341 a_4088_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2833 a_2623_12335 _157_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2834 tdc1.w_ring_int_norsz9 net41 a_20273_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2835 VGND _197_ _037_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2837 tdc1.w_ring_norsz16 tdc1.w_ring_int_norsz16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2838 VPWR _162_ a_1113_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2839 _624_.X a_15904_11445 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2840 VPWR net25 a_12897_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2841 a_28047_21237 net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2843 VGND a_7442_12671 a_7400_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2845 a_27159_11989 a_26964_12131 a_27469_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X2846 VGND a_19355_13103 _022_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X2847 VPWR net27 a_7479_17461 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2848 VPWR tdc1.r_ring_ctr0 _016_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2850 a_6913_15823 tdc0.w_ring_buf29 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2851 a_13809_9845 a_13643_9845 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2852 VGND a_17567_10099 net16 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2853 a_15603_14013 a_14821_13647 a_15519_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2855 uo_out[6] a_13344_20693 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2856 a_17027_10749 _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2857 tdc0.r_dly_store_ring26 a_11915_15003 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2859 VGND tdc0.w_ring_norsz0 tdc0.w_ring_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2860 a_22067_13335 a_22358_13225 a_22309_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2861 a_6445_14735 a_5455_14735 a_6319_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2864 _061_ net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2867 a_12240_11305 a_11325_10933 a_11893_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2868 VPWR a_28078_16885 a_28007_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X2870 VPWR a_2479_16885 a_2466_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2871 VPWR tdc1.w_ring_norsz5 a_18233_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2872 a_10402_20541 a_9963_20175 a_10317_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2874 a_7079_11231 a_6904_11305 a_7258_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2875 a_12805_17161 tdc0.r_dly_store_ctr4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2877 _148_ _145_ a_13097_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
R40 VPWR tdc1.g_ring322.stg01_69.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2879 a_14032_16911 _117_ a_14300_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2880 net10 a_26615_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2881 VGND a_2479_16885 a_2413_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2882 VGND a_6987_12247 _154_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2883 VPWR net10 a_29099_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2884 VPWR a_9839_17715 net39 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2885 VPWR a_30263_12319 tdc1.r_ring_ctr1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2886 VGND a_12007_17179 a_11965_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2887 tdc0.r_dly_store_ring14 a_7775_20443 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2888 a_26747_18863 a_26431_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2891 a_26851_19863 a_27142_19753 a_27093_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2893 VGND _127_ a_12618_21039 VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.185 ps=1.22 w=0.65 l=0.15
X2895 tdc1.w_ring_norsz13 tdc1.w_ring_int_norsz13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2897 VPWR a_22603_21629 a_22771_21531 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2899 VGND a_13019_12827 a_12977_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2901 tdc0.w_ring_norsz13 net22 a_7289_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2903 VPWR a_25203_10357 a_25190_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2904 _180_ _179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2905 VPWR a_23323_19355 a_23239_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2906 a_30791_16367 a_29927_16373 a_30534_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2907 net37 a_29099_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2908 VPWR a_22070_11583 a_21997_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2909 a_24736_13647 _027_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2910 a_29185_19337 tdc1.w_ring_norsz30 a_29101_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2911 VGND _033_ a_14421_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2912 VPWR net7 a_3431_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2914 a_5161_15823 a_4995_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2915 a_14560_20425 _143_ a_14172_20149 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2916 a_7699_12925 a_6835_12559 a_7442_12671 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2917 a_15196_16073 _108_ a_15027_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X2918 _197_ a_5087_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2919 a_30461_16367 a_29927_16373 a_30366_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2921 tdc0.r_dly_store_ring2 a_15319_19355 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2922 a_9301_20719 a_8767_20725 a_9206_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2923 tdc1.r_ring_ctr12 a_17659_10357 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X2924 a_17287_11471 a_16771_11471 a_17192_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2925 a_18383_17076 tdc1.w_ring_norsz20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2926 a_21844_12393 a_21445_12021 a_21718_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2927 a_5805_13647 a_5639_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2928 a_7369_12925 a_6835_12559 a_7274_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2930 VPWR a_19770_11583 a_19697_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2933 a_23403_9839 _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2934 VGND a_6119_17179 a_6077_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2936 VPWR a_29741_11989 a_29631_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2937 VPWR net16 _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2938 VPWR a_18731_17063 _133_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X2939 tdc1.r_dly_store_ctr8 a_20195_11739 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2941 tdc0.w_dly_stop5 a_3707_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2942 a_17309_17455 tdc1.w_ring_buf22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2943 VGND a_4595_14709 a_4529_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2944 a_13641_9545 tdc0.r_ring_ctr0 a_13559_9545 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2945 a_13905_17999 tdc0.w_ring_buf4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2946 a_7465_18543 tdc0.w_ring_buf13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X2948 tdc1.r_dly_store_ctr9 a_22495_11739 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2949 VPWR a_15170_11989 a_15097_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X2950 a_30434_14013 a_29357_13647 a_30272_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2951 a_13993_16073 tdc0.r_dly_store_ring3 a_13909_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2952 VGND a_5087_11471 _197_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2953 a_26667_21237 ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2954 tdc1.w_ring_int_norsz20 tdc1.w_ring_norsz19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2955 tdc0.w_ring_buf14 a_6283_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2956 a_2953_11247 tdc0.r_ring_ctr8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2957 a_18961_10383 a_18795_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2959 a_16991_14191 a_16127_14197 a_16734_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2960 a_6244_11293 _013_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2961 a_24831_13647 a_24315_13647 a_24736_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2962 a_17010_16341 a_16842_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X2964 a_17243_21097 a_17114_20841 a_16823_20951 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X2966 a_19743_16367 a_18961_16373 a_19659_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2967 VGND net70 tdc1.w_ring_int_norsz23 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2968 net2 a_29559_21263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2969 tdc1.w_ring_norsz23 tdc1.w_ring_norsz7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2971 VGND _166_ _005_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2972 VPWR _116_ a_13861_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X2973 a_16661_14191 a_16127_14197 a_16566_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2975 net42 a_27679_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2976 a_23891_20719 a_23027_20725 a_23634_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2977 VPWR net28 a_6559_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2979 a_9121_15823 tdc0.w_ring_buf21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2980 VPWR _065_ a_26426_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X2982 a_27622_14735 a_27307_14887 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X2985 VGND tdc1.w_ring_int_norsz12 tdc1.w_ring_norsz12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2986 VGND a_24738_15935 a_24696_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X2987 a_24995_16189 a_24131_15823 a_24738_15935 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X2989 VPWR tdc1.w_ring_buf15 a_28885_21097 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X2990 VPWR _160_ _161_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2991 a_28977_15657 a_28430_15401 a_28630_15556 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X2992 a_23561_20719 a_23027_20725 a_23466_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X2993 VGND a_15196_16073 uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2994 tdc1.w_ring_int_norsz8 tdc1.w_ring_norsz7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2995 a_5859_16189 a_5161_15823 a_5602_15935 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2996 a_5434_16189 a_4995_15823 a_5349_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2997 a_15719_21237 net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2999 a_17804_15279 _192_ a_17720_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3000 VGND tdc0.w_ring_norsz13 a_6927_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3001 tdc1.w_ring_int_norsz25 tdc1.w_ring_norsz24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3003 VGND a_14172_20149 uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X3004 a_24665_16189 a_24131_15823 a_24570_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3005 tdc0.w_ring_int_norsz18 net47 a_5921_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3006 a_27017_19337 _067_ a_26933_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3007 a_4165_11989 a_3947_12393 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3008 a_15553_20009 a_14563_19637 a_15427_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3009 VGND tdc1.w_ring_norsz30 a_29743_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3010 VPWR a_28630_15556 a_28559_15657 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3014 a_8010_14191 a_7571_14197 a_7925_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3015 _056_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3018 VPWR a_30534_16341 a_30461_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3019 a_30549_17999 a_29559_17999 a_30423_18365 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3020 VPWR a_9374_20693 a_9301_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3022 VGND net29 a_10975_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3023 a_24477_19087 tdc1.r_dly_store_ring31 a_24131_19337 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3024 net13 a_5087_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3025 tdc0.r_dly_store_ring15 a_5935_19355 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3026 tdc1.r_dly_store_ring20 a_17435_16341 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3027 a_18939_20327 _084_ a_19267_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3028 a_17094_12925 a_16017_12559 a_16932_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3029 VGND net20 _045_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3030 a_27518_16189 a_27271_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3031 VPWR _082_ a_22256_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X3033 VGND a_9466_12671 a_9424_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3034 a_9677_19337 net50 tdc0.w_ring_int_norsz21 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3036 VGND a_2571_15797 a_2505_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3037 tdc1.r_dly_store_ring17 a_22771_21531 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3038 VGND tdc1.w_ring_int_norsz0 tdc1.w_ring_norsz0 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3039 VPWR net27 a_7111_18549 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3040 VPWR tdc0.w_ring_norsz3 a_10147_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3041 VPWR _026_ a_27814_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3043 VGND tdc0.w_ring_norsz9 tdc0.w_ring_int_norsz10 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3044 a_29469_19337 tdc1.w_ring_int_norsz30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3046 tdc0.r_dly_store_ctr4 a_11547_12827 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3047 tdc0.r_dly_store_ring7 a_12559_21531 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3049 VGND tdc1.w_ring_norsz6 tdc1.w_ring_int_norsz7 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3050 VGND a_24915_15511 tdc1.r_dly_store_ring16 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3051 VPWR a_14623_16627 _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3052 a_4404_19061 net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3053 VPWR a_7975_18543 a_8143_18517 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3055 a_10405_15823 a_10239_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3056 tdc1.w_ring_buf3 a_20911_17455 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3059 a_20819_11471 tdc1.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X3060 VGND _038_ a_7245_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3061 a_3788_15599 tdc0.r_ring_ctr12 a_3485_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X3062 a_25103_16599 _084_ a_25431_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3063 VGND a_7975_18543 a_8143_18517 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3064 a_22615_16599 tdc1.r_dly_store_ring3 a_22855_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X3065 a_13669_16705 tdc0.r_dly_store_ctr12 a_13583_16705 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X3066 a_29427_20693 net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X3067 a_21886_11989 a_21718_12015 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3068 a_20713_14735 tdc1.w_ring_buf8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3069 VPWR _185_ a_17691_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X3070 VPWR a_16734_14165 a_16661_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3071 a_30124_17999 a_29725_17999 a_29998_18365 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3074 a_11877_19631 a_11343_19637 a_11782_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3076 tdc1.r_dly_store_ctr15 a_23231_13915 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3077 VGND a_26031_16885 net41 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3078 a_4512_12393 a_3597_12021 a_4165_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3079 _194_ a_20911_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X3080 VGND a_12375_13915 a_12333_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3081 VPWR a_15427_20719 a_15595_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3082 a_16569_10383 a_16403_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3083 a_9723_12925 a_8859_12559 a_9466_12671 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3084 VPWR a_23634_20693 a_23561_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3085 VGND tdc0.w_ring_int_norsz8 tdc0.w_ring_norsz8 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3086 VPWR _079_ a_13817_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3087 a_17129_14985 _089_ a_17213_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3089 a_19567_12015 a_18869_12021 a_19310_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3090 tdc0.w_ring_buf30 a_6651_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3091 _057_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3093 VPWR a_27894_14709 a_27823_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3094 VPWR a_24738_15935 a_24665_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3095 a_11325_10933 a_11159_10933 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3096 VGND a_22995_10357 a_22929_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3097 a_9393_12925 a_8859_12559 a_9298_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3098 VGND a_17208_20149 uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3099 a_17027_10749 a_16403_10383 a_16919_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3100 _068_ a_25287_18517 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3101 a_19694_14191 a_19255_14197 a_19609_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3102 a_24927_13647 a_24481_13647 a_24831_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3103 a_5434_16189 a_5161_15823 a_5349_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3104 tdc1.w_ring_norsz16 net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3108 a_22178_21629 a_21905_21263 a_22093_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3110 a_16734_18517 a_16566_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3111 a_1297_14197 a_1131_14197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3112 a_7737_14197 a_7571_14197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3113 VGND tdc0.r_dly_store_ctr14 a_13277_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X3114 a_18030_20175 _078_ a_17208_20149 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3115 tdc1.r_dly_store_ctr11 a_22311_11989 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3116 VGND tdc0.w_ring_norsz5 tdc0.w_ring_norsz21 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3117 VPWR tdc0.r_ring_ctr0 a_13551_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X3118 a_25111_20327 net24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X3120 a_21905_16911 a_21739_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3121 a_17208_20149 _091_ a_17678_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3122 tdc0.w_dly_stop5 a_3707_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3123 a_25295_15497 net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3124 tdc1.r_dly_store_ctr11 a_22311_11989 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3125 VGND a_16656_16885 uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3128 a_13615_17571 _114_ a_13543_17571 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3130 VGND _152_ a_6244_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3131 a_8562_15279 a_8123_15285 a_8477_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3134 a_24777_20425 _139_ a_24681_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3135 a_27135_19849 net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3136 a_9004_20149 net22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3138 VGND a_17903_16599 _111_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3139 a_17478_16911 _095_ a_16656_16885 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3140 a_10654_10749 a_9577_10383 a_10492_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3142 a_17673_13109 a_17507_13109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3143 a_18383_17076 tdc1.w_ring_norsz20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3145 a_15027_15823 _103_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3146 a_14555_10901 a_14399_11169 a_14700_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X3147 VGND a_3946_15935 a_3904_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3148 a_3786_14191 _163_ a_3483_14423 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3149 a_12415_11231 a_12240_11305 a_12594_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3150 tdc0.w_ring_norsz24 net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3152 VGND net21 tdc0.w_ring_norsz19 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3153 VGND net3 _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3155 a_27761_11471 a_27717_11713 a_27595_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3157 a_29357_13647 a_29191_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3159 a_10873_13897 net23 tdc0.w_ring_norsz9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3160 _076_ a_13735_21263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3161 VGND net10 a_29099_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3162 a_3873_16189 a_3339_15823 a_3778_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3163 VGND a_11915_18267 a_11873_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3164 VGND a_6246_13759 a_6204_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3165 a_13583_19115 tdc0.r_dly_store_ring23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X3166 a_20621_16911 tdc1.w_ring_buf19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3167 a_19685_21263 a_19138_21537 a_19338_21237 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3168 a_24694_11517 _179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X3169 a_24030_13647 _170_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X3170 VGND a_29642_20149 a_29571_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
R41 VGND net51 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3171 VPWR a_21327_10071 _181_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X3173 VGND a_14623_16627 _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
R42 tdc0.g_ring326.stg01_55.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3175 a_22855_16687 _086_ a_22748_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3176 a_24021_14735 a_23855_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3177 VPWR a_15196_16073 uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3178 VGND a_20195_11739 a_20153_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3179 VPWR a_9466_12671 a_9393_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3180 VPWR a_23967_17429 a_23883_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3181 VGND a_20131_20340 tdc1.w_ring_buf2 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3182 tdc1.w_ring_int_norsz19 net66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3183 a_9299_11837 a_8675_11471 a_9191_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3184 VGND a_20119_14191 a_20287_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3185 VPWR tdc0.r_ring_ctr12 a_945_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3188 VPWR _034_ a_14700_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X3189 VPWR tdc0.r_ring_ctr2 a_13603_11445 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X3190 VPWR net26 a_6559_13109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3191 VGND a_13879_10901 tdc0.r_ring_ctr2 VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3192 a_30366_14191 a_29927_14197 a_30281_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3193 a_1485_12809 tdc0.r_ring_ctr10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3194 VPWR a_4404_19061 net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3195 VGND a_28239_11445 tdc1.r_ring_ctr0 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3196 VPWR a_7423_13103 a_7591_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3197 VPWR tdc1.w_ring_norsz7 a_16679_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3200 a_15553_12393 a_14563_12021 a_15427_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3201 a_29473_17455 tdc1.w_ring_norsz28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3202 VGND net35 a_22935_17461 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3203 a_11049_17999 a_10883_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3204 VGND net16 _058_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3205 VGND a_7423_13103 a_7591_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3206 a_19237_18249 tdc1.w_ring_norsz21 a_19153_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3209 tdc0.r_dly_store_ctr7 a_7867_12827 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3210 a_11697_13647 tdc0.w_ring_buf24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3212 a_12793_14511 tdc0.r_dly_store_ring24 a_12447_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3213 _064_ a_25971_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X3214 a_18337_16687 _083_ a_17903_16599 VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3215 a_28814_13423 tdc1.r_ring_ctr0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X3216 tdc1.w_ring_buf7 a_16679_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3217 VGND _141_ a_24546_20327 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X3218 VPWR a_29791_20938 tdc1.w_ring_buf15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3219 a_27587_16885 a_27878_17185 a_27829_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X3220 a_17393_16745 a_16403_16373 a_17267_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3223 VGND _150_ _153_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3224 VGND tdc1.w_ring_norsz23 tdc1.w_ring_int_norsz24 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3225 _007_ tdc0.r_ring_ctr0 a_13809_9295 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X3226 a_24920_11471 tdc1.r_ring_ctr7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3227 VPWR a_21463_15823 _089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3228 VGND tdc1.w_ring_buf1 a_19685_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X3229 a_27003_11169 net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3230 VPWR a_1865_14165 a_1755_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3231 a_28358_15645 a_28043_15511 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3232 VGND a_27307_14887 tdc1.r_dly_store_ctr0 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3234 a_22730_19453 a_22457_19087 a_22645_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3235 a_13955_12015 a_13091_12021 a_13698_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3237 _192_ a_17047_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X3239 a_9004_20149 net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3240 VGND net39 tdc0.w_ring_int_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3241 a_29393_16189 a_29055_15975 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3242 a_11580_11293 _009_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3244 a_9756_11471 a_8675_11471 a_9409_11713 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3245 tdc1.r_ring_ctr7 a_25571_12319 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3247 _000_ tdc0.r_ring_ctr0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3249 a_8493_14985 tdc0.w_ring_int_norsz27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R43 uio_oe[6] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3250 a_15983_19414 a_15801_19414 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3251 VPWR tdc1.r_ring_ctr2 a_28455_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X3252 _069_ a_14623_16627 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3254 VGND _028_ a_27722_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3255 net29 a_14799_11445 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3256 VPWR net20 _043_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3257 VPWR a_3946_15935 a_3873_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3258 net12 a_5455_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3259 _037_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3260 VGND _163_ a_3701_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X3262 VPWR tdc1.w_ring_int_norsz22 a_18225_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3263 a_29055_15975 a_29151_15797 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3269 VGND _052_ a_26813_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X3270 a_27403_17973 _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X3271 a_17661_21097 a_17114_20841 a_17314_20996 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3272 a_17137_10625 a_16919_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
R44 VPWR tt_um_hpretl_tt06_tdc_v2_83.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3274 a_19517_11471 tdc1.r_ring_ctr8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3275 a_23075_18762 tdc1.w_ring_norsz10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3278 a_15519_14013 a_14655_13647 a_15262_13759 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3279 VPWR a_13344_20693 uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3280 a_23101_10933 a_22935_10933 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3281 VPWR net16 a_18243_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3282 VGND tdc0.w_ring_norsz11 a_7847_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3283 a_14415_18365 a_13717_17999 a_14158_18111 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3287 VPWR a_17314_20996 a_17243_21097 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3288 a_11103_16189 a_10239_15823 a_10846_15935 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3289 a_2466_17277 a_1389_16911 a_2304_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3291 a_21817_11471 tdc1.r_ring_ctr9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3294 a_13173_14511 tdc0.r_dly_store_ctr11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3295 a_15189_14013 a_14655_13647 a_15094_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3296 a_24021_14735 a_23855_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3297 a_7350_20287 a_7182_20541 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3298 a_9374_15935 a_9206_16189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3300 a_12907_16367 _072_ a_12989_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3301 VPWR a_18939_20327 _132_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X3303 tdc1.w_ring_buf16 a_25787_20719 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3304 a_8178_14165 a_8010_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3305 a_15262_13759 a_15094_14013 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3307 a_11540_16911 a_11141_16911 a_11414_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3308 a_16293_18549 a_16127_18549 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3311 a_17029_13647 a_16863_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3312 VGND net45 tdc0.w_ring_int_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3314 a_22603_21629 a_21905_21263 a_22346_21375 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3315 a_9309_19337 net40 tdc0.w_ring_int_norsz6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3316 VPWR a_14377_9813 a_14267_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3317 a_13551_15279 _075_ a_13633_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3318 net9 a_25932_12533 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3319 a_7289_17455 tdc0.w_ring_norsz29 a_7205_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3322 VGND _197_ _033_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3323 a_12552_12559 a_12153_12559 a_12426_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3324 VGND net28 a_6559_19637 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3326 tdc1.w_ring_norsz8 net14 a_19617_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3327 VGND net16 _062_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3328 a_24831_12393 a_24481_12021 a_24736_12381 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3331 _120_ a_13459_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X3332 a_19329_11471 a_19163_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3333 a_8497_11721 _150_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3334 a_11505_12559 a_10515_12559 a_11379_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3335 tdc1.r_ring_ctr5 a_25571_13621 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3336 VPWR net26 a_4995_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3338 tdc1.r_dly_store_ring10 a_23323_19355 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3340 a_14555_10901 a_14360_11043 a_14865_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
R45 VGND net57 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3342 VGND net20 a_5087_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3343 a_14917_12015 tdc0.r_ring_ctr1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3345 a_12618_21039 _130_ a_12864_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=2.77 as=0.125 ps=1.25 w=1 l=0.15
X3346 VPWR tdc0.w_ring_norsz20 a_9677_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3347 a_3947_13481 a_3597_13109 a_3852_13469 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3348 VPWR a_15151_19453 a_15319_19355 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3350 VPWR _142_ a_14560_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X3351 tdc1.w_ring_buf23 a_21923_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3352 VPWR a_27346_17687 _123_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X3354 tdc1.w_ring_norsz25 tdc1.w_ring_int_norsz25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3356 a_6461_18543 tdc0.w_ring_norsz14 a_6377_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3357 a_26627_18543 _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X3358 VPWR tdc0.w_ring_norsz31 a_6007_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3359 a_9850_15101 a_9577_14735 a_9765_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3360 VGND a_20051_10357 a_19985_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3362 tdc0.w_ring_int_norsz17 net46 a_4357_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3363 VPWR _198_ _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3364 VGND tdc0.w_ring_int_norsz15 tdc0.w_ring_norsz15 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3365 a_4209_13469 a_4165_13077 a_4043_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3367 VGND a_28915_10927 _198_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3369 _125_ a_20258_16073 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X3370 a_5652_16911 a_5253_16911 a_5526_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3371 _039_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3373 VGND a_8178_14165 a_8136_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3374 a_12494_9839 a_11417_9845 a_12332_10217 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3375 a_23615_19631 a_22917_19637 a_23358_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3376 a_23189_13647 a_22199_13647 a_23063_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3379 tdc0.r_dly_store_ctr15 a_4279_17179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3381 VGND _034_ a_14117_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X3382 VPWR a_19860_15797 _080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3383 VGND a_22346_17023 a_22304_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3384 a_22603_17277 a_21739_16911 a_22346_17023 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3385 a_24385_18249 a_24635_17973 _072_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3386 a_8385_13103 tdc0.r_ring_ctr9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3387 a_13909_16073 _076_ a_13827_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3388 a_8343_17455 a_7645_17461 a_8086_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3389 a_1551_15253 tdc0.r_ring_ctr12 a_1949_15645 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X3391 tdc0.w_ring_norsz18 net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3392 VGND net39 tdc0.w_ring_int_norsz15 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3393 a_11881_21263 tdc0.w_ring_buf7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3395 VGND tdc0.r_ring_ctr8 a_2703_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3396 VGND a_30355_12533 a_30289_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3397 VPWR net9 a_18795_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3399 a_13077_13103 tdc0.r_ring_ctr2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3400 a_22273_17277 a_21739_16911 a_22178_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3401 a_11839_12015 a_11141_12021 a_11582_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3402 VPWR tdc0.r_ring_ctr15 a_1129_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3403 VGND a_10287_20938 tdc0.w_ring_buf22 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3404 a_19659_16367 a_18795_16373 a_19402_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3405 a_3962_16367 a_3523_16373 a_3877_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3408 a_11414_12015 a_10975_12021 a_11329_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3409 VGND tdc1.w_ring_norsz7 a_16679_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3410 a_12889_16073 tdc0.r_dly_store_ctr5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3411 a_6998_19631 a_6725_19637 a_6913_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3412 VPWR _198_ _048_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3413 VGND a_18114_13077 a_18072_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3415 a_1736_15823 _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3416 a_29631_12015 _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3417 a_12507_10143 a_12332_10217 a_12686_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3418 a_10287_20938 tdc0.w_ring_norsz22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3419 a_28829_18543 tdc1.w_ring_norsz29 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3420 tdc0.r_ring_ctr7 a_7079_11231 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3421 a_22453_11471 a_21463_11471 a_22327_11837 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3422 a_16991_14191 a_16293_14197 a_16734_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3423 VGND a_17468_15797 _079_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X3424 tdc1.w_ring_buf7 a_16679_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3425 a_21223_15101 a_20525_14735 a_20966_14847 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3426 VPWR _185_ a_18051_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3427 a_6262_14191 a_5823_14197 a_6177_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3428 VPWR _089_ a_12448_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
X3429 VGND _198_ _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3430 VPWR tdc1.w_ring_norsz8 a_20083_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3431 VPWR _067_ a_25643_18775 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3432 a_18371_13103 a_17673_13109 a_18114_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3433 VPWR net30 a_14655_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3434 a_17117_14569 a_16127_14197 a_16991_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3435 _078_ a_15577_16483 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3436 tdc1.r_dly_store_ring30 a_30683_17429 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3437 VPWR a_9963_19631 net40 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3438 VGND _076_ a_14366_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X3439 a_29817_17461 a_29651_17461 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3440 _198_ a_28915_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3441 VPWR a_20316_18151 _126_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X3442 a_7723_10357 a_7548_10383 a_7902_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3443 a_26920_12015 a_26483_11989 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3444 tdc1.r_dly_store_ring30 a_30683_17429 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3445 a_28418_11471 _048_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3446 a_25317_13103 _174_ _027_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3447 a_18114_13077 a_17946_13103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3451 VPWR tdc0.w_ring_int_norsz9 a_10957_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3452 VPWR tdc0.r_ring_ctr0 a_13323_11159 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X3453 a_26755_19863 a_26851_19863 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3454 a_5510_19199 a_5342_19453 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3455 VPWR a_25203_10357 tdc1.r_ring_ctr8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3456 a_29631_12015 a_29007_12021 a_29523_12393 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3457 VGND a_5767_19453 a_5935_19355 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3458 a_25396_12393 a_24315_12021 a_25049_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3459 VGND tdc0.w_ring_norsz19 tdc0.w_ring_int_norsz20 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3460 a_10275_15101 a_9577_14735 a_10018_14847 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3461 a_1137_16073 _165_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3462 a_22346_21375 a_22178_21629 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3463 a_13361_19951 tdc0.r_dly_store_ring15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X3464 a_29357_13647 a_29191_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3466 a_24849_20425 _140_ a_24777_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3467 a_20038_10749 a_18961_10383 a_19876_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3468 a_4512_13481 a_3431_13109 a_4165_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3469 tdc1.w_ring_norsz0 tdc1.w_ring_norsz16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3470 VPWR tdc0.w_ring_norsz4 a_10137_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3471 tdc0.w_ring_int_norsz10 net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3472 a_30791_15279 a_30093_15285 a_30534_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3473 a_1552_13469 _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3474 VGND a_11379_12925 a_11547_12827 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3475 VPWR a_12391_21629 a_12559_21531 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3476 a_23075_18762 tdc1.w_ring_norsz10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3477 tdc1.w_ring_int_norsz7 net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3481 VPWR net34 a_22291_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3482 tdc1.w_ring_buf29 a_30295_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3483 VGND tdc1.w_ring_int_norsz4 tdc1.w_ring_norsz4 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3484 VPWR a_23615_19631 a_23783_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3485 a_4209_12381 a_4165_11989 a_4043_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3486 a_4043_13481 a_3597_13109 a_3947_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3487 net20 a_4443_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3490 VPWR net9 a_16771_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3491 a_25431_16367 tdc1.r_dly_store_ring26 a_25229_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3492 VGND a_28239_11445 a_28173_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3493 VGND a_23615_19631 a_23783_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3494 VPWR a_22346_17023 a_22273_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R46 VPWR tdc0.g_ring318.stg01_47.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3495 a_15118_10927 a_14399_11169 a_14555_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3496 a_30599_17455 a_29817_17461 a_30515_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3497 VGND _048_ a_27761_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3498 VPWR tdc1.r_ring_ctr13 a_17691_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3499 VGND net41 tdc1.w_ring_int_norsz2 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3500 a_7745_10927 _153_ _012_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3501 VPWR a_21299_17179 a_21215_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3502 a_28885_21097 a_28331_20937 a_28538_20996 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3503 a_25932_12533 tdc1.w_ring_buf0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3504 a_24209_14735 tdc1.r_ring_ctr7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3506 VGND _087_ a_21397_15617 VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3508 VGND a_15427_20719 a_15595_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3509 VGND net15 tdc1.w_ring_norsz2 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3510 VGND a_8730_15253 a_8688_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3511 VPWR net37 a_29651_17461 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3512 a_13990_18365 a_13551_17999 a_13905_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
R47 tdc0.g_ring331.stg01_60.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3513 VPWR _064_ a_24635_17973 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3514 a_22806_13759 a_22638_14013 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3515 VGND tdc0.w_ring_int_norsz2 tdc0.w_ring_norsz2 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3517 tdc1.w_ring_norsz28 tdc1.w_ring_norsz12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3520 VPWR _198_ _053_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3521 _063_ net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3523 _035_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3527 a_29105_17455 tdc1.w_ring_norsz12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3528 a_11923_12015 a_11141_12021 a_11839_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3529 VGND _172_ a_24745_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3530 a_11908_13647 a_11509_13647 a_11782_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3534 a_24831_12393 a_24315_12021 a_24736_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3535 a_9466_12671 a_9298_12925 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3536 a_21131_17277 a_20433_16911 a_20874_17023 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3537 VPWR a_18243_17999 net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3538 a_21886_18517 a_21718_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3539 a_5989_14197 a_5823_14197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3541 VPWR tdc1.w_ring_buf12 a_29989_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3544 VPWR tdc1.w_ring_norsz19 a_19991_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3545 a_7918_17455 a_7645_17461 a_7833_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3546 tdc1.w_ring_norsz9 net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3548 VPWR a_25396_12393 a_25571_12319 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3549 VPWR a_30272_13647 a_30447_13621 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3550 tdc1.r_dly_store_ring28 a_30959_16341 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3551 a_28253_20425 tdc1.w_ring_norsz15 a_28169_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3552 a_17852_11471 a_16771_11471 a_17505_11713 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3553 VGND a_25502_15556 a_25431_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3554 VPWR a_26297_20340 tdc1.w_ring_buf0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3555 a_3947_13481 a_3431_13109 a_3852_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3556 tdc1.r_dly_store_ring28 a_30959_16341 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3557 VGND _075_ a_17485_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X3558 VGND net5 a_25251_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3559 VGND a_22327_11837 a_22495_11739 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3560 tdc1.w_ring_int_norsz29 net76 a_29473_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3561 a_18869_14985 tdc1.r_dly_store_ctr6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3562 a_14557_14735 tdc0.r_dly_store_ring19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X3563 VPWR tdc1.w_ring_buf27 a_27689_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X3564 a_24641_16705 _071_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X3565 a_22615_16599 _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X3566 a_23615_19631 a_22751_19637 a_23358_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3568 VPWR a_22351_13321 a_22358_13225 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3569 VPWR a_11985_9813 a_11875_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3570 a_25230_15645 a_24915_15511 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3571 a_19751_15279 a_18887_15285 a_19494_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3572 VPWR a_19338_21237 a_19267_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3573 a_25251_19951 net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X3574 a_16155_15975 tdc0.r_dly_store_ctr1 a_16301_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X3575 a_17678_20175 _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X3576 VPWR a_25295_15497 a_25302_15401 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3577 a_27689_15823 a_27135_15797 a_27342_15797 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3579 uo_out[2] a_16656_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3580 VPWR a_17659_10357 tdc1.r_ring_ctr12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3583 a_27271_15823 a_27142_16097 a_26851_15797 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X3584 a_23285_19631 a_22751_19637 a_23190_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3585 a_12153_12559 a_11987_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3586 a_30129_18543 a_29791_18775 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X3587 VGND a_30534_14165 a_30492_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3588 a_25028_10383 a_24113_10383 a_24681_10625 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3589 VGND tdc0.w_ring_norsz17 tdc0.w_ring_norsz1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3590 VPWR tdc1.r_ring_ctr8 a_21331_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X3591 VGND a_25111_20327 _139_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3592 a_16293_14197 a_16127_14197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3596 a_14032_16911 _112_ a_13948_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3597 VGND net33 a_17507_13109 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3598 tdc0.r_dly_store_ctr13 a_6027_16091 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3600 VGND _075_ a_21912_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X3601 a_10827_20541 a_10129_20175 a_10570_20287 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3602 a_12993_15599 _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X3603 a_27159_10901 a_27003_11169 a_27304_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X3604 a_12161_16073 tdc0.r_dly_store_ctr13 a_12079_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3605 VPWR tdc1.r_dly_store_ctr10 a_24467_16599 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3606 a_22199_12559 _172_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3607 VPWR tdc0.r_ring_ctr14 a_1551_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
R48 VGND net67 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3610 tdc0.r_dly_store_ring8 a_17159_14165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3611 a_16097_16911 a_15543_16885 a_15750_16885 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X3612 a_20861_12559 a_20817_12801 a_20695_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
R49 VPWR tdc0.g_ring327.stg01_56.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3613 tdc1.r_dly_store_ring17 a_22771_21531 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3614 tdc1.w_dly_stop2 a_15575_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3615 a_1113_13647 tdc0.r_ring_ctr12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3617 a_29815_14013 a_29191_13647 a_29707_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3618 a_16932_12559 a_16017_12559 a_16585_12801 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3619 VGND _197_ _040_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3620 tdc1.w_ring_norsz18 tdc1.w_ring_norsz2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3621 tdc0.r_dly_store_ctr4 a_11547_12827 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3623 a_24368_10383 _030_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3624 a_8933_17277 a_8399_16911 a_8838_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3627 VPWR a_23231_13915 a_23147_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3628 a_11329_15279 tdc0.w_ring_buf19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3629 tdc1.r_dly_store_ring18 a_24059_20693 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3630 VPWR a_22711_12533 _185_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X3631 tdc0.r_dly_store_ring19 a_12007_15253 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3632 VGND tdc0.w_ring_norsz13 tdc0.w_ring_int_norsz14 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3634 VPWR a_15196_16073 uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3636 a_16187_19891 _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X3638 tdc0.r_dly_store_ring19 a_12007_15253 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3639 a_15262_13759 a_15094_14013 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3640 VPWR a_4165_13077 a_4055_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3641 a_17029_13647 a_16863_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3642 a_28043_14735 a_27823_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3644 a_29520_12559 _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3645 a_28415_21237 ui_in[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X3646 a_20798_15101 a_20359_14735 a_20713_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3647 a_22527_20327 _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X3648 VPWR _138_ a_14560_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3649 VGND _070_ a_15577_16483 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3650 VPWR net26 a_8859_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3651 a_12029_10205 a_11985_9813 a_11863_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3653 a_21729_11293 tdc1.r_ring_ctr9 a_21623_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X3654 a_24678_14557 a_24363_14423 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3655 a_17838_10383 _060_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3656 a_11950_19605 a_11782_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
R50 VGND net44 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3657 VGND _076_ a_13459_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3658 VGND a_26483_10901 tdc1.r_ring_ctr9 VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3659 a_5809_14735 tdc0.w_ring_buf16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3661 a_30093_15285 a_29927_15285 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3662 VGND net12 tdc0.w_ring_int_norsz2 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3663 VGND net33 a_18703_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3664 a_27587_16885 a_27871_16885 a_27806_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3665 a_12383_19453 a_11601_19087 a_12299_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3666 tdc1.w_ring_int_norsz28 net75 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3667 _017_ _181_ a_21353_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X3671 VPWR a_23363_12711 _177_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3672 a_27687_14709 net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3674 VGND tdc1.r_ring_ctr2 _167_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3675 tdc1.r_ring_ctr0 a_28239_11445 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X3676 a_28331_20937 net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3678 net27 a_8912_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3679 a_7442_12671 a_7274_12925 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3680 a_6503_14013 a_5639_13647 a_6246_13759 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X3681 VGND _080_ a_18324_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3682 VGND tdc1.w_ring_norsz8 a_20083_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3683 a_13909_16073 _089_ a_13993_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3684 VPWR net9 a_21739_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3685 _058_ net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3686 a_26581_18145 _123_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X3688 VGND a_7699_12925 a_7867_12827 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3690 a_29741_11989 a_29523_12393 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3691 VPWR a_7423_16189 a_7591_16091 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3692 a_13611_20327 tdc0.r_dly_store_ring14 a_13785_20203 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3693 VPWR _064_ a_24087_18775 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0662 ps=0.735 w=0.42 l=0.15
X3694 a_3963_10927 a_3339_10933 a_3855_11305 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3695 _014_ _156_ a_2953_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X3696 VPWR a_23358_19605 a_23285_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3697 a_17075_14191 a_16293_14197 a_16991_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3700 a_22595_14887 tdc1.r_dly_store_ctr0 a_22741_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X3701 a_25121_15823 a_24131_15823 a_24995_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3702 a_6173_14013 a_5639_13647 a_6078_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3703 a_25953_14735 a_25787_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3705 _011_ _151_ a_8497_11721 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3706 VGND net68 tdc1.w_ring_int_norsz21 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3707 VPWR tdc1.w_ring_int_norsz16 a_27333_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3708 VGND _188_ _021_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3709 a_28537_20425 net18 tdc1.w_ring_norsz15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3710 VGND a_27127_16885 net18 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3711 VGND a_15227_13077 a_15185_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3714 a_24927_12393 a_24481_12021 a_24831_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3715 _091_ a_16607_20502 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X3716 _089_ a_21463_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3717 a_17121_17461 a_16955_17461 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3718 a_14700_10927 a_14486_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X3720 VGND tdc1.w_ring_int_norsz19 tdc1.w_ring_norsz19 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3722 VGND tdc1.r_dly_store_ring9 a_22937_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X3724 a_11509_19637 a_11343_19637 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3725 a_13656_12393 a_13257_12021 a_13530_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3727 a_29791_15823 a_29571_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X3728 tdc0.w_ring_int_norsz16 net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3729 a_25001_19337 _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
R51 VPWR tt_um_hpretl_tt06_tdc_v2_91.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3731 a_28609_13647 tdc1.r_ring_ctr0 a_28537_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3732 a_18881_18249 tdc1.w_ring_norsz5 a_18797_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3733 a_25079_16189 a_24297_15823 a_24995_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3735 VGND a_17159_14165 a_17117_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3736 tdc0.r_dly_store_ring23 a_12375_19605 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3737 a_17567_10099 tdc1.w_dly_stop5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3738 a_9757_21097 a_8767_20725 a_9631_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3739 a_22995_10357 a_22820_10383 a_23174_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3740 VGND tdc0.w_ring_norsz3 a_10147_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3741 VGND _075_ a_14265_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X3743 a_9757_15823 a_8767_15823 a_9631_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3744 a_27342_19908 a_27142_19753 a_27491_19997 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X3745 a_19407_10383 a_18961_10383 a_19311_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3747 net17 a_27772_16341 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3748 tdc0.r_ring_ctr3 a_12415_11231 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3749 a_25049_13889 a_24831_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3750 a_16272_12559 _021_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3752 VGND _035_ a_11937_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3753 VPWR a_29055_15975 tdc1.r_dly_store_ring12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3754 VGND _198_ _056_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3755 VGND _075_ a_17128_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3756 VPWR net19 _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3757 a_18072_15279 _084_ a_17804_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3758 VPWR a_1368_17429 net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3760 a_22281_12559 _170_ a_22199_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
R52 VGND uio_out[0] sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3761 VGND net30 a_14655_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3762 a_8849_14985 net39 tdc0.w_ring_int_norsz11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3763 a_27722_12015 a_27003_12257 a_27159_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3764 a_17559_11159 _187_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X3766 a_6430_14165 a_6262_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X3767 _080_ a_19860_15797 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3768 VPWR a_9279_21237 net28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3769 _025_ _171_ a_28737_12809 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3770 a_27307_14887 a_27403_14709 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X3771 a_27759_17775 a_27705_17687 a_27659_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X3772 VPWR _069_ a_13173_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3774 a_5989_10933 a_5823_10933 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3776 tdc0.w_ring_buf30 a_6651_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3777 a_14729_12021 a_14563_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3779 a_6262_14191 a_5989_14197 a_6177_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3780 a_16757_16367 tdc1.w_ring_buf20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3781 _048_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3782 VPWR tdc1.w_ring_norsz26 a_23671_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3783 a_13879_10901 a_14082_11059 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X3784 VGND tdc0.w_ring_int_norsz5 tdc0.w_ring_norsz5 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3785 a_7723_10357 _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3786 a_17549_11471 a_17505_11713 a_17383_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3790 VPWR a_11950_13759 a_11877_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3791 VGND net31 a_16127_18549 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3792 a_16180_21237 net32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3793 a_11509_13647 a_11343_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3794 a_27687_14709 net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3795 a_4117_14735 a_4073_14977 a_3951_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3796 VPWR _173_ a_25317_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3797 VPWR a_6246_13759 a_6173_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3799 a_1755_14191 a_1131_14197 a_1647_14569 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3801 VGND tdc1.w_ring_norsz19 a_19991_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3803 _033_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3804 VPWR a_4130_16341 a_4057_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3805 a_19617_19337 tdc1.w_ring_norsz24 a_19533_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3806 VGND a_21331_10901 _182_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X3807 _147_ a_11763_11445 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3810 VPWR tdc0.w_ring_norsz16 a_5087_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3811 VGND a_6430_14165 a_6388_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3812 a_25953_14735 a_25787_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3815 _075_ a_15451_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3816 VGND tdc1.w_ring_int_norsz20 tdc1.w_ring_norsz20 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3817 tdc0.r_ring_ctr12 a_2387_14495 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X3818 tdc0.r_dly_store_ctr7 a_7867_12827 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3819 a_23947_13897 tdc1.r_ring_ctr4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X3820 VPWR a_9004_20149 net21 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3821 a_9401_18543 net21 tdc0.w_ring_norsz5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3822 a_25229_16367 _066_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X3823 VPWR a_15595_20693 a_15511_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3824 a_13183_19631 net24 a_13361_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X3825 a_17383_11471 a_16937_11471 a_17287_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3826 a_2743_12711 _156_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X3828 a_6377_18543 tdc0.w_ring_int_norsz30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3830 VGND tdc0.w_ring_norsz16 tdc0.w_ring_norsz0 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3831 VGND a_24995_16189 a_25163_16091 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3832 VGND a_16175_20938 tdc0.w_ring_buf1 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3833 a_27815_17429 _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X3834 VPWR _076_ a_16269_19414 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.0767 ps=0.785 w=0.42 l=0.15
X3835 _050_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3836 tdc1.r_dly_store_ring8 a_21391_15003 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3837 tdc0.w_ring_norsz15 tdc0.w_ring_norsz31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3838 tdc0.r_ring_ctr9 a_4687_12319 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3840 _198_ a_28915_10927 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3841 a_11417_15101 a_10883_14735 a_11322_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3842 VGND _197_ _034_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3844 VPWR _071_ a_13583_16705 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3845 VPWR tdc0.w_ring_int_norsz28 a_7369_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3846 VGND a_17107_20937 a_17114_20841 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3847 tdc1.r_dly_store_ring2 a_15595_19605 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3848 _103_ a_13827_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X3849 VPWR net37 a_29927_16373 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3850 a_18847_21237 a_19131_21237 a_19066_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X3852 a_11490_14847 a_11322_15101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X3853 a_30263_12319 _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3854 a_28885_21097 a_28338_20841 a_28538_20996 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3855 a_23592_21097 a_23193_20725 a_23466_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3856 VGND tdc0.w_ring_norsz2 tdc0.w_ring_norsz18 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3857 a_21331_10901 _179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X3858 VPWR a_5875_11623 _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X3859 tdc0.w_ring_int_norsz15 tdc0.w_ring_norsz14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3860 a_7657_10383 a_6467_10383 a_7548_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3861 VGND a_14899_10143 a_14833_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3862 a_28254_17277 a_28007_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X3863 a_18130_19631 a_17691_19637 a_18045_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3864 tdc1.w_ring_norsz27 net17 a_27161_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3865 VPWR net32 a_16403_16373 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3866 a_25381_17429 a_25551_17545 a_25509_17571 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3867 VPWR a_24455_17687 _081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3868 a_14486_10927 a_14399_11169 a_14082_11059 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X3869 a_6273_17455 net39 tdc0.w_ring_int_norsz13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3872 a_1129_16367 _165_ a_1047_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3873 tdc1.w_ring_norsz25 net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3874 VPWR _079_ a_13717_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X3875 a_29989_15823 a_29442_16097 a_29642_15797 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X3876 VPWR tdc1.w_ring_norsz18 a_21647_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3877 VPWR net7 a_3339_10933 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3878 tdc0.w_ring_norsz7 tdc0.w_ring_int_norsz7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3879 a_20568_15823 _086_ a_20448_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X3880 VPWR a_28538_20996 a_28467_21097 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X3881 a_4582_15101 a_3505_14735 a_4420_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3882 a_6987_12247 tdc0.r_ring_ctr7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X3883 VGND a_17314_20996 a_17243_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X3884 VPWR net7 a_1223_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3885 a_19602_11837 a_19163_11471 a_19517_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3886 a_6020_14735 a_5621_14735 a_5894_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3887 a_20706_17277 a_20433_16911 a_20621_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X3888 tdc1.w_ring_int_norsz13 net42 a_29105_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3889 _079_ a_17468_15797 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3890 VGND _064_ a_27019_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X3892 a_2093_15823 a_2049_16065 a_1927_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3893 a_11141_16911 a_10975_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3894 tdc0.r_ring_ctr15 a_2479_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3895 _052_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3896 VPWR a_23211_14735 net33 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3897 VPWR a_21971_13335 tdc1.r_dly_store_ctr6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3898 _006_ a_1047_16367 a_1297_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X3900 a_21518_12559 _063_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3901 a_17042_21085 a_16727_20951 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X3902 a_4287_16189 a_3505_15823 a_4203_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3903 tdc0.w_ring_buf15 a_4903_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3904 a_16180_21237 net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3906 a_12153_12559 a_11987_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3908 a_14799_11445 net32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X3909 a_10317_20175 tdc0.w_ring_buf22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3910 VGND tdc0.r_ring_ctr1 a_13559_9545 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3913 VGND a_17470_13759 a_17428_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3914 a_11923_17277 a_11141_16911 a_11839_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3915 a_11908_20009 a_11509_19637 a_11782_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3917 a_15511_19631 a_14729_19637 a_15427_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3918 VGND tdc0.w_ring_norsz21 tdc0.w_ring_int_norsz22 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3919 a_30342_12925 a_29265_12559 a_30180_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3920 VPWR a_26755_19863 tdc1.r_dly_store_ring31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3921 a_9299_11837 _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3922 tdc0.r_dly_store_ctr3 a_14123_11989 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3923 a_3485_15253 tdc0.r_ring_ctr13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X3925 a_13717_17999 a_13551_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3926 VGND a_29427_20693 net38 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3929 tdc0.r_dly_store_ctr3 a_14123_11989 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3930 a_24481_13647 a_24315_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3931 a_13717_14985 tdc0.r_dly_store_ctr0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3932 tdc0.w_ring_int_norsz20 net49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3936 _088_ a_21311_15617 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X3939 VPWR tdc1.r_ring_ctr6 a_24591_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3940 VGND tdc1.w_ring_norsz18 tdc1.w_ring_int_norsz19 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3941 a_5253_16911 a_5087_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3943 a_8477_15279 tdc0.w_ring_buf11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
R53 net69 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3945 net20 a_4443_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3946 VPWR a_8511_17429 a_8427_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3947 a_14549_13103 tdc0.w_ring_buf25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3948 tdc0.w_ring_int_norsz1 net40 a_4909_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3949 VGND tdc0.w_dly_stop5 a_7111_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3950 a_17811_14013 a_17029_13647 a_17727_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3951 VGND a_21339_12533 a_21273_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3952 VPWR a_8603_14165 a_8519_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3954 tdc1.w_ring_norsz4 tdc1.w_ring_norsz20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3955 VGND a_22527_20327 _085_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X3957 a_22517_10383 a_22473_10625 a_22351_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3958 VGND a_26394_14847 a_26352_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X3960 VGND _063_ a_20861_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3961 a_28078_16885 a_27871_16885 a_28254_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3963 VPWR a_7591_13077 a_7507_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3964 VGND a_28599_15797 net36 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3966 VPWR a_13330_13077 a_13257_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X3967 VGND net26 a_8859_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3969 tdc0.r_ring_ctr6 a_7723_10357 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3970 VPWR net35 a_21279_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3971 a_8013_14985 tdc0.w_ring_norsz27 a_7929_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3972 net35 a_23907_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3973 a_21397_15617 _086_ a_21311_15617 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X3974 VGND net27 a_7479_17461 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3975 a_29642_20149 a_29435_20149 a_29818_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X3977 a_24397_19631 _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X3978 a_11697_19631 tdc0.w_ring_buf23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X3979 a_20901_11471 tdc1.r_ring_ctr8 a_20819_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X3981 VPWR tdc0.w_ring_int_norsz6 a_9209_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3982 VGND net34 a_21279_19637 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3983 a_15118_10927 a_14360_11043 a_14555_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X3984 VGND a_27003_12257 a_26964_12131 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3985 a_22093_21263 tdc1.w_ring_buf17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3986 a_7737_16367 tdc0.w_ring_norsz28 a_7653_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3987 _072_ _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3988 VGND tdc1.w_ring_int_norsz5 tdc1.w_ring_norsz5 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3989 VPWR _198_ _049_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3990 a_14039_12015 a_13257_12021 a_13955_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3991 a_19057_12015 tdc1.r_ring_ctr13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X3992 a_29571_20175 a_29435_20149 a_29151_20149 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X3994 a_20989_11471 tdc1.r_ring_ctr9 a_20901_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X3995 a_25571_13621 _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3996 VGND a_9799_20693 a_9757_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3997 a_22711_12533 _170_ a_23109_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X3998 VGND a_4203_16189 a_4371_16091 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3999 VPWR a_30791_16367 a_30959_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4000 a_28169_20425 net18 tdc1.w_ring_norsz31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4001 a_30447_13621 _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4002 a_11509_12015 a_10975_12021 a_11414_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4003 _143_ a_14583_21590 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X4008 VGND net18 tdc1.w_ring_norsz17 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4009 a_27499_11471 a_27149_11471 a_27404_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4010 a_25251_19951 net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4012 a_15926_17277 a_15679_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4014 a_20635_13897 _080_ a_20717_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4016 VPWR a_23063_14013 a_23231_13915 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4017 a_14583_21590 tdc0.r_dly_store_ring7 a_14583_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4018 a_6319_15101 a_5621_14735 a_6062_14847 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4019 a_1644_16911 _006_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4020 VPWR a_18751_21415 tdc1.r_dly_store_ring1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4021 VGND tdc0.w_ring_norsz4 tdc0.w_ring_norsz20 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4023 a_15117_14741 _093_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4024 a_12867_15511 _129_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4025 VGND a_15170_11989 a_15128_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4026 VGND a_7591_19605 a_7549_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4028 a_19355_13103 _188_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4030 VPWR tdc0.w_ring_norsz6 a_8757_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
R54 VGND net74 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4032 tdc1.w_ring_buf23 a_21923_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4033 a_24694_11517 _179_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4034 VPWR net29 a_11987_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4035 VPWR _113_ a_13615_17571 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4036 VPWR a_26426_17687 _104_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.26 ps=2.52 w=1 l=0.15
X4037 a_4674_12015 a_3597_12021 a_4512_12393 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4038 VGND a_4595_11231 a_4529_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4040 VGND tdc0.w_ring_norsz31 a_6007_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4041 VPWR tdc1.r_ring_ctr4 a_26521_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4043 VGND a_12042_19199 a_12000_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4044 VPWR tdc1.r_dly_store_ctr3 a_22281_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X4045 a_5273_17455 tdc0.w_ring_int_norsz17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4046 VPWR net30 a_16127_14197 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4047 a_21718_19631 a_21445_19637 a_21633_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4048 VPWR a_5767_19453 a_5935_19355 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4049 a_22995_10357 _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4051 VPWR a_5859_16189 a_6027_16091 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4053 a_12815_17455 _071_ a_12897_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4054 VPWR a_16991_14191 a_17159_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4055 VPWR a_24462_14847 a_24389_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4056 a_10521_16367 tdc0.w_ring_norsz18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4057 tdc1.r_dly_store_ring18 a_24059_20693 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4059 a_17773_19337 net14 tdc1.w_ring_norsz6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4060 VPWR a_25932_12533 net9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4061 _022_ _188_ a_19605_13423 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X4063 VPWR a_18539_13077 a_18455_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4064 VPWR tdc0.w_ring_norsz5 a_10331_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4065 tdc1.r_ring_ctr1 a_30263_12319 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X4066 VPWR a_11379_12925 a_11547_12827 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4067 uo_out[7] a_14172_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X4069 VPWR net9 a_26983_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4070 a_19395_17076 tdc1.w_ring_norsz5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4071 a_7975_18543 a_7111_18549 a_7718_18517 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4072 a_22353_12559 _172_ a_22281_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4073 VPWR a_23891_20719 a_24059_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4074 VPWR tdc1.w_ring_buf29 a_30725_18921 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4077 VGND a_27894_14709 a_27823_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X4079 VGND a_863_13897 _003_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X4080 a_21768_14191 _193_ a_21666_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4081 VPWR a_11839_15279 a_12007_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4083 tdc0.w_ring_int_norsz14 net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4084 a_13551_10633 tdc0.r_ring_ctr1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X4085 VPWR a_19876_10383 a_20051_10357 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4087 VGND a_11839_15279 a_12007_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4088 VGND a_13603_11445 _146_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X4089 a_15282_16073 _103_ a_15196_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4090 a_11509_13647 a_11343_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4091 VPWR net8 a_9411_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4092 _051_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4093 a_17107_12533 a_16932_12559 a_17286_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4094 a_7645_18543 a_7111_18549 a_7550_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4095 a_14560_20425 _138_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4096 _193_ a_20635_13897 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4099 a_14172_20149 _089_ a_14560_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4100 VPWR tdc1.r_ring_ctr15 a_19437_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4102 VPWR tdc1.r_ring_ctr4 a_25297_14569 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4103 VGND _089_ a_14300_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X4104 a_4687_13407 a_4512_13481 a_4866_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4105 a_15750_16885 a_15543_16885 a_15926_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X4106 a_27679_21237 net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X4108 a_12299_19453 a_11435_19087 a_12042_19199 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4109 tdc1.r_ring_ctr15 a_21339_12533 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4110 a_20874_17023 a_20706_17277 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4111 a_3601_12559 tdc0.r_ring_ctr9 a_3513_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4112 _190_ a_12447_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4114 a_7258_11293 _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4116 VGND tdc1.r_dly_store_ring16 a_23029_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4117 a_24939_12015 _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4118 a_16658_15279 a_16481_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X4119 VGND tdc1.w_ring_norsz4 tdc1.w_ring_int_norsz5 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4120 a_2965_14735 tdc0.r_ring_ctr13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R55 VGND net49 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4121 VGND _045_ a_4117_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4124 a_16301_16073 _069_ a_16155_15975 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X4125 _138_ a_13921_19747 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X4126 VPWR tdc0.w_ring_norsz25 a_11067_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4127 a_15679_16911 a_15543_16885 a_15259_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4128 a_16823_20951 a_17107_20937 a_17042_21085 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4129 a_11237_14735 tdc0.w_ring_buf26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4130 VPWR a_2212_13481 a_2387_13407 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4131 tdc0.r_dly_store_ring10 a_10443_15003 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4132 a_13173_14191 tdc0.r_dly_store_ring27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4133 VGND net36 a_25787_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4135 tdc1.w_ring_int_norsz21 tdc1.w_ring_norsz20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4136 _136_ a_12815_17455 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X4137 _021_ _189_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4138 net18 a_27127_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4140 a_14560_20425 _089_ a_14172_20149 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X4141 a_13459_18543 _089_ a_13637_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4142 a_27304_10927 a_27090_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X4143 VPWR a_22327_11837 a_22495_11739 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4144 VPWR tdc0.w_dly_stop5 a_4443_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4146 a_7548_10383 a_6633_10383 a_7201_10625 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4148 tdc1.w_ring_norsz19 tdc1.w_ring_norsz3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4149 a_19419_10749 a_18795_10383 a_19311_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4150 VGND net27 a_7111_18549 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4151 tdc0.r_dly_store_ring9 a_15687_13915 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4152 a_24777_17821 _065_ a_24677_17821 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X4157 a_18797_18249 tdc1.w_ring_int_norsz21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4158 tdc0.w_ring_norsz29 net22 a_6921_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4159 tdc1.w_ring_buf29 a_30295_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4160 a_23653_10159 tdc1.r_ring_ctr8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4162 a_14545_14985 tdc0.r_dly_store_ctr3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4164 a_15427_19631 a_14729_19637 a_15170_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4165 a_14797_21590 tdc0.r_dly_store_ring7 a_14583_21590 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X4166 a_15002_20719 a_14729_20725 a_14917_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4167 a_4055_13103 a_3431_13109 a_3947_13481 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4170 tdc1.w_ring_norsz7 net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4171 VGND _173_ _176_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4172 VPWR a_13735_21263 _076_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4174 VPWR a_3295_19252 tdc0.w_dly_stop1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4175 a_17804_15279 _084_ a_18072_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4176 _047_ net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4177 VGND tdc1.w_ring_buf4 a_16097_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4178 net7 a_1368_17429 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4179 VPWR a_7718_18517 a_7645_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4182 VPWR tdc0.w_ring_norsz12 a_6273_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4183 a_6725_15823 a_6559_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4184 VPWR a_3851_13621 _002_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X4185 net28 a_9279_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4186 a_14641_19087 tdc0.w_ring_buf2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4188 a_26933_19337 _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X4191 a_28713_18249 tdc1.w_ring_norsz13 a_28629_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4192 a_3877_16367 tdc0.r_ring_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4193 a_19876_10383 a_18795_10383 a_19529_10625 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4194 VGND _046_ a_2093_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4195 a_19267_20425 tdc1.r_dly_store_ring6 a_19065_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4197 _045_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4198 VPWR a_12507_10143 tdc0.r_ring_ctr0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4199 VPWR _069_ a_12161_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4200 a_4088_16745 a_3689_16373 a_3962_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4201 VGND a_26297_20340 tdc1.w_ring_buf0 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4202 tdc1.r_dly_store_ring23 a_23783_19605 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4203 a_24481_13647 a_24315_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4205 a_4687_12319 a_4512_12393 a_4866_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4206 VPWR net34 a_21739_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4207 a_21817_11471 tdc1.r_ring_ctr9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4208 tdc1.r_dly_store_ring23 a_23783_19605 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4209 VGND _036_ a_10189_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4211 VPWR _191_ a_17720_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X4212 VPWR a_12415_11231 a_12402_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4214 a_23542_10901 a_23374_10927 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4215 VGND net9 a_16403_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4216 a_9773_19631 tdc0.w_ring_norsz7 a_9689_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4217 a_1297_14197 a_1131_14197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4218 a_24738_15935 a_24570_16189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4219 _075_ a_15451_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X4220 a_20798_15101 a_20525_14735 a_20713_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4221 a_17395_11837 a_16771_11471 a_17287_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4223 VPWR a_25623_11247 _031_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X4224 a_25295_15497 net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4226 VPWR net36 a_25787_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
R56 tdc0.g_ring322.stg01_51.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4229 a_3854_17023 a_3686_17277 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4230 VPWR a_25221_19605 _087_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4231 VPWR a_7699_12925 a_7867_12827 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4232 VGND net29 a_10883_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4234 a_4529_11305 a_3339_10933 a_4420_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4236 a_29791_20938 tdc1.w_ring_norsz15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4237 _046_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4238 VGND a_10846_15935 a_10804_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4239 VPWR a_27403_17973 net24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4242 tdc0.w_ring_norsz0 tdc0.w_ring_int_norsz0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4243 tdc1.w_ring_norsz30 net17 a_29553_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R57 net62 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4244 a_6913_19631 tdc0.w_ring_buf31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4245 a_13344_20693 _132_ a_13732_21039 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4248 a_14724_10217 a_13809_9845 a_14377_9813 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4251 VGND a_7607_20541 a_7775_20443 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4252 _009_ _148_ a_11533_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4253 tdc1.w_dly_stop2 a_15575_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4254 a_17691_12559 tdc1.r_ring_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X4255 a_28241_14735 a_27694_15009 a_27894_14709 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4256 tdc0.r_dly_store_ring21 a_9799_16091 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4257 a_10773_16189 a_10239_15823 a_10678_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4258 VGND _058_ a_22517_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4259 a_21629_11471 a_21463_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4260 VGND tdc1.w_ring_norsz21 tdc1.w_ring_int_norsz22 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4261 a_13583_16705 tdc0.r_dly_store_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4262 a_7369_16367 tdc0.w_ring_norsz12 a_7285_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4263 a_5893_19087 a_4903_19087 a_5767_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4264 _113_ a_13583_16705 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X4266 tdc1.r_dly_store_ctr12 a_17895_13915 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4267 a_1939_16189 a_1315_15823 a_1831_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4270 a_30281_16367 tdc1.w_ring_buf28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4271 VPWR a_15719_21237 net32 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4273 VPWR net8 a_11159_10933 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4274 VPWR tdc0.w_ring_norsz7 a_11251_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4275 VPWR a_24546_20327 _142_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X4276 a_27090_10927 a_27003_11169 a_26686_11059 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X4278 a_22729_21263 a_21739_21263 a_22603_21629 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4279 tdc0.w_dly_stop2 a_2971_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4280 _031_ _180_ a_25953_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X4281 a_12079_16073 _080_ a_12161_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X4282 VGND a_6027_16091 a_5985_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4284 a_27561_13469 a_27182_13103 a_27489_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4286 a_6987_12247 tdc0.r_ring_ctr6 a_7161_12353 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4287 a_19395_17076 tdc1.w_ring_norsz5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4291 VGND _076_ a_17047_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4292 VGND tdc0.w_ring_norsz25 a_11067_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4293 a_27772_16341 net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4294 a_16629_12559 a_16585_12801 a_16463_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4295 VPWR a_7159_17076 tdc0.w_ring_buf29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4296 a_26747_18863 tdc1.r_dly_store_ring21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X4297 a_11881_21263 tdc0.w_ring_buf7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4299 VGND net31 a_10975_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4300 a_14116_17999 a_13717_17999 a_13990_18365 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4302 a_17010_16341 a_16842_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4303 net33 a_23211_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X4304 a_9765_14735 tdc0.w_ring_buf10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4305 a_9347_17277 a_8565_16911 a_9263_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4307 _173_ a_24347_13441 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X4308 VGND a_19735_11989 a_19693_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4309 a_12618_21039 tdc0.r_dly_store_ring6 a_12537_21039 VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.0829 ps=0.905 w=0.65 l=0.15
X4310 VGND a_17208_20149 uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X4311 VGND net29 a_11987_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4312 a_24409_18909 _065_ a_24309_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X4317 a_16301_15823 net25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X4318 a_25149_12809 tdc1.r_ring_ctr6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4319 a_15427_19631 a_14563_19637 a_15170_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4320 a_9409_11713 a_9191_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4322 VGND a_24251_19863 _097_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4324 net38 a_29427_20693 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R58 uio_oe[3] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4325 a_27491_19997 a_27271_20009 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X4326 tdc1.w_ring_int_norsz18 net65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4327 VPWR a_6855_14165 a_6771_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4328 _036_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4329 _042_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4330 VPWR net10 a_24315_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4331 _116_ a_13461_17571 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X4332 a_8469_17833 a_7479_17461 a_8343_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4333 tdc1.r_dly_store_ring19 a_21299_17179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4334 VGND _089_ a_17678_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4336 a_18059_17161 _109_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X4337 a_11509_17277 a_10975_16911 a_11414_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4338 a_15097_19631 a_14563_19637 a_15002_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4339 a_21331_10901 tdc1.r_ring_ctr9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X4340 VPWR tdc0.w_ring_int_norsz31 a_5529_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4342 VPWR net29 a_10883_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4344 VPWR a_10846_15935 a_10773_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4345 VGND net27 a_5087_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4346 a_11693_21263 a_11527_21263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4347 a_24546_20327 _141_ a_24849_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X4348 VGND tdc0.w_ring_norsz6 tdc0.w_ring_norsz22 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4350 tdc0.w_ring_buf4 a_12355_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4353 _007_ a_13559_9545 a_13809_9545 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X4354 VPWR tdc0.w_ring_norsz22 a_9769_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4355 a_15002_19631 a_14563_19637 a_14917_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4356 tdc1.w_ring_buf28 a_29743_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4357 a_4073_10901 a_3855_11305 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4358 a_10601_13897 tdc0.w_ring_norsz9 a_10517_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4360 a_17727_14013 a_16863_13647 a_17470_13759 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4361 tdc1.w_ring_buf9 a_20727_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4362 a_15427_12015 a_14729_12021 a_15170_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4363 a_12291_14013 a_11509_13647 a_12207_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4366 a_21349_14735 a_20359_14735 a_21223_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4368 tdc0.w_ring_int_norsz19 net48 a_10521_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4371 net36 a_28599_15797 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4372 a_18497_13481 a_17507_13109 a_18371_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4373 a_945_13897 _162_ a_863_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4375 a_17397_14013 a_16863_13647 a_17302_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4376 a_17267_16367 a_16569_16373 a_17010_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4377 a_14729_20725 a_14563_20725 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4379 a_7929_14985 net23 tdc0.w_ring_norsz11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4381 VGND a_29467_15287 _627_.X VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4383 a_7925_14191 tdc0.w_ring_buf27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4384 a_1865_13077 a_1647_13481 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4385 a_23316_20009 a_22917_19637 a_23190_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4386 a_25892_19951 net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4387 net19 a_4404_19061 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4391 VGND a_24835_13335 _172_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X4392 a_12594_11293 _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4393 VPWR _028_ a_27722_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X4394 a_5621_14735 a_5455_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4395 a_17470_13759 a_17302_14013 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4396 a_9209_19631 tdc0.w_ring_norsz22 a_9125_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4397 a_17946_13103 a_17673_13109 a_17861_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4398 a_22281_14191 _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
R59 VPWR tt_um_hpretl_tt06_tdc_v2_87.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4399 a_24131_19337 _072_ a_24213_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4400 a_29151_20149 a_29442_20449 a_29393_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X4403 a_23500_17833 a_23101_17461 a_23374_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4404 a_25085_19337 _065_ a_25001_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4405 a_11448_14735 a_11049_14735 a_11322_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4408 VPWR a_22311_19605 a_22227_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4410 a_26651_15101 a_25787_14735 a_26394_14847 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4411 VGND _076_ a_15801_19414 VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X4412 VPWR tdc1.r_ring_ctr1 a_28455_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4413 a_21934_20221 _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4414 tdc1.w_ring_int_norsz24 net71 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4415 VPWR a_24087_18775 _129_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4416 a_2479_16885 a_2304_16911 a_2658_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4417 VPWR a_24819_17776 a_24455_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X4419 VGND a_9263_17277 a_9431_17179 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4420 VPWR a_10570_20287 a_10497_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4421 VGND a_11490_18111 a_11448_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4424 a_30534_16341 a_30366_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4425 a_27499_11471 a_26983_11471 a_27404_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4426 a_27518_19631 a_27271_20009 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X4427 a_30917_15657 a_29927_15285 a_30791_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4428 VGND tdc1.w_ring_norsz26 a_23671_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4430 tdc0.r_dly_store_ctr1 a_15595_11989 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4431 VGND a_7166_15935 a_7124_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4432 a_7423_16189 a_6559_15823 a_7166_15935 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4433 a_22741_14735 _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X4436 tdc1.w_ring_int_norsz10 net41 a_21009_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4438 VGND tdc1.w_dly_stop3 a_16311_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4439 a_17562_17429 a_17394_17455 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4440 VPWR a_16656_16885 uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4441 a_9025_10633 tdc0.r_ring_ctr4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4443 a_9927_10383 a_9411_10383 a_9832_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4444 a_14899_10143 a_14724_10217 a_15078_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4445 a_3597_13109 a_3431_13109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4446 VGND _094_ a_15117_14741 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4447 a_22411_11837 a_21629_11471 a_22327_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4448 VPWR a_5875_13077 _160_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X4449 a_7093_16189 a_6559_15823 a_6998_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4451 _043_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4452 VPWR net33 a_19255_14197 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4453 VGND a_12415_11231 a_12349_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4454 a_17394_17455 a_17121_17461 a_17309_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4455 a_23105_19631 tdc1.w_ring_buf23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4456 VPWR _068_ a_13349_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X4457 VPWR a_8730_15253 a_8657_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4458 VPWR a_21463_15823 _089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4459 VGND tdc0.w_ring_norsz16 a_5087_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4460 a_14570_17494 _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X4461 a_11831_18365 a_11049_17999 a_11747_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4463 a_24455_17687 a_24819_17776 a_24777_17821 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4465 VGND _194_ a_21337_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X4466 VPWR a_17137_10625 a_17027_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X4467 a_26895_17429 _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X4468 VGND tdc1.r_dly_store_ring6 a_19349_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X4470 a_7825_12559 a_6835_12559 a_7699_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4472 tdc0.w_dly_stop2 a_2971_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4474 _141_ a_23855_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4475 tdc0.w_ring_norsz27 net23 a_8577_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4477 tdc0.r_dly_store_ctr2 a_13755_13077 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4479 _171_ _168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4480 _137_ a_13183_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4481 a_4595_14709 a_4420_14735 a_4774_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4482 a_21257_16911 a_20267_16911 a_21131_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4483 a_16825_15797 _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X4484 tdc0.w_ring_buf20 a_10331_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4486 VPWR tdc0.r_ring_ctr9 a_2623_12335 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X4487 a_11379_12925 a_10681_12559 a_11122_12671 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4489 a_15511_12015 a_14729_12021 a_15427_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4490 VGND a_22247_20938 tdc1.w_ring_buf17 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4491 VGND tdc1.w_ring_norsz0 tdc1.w_ring_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4492 a_23925_11305 a_22935_10933 a_23799_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4493 VGND net25 a_13069_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4495 a_13485_11293 tdc0.r_ring_ctr2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X4496 a_29791_18775 a_29887_18775 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4498 a_15110_16073 _102_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X4499 a_19065_20425 _075_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X4500 a_27659_17775 _067_ a_27555_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X4502 VPWR net33 a_16863_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4503 VPWR a_25103_16599 _098_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X4504 a_7645_17461 a_7479_17461 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4505 a_22247_20938 tdc1.w_ring_norsz17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4506 VPWR a_19310_11989 a_19237_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4507 a_22343_15975 _081_ a_22671_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4508 a_13633_15279 tdc0.r_dly_store_ring10 a_13551_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4509 _175_ a_24591_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X4510 tdc0.w_ring_norsz16 net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4511 a_5621_14735 a_5455_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4513 a_22487_13481 a_22351_13321 a_22067_13335 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X4514 a_26813_13469 a_26778_13235 a_26575_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X4515 a_18239_16073 _084_ a_18021_15797 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4516 a_17394_17455 a_16955_17461 a_17309_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4519 VPWR net33 a_19163_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4521 VPWR tdc1.w_dly_stop2 a_15759_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4522 VGND tdc1.w_ring_norsz13 tdc1.w_ring_int_norsz14 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4524 VGND a_16182_14847 a_16140_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4525 VGND a_16734_18517 a_16692_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X4527 a_14300_16911 _117_ a_14032_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4528 VPWR a_27135_19849 a_27142_19753 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4529 a_5349_15823 tdc0.r_ring_ctr13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4530 net39 a_9839_17715 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4531 VGND a_26615_13647 net10 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4532 tdc0.w_ring_buf15 a_4903_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4533 a_29265_12559 a_29099_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4536 a_5875_13077 tdc0.r_ring_ctr8 a_6273_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X4538 VGND a_7159_17076 tdc0.w_ring_buf29 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4539 a_17107_20937 net34 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4540 a_20316_18151 _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X4541 VPWR a_7166_15935 a_7093_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X4542 a_16991_18543 a_16293_18549 a_16734_18517 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4543 VGND tdc1.w_ring_norsz29 tdc1.w_ring_norsz13 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4545 a_20635_13897 _080_ a_20717_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4546 a_3760_14735 _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4547 _076_ a_13735_21263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X4548 VPWR net20 _044_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4550 a_29723_12925 a_29099_12559 a_29615_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X4551 a_17117_18921 a_16127_18549 a_16991_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X4553 _022_ a_19355_13103 a_19605_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X4554 VPWR tdc1.r_ring_ctr8 _180_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4555 a_14802_13077 a_14634_13103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4556 a_2387_13407 _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4557 a_29057_21428 ui_in[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4558 a_30875_16367 a_30093_16373 a_30791_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4559 a_21718_18543 a_21279_18549 a_21633_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4560 a_27517_18543 a_27351_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X4561 tdc1.w_ring_norsz14 net17 a_29185_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4562 a_21729_16367 tdc1.r_dly_store_ring27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X4563 a_14428_17687 tdc0.r_dly_store_ring4 a_14570_17494 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
R60 VPWR tdc1.g_ring317.stg01_64.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4564 a_9715_20719 a_8933_20725 a_9631_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4565 a_3597_12021 a_3431_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4566 a_22327_11837 a_21629_11471 a_22070_11583 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4568 VPWR tdc0.r_ring_ctr7 a_6340_11721 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X4569 VPWR a_15319_19355 a_15235_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4572 VGND a_5087_11471 _197_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4575 VGND a_15519_14013 a_15687_13915 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4576 a_18146_12335 tdc1.r_ring_ctr12 _189_ VGND sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.106 ps=0.975 w=0.65 l=0.15
X4578 a_15002_12015 a_14563_12021 a_14917_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4579 a_2571_15797 a_2396_15823 a_2750_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4580 net20 a_4443_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4581 a_21971_13335 a_22067_13335 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X4582 net34 a_23264_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4583 a_23363_12711 tdc1.r_ring_ctr7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X4585 VGND tdc1.r_ring_ctr8 a_23403_9839 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4586 a_1747_15645 _162_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X4587 net30 a_16162_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4588 VGND tdc1.w_ring_norsz15 tdc1.w_ring_int_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4591 a_3431_12559 tdc0.r_ring_ctr10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X4592 VPWR a_23996_16599 _099_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X4596 tdc1.w_ring_buf28 a_29743_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4597 a_28007_16911 a_27878_17185 a_27587_16885 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4600 a_10528_20175 a_10129_20175 a_10402_20541 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4601 net40 a_9963_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4602 a_22645_19087 tdc1.w_ring_buf10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4603 VGND net37 a_29651_17461 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4604 VPWR tdc1.r_dly_store_ring17 a_22653_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X4605 VGND a_9891_12827 a_9849_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4607 a_27645_15101 a_27307_14887 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4608 a_14117_11293 a_14082_11059 a_13879_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X4609 a_8470_13103 a_8031_13109 a_8385_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4610 VGND a_8511_17429 a_8469_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4611 VPWR net4 a_25287_18517 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X4613 VPWR _165_ a_1297_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4614 a_17505_11713 a_17287_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4615 a_6059_11989 _155_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X4618 a_28629_18249 net17 tdc1.w_ring_norsz29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4619 a_13625_18543 tdc0.r_dly_store_ring13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X4620 VGND _175_ a_24920_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X4621 a_13162_13103 a_12723_13109 a_13077_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4622 VGND a_22311_19605 a_22269_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4623 a_23975_20719 a_23193_20725 a_23891_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
R61 net65 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4624 a_21718_12015 a_21445_12021 a_21633_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4625 a_16941_15279 a_16764_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X4626 a_19065_20425 _089_ a_19267_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4628 VGND net43 a_9963_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X4629 a_12686_10205 _032_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4630 VGND net10 a_24315_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4634 VPWR tdc1.w_ring_norsz6 a_18509_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4635 VPWR _178_ a_23211_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4636 _038_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4637 a_13633_14985 _083_ a_13717_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R62 net56 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4639 VPWR a_10443_15003 a_10359_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4640 a_28047_20951 a_28331_20937 a_28266_21085 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4642 VGND a_26575_13077 tdc1.r_ring_ctr4 VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X4643 a_17720_15279 _192_ a_17804_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4644 VPWR tdc0.w_ring_int_norsz11 a_8013_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4645 a_9689_19631 tdc0.w_ring_int_norsz23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4647 a_17405_19631 net14 tdc1.w_ring_norsz23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4648 a_7902_10383 _038_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4649 VPWR net34 a_17691_19637 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4650 VPWR _147_ a_8767_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X4651 VGND _172_ a_24433_13441 VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4652 a_12349_11305 a_11159_10933 a_12240_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4653 a_14361_13109 a_14195_13109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4654 a_16824_10383 _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4655 a_18249_12335 tdc1.r_ring_ctr13 a_18146_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X4656 a_2785_10927 _156_ a_2703_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4657 VGND a_25295_15497 a_25302_15401 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4658 VPWR a_17107_12533 a_17094_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4659 VGND a_28415_21237 net3 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4660 VPWR a_12875_20327 _128_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4661 tdc0.w_ring_buf20 a_10331_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4662 _095_ a_15117_14741 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X4663 VPWR a_18555_19631 a_18723_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4664 VPWR net33 a_22935_10933 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4665 VPWR tdc1.r_dly_store_ctr2 a_25229_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X4666 a_19131_21237 net34 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4667 VGND a_18555_19631 a_18723_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4668 a_16055_19087 a_15801_19414 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.145 ps=1.11 w=0.42 l=0.15
X4669 tdc0.w_ring_norsz2 tdc0.w_ring_norsz18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4672 a_16293_14197 a_16127_14197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4673 a_19089_21629 a_18751_21415 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4674 a_7277_18549 a_7111_18549 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4676 VGND a_12507_10143 a_12441_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4679 a_12989_16367 tdc0.r_dly_store_ring17 a_12907_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4680 a_20621_16911 tdc1.w_ring_buf19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4681 tdc0.r_dly_store_ring13 a_8143_18517 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4682 VGND a_30959_15253 a_30917_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4683 VGND tdc0.w_ring_norsz5 a_10331_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4684 a_21185_10633 _181_ a_21103_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4685 _033_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4686 tdc1.w_ring_int_norsz22 net69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4687 tdc0.r_dly_store_ring13 a_8143_18517 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4688 VPWR _083_ a_14197_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4690 uo_out[0] a_17804_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4691 a_14453_19087 a_14287_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4692 VPWR _184_ a_17862_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X4693 VPWR net29 a_13091_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4694 net32 a_15719_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4695 VGND tdc1.w_ring_norsz14 tdc1.w_ring_int_norsz15 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4696 a_3852_12381 _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X4697 a_30258_17429 a_30090_17455 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4698 a_26851_15797 a_27135_15797 a_27070_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X4699 _065_ a_27259_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4700 VGND a_7723_10357 a_7657_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4702 VGND tdc1.w_ring_int_norsz2 tdc1.w_ring_norsz2 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4704 _062_ net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4705 VGND _182_ a_20169_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4706 VGND a_6796_17973 net22 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X4707 a_30090_17455 a_29817_17461 a_30005_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4709 a_5560_15823 a_5161_15823 a_5434_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4712 a_14195_18863 _120_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X4714 a_9807_12925 a_9025_12559 a_9723_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4715 a_14726_19453 a_14287_19087 a_14641_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4716 a_10613_18249 tdc0.w_ring_norsz2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4717 a_14570_17821 _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X4718 VPWR _126_ a_14372_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.14 ps=1.28 w=1 l=0.15
X4720 a_26513_20719 net18 tdc1.w_ring_norsz0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4722 a_8136_14569 a_7737_14197 a_8010_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4723 a_30093_15285 a_29927_15285 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4724 net41 a_26031_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4725 a_18555_19631 a_17691_19637 a_18298_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4727 a_1368_17429 tdc0.w_ring_buf0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4728 a_26805_16367 tdc1.w_ring_norsz26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4729 VGND a_26651_15101 a_26819_15003 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4730 uo_out[1] a_17208_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4732 tdc1.r_dly_store_ring24 a_20287_14165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4734 VGND _057_ a_26721_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X4735 VPWR a_9103_12247 _149_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4737 a_9096_11471 _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X4738 a_8059_18543 a_7277_18549 a_7975_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4739 a_24467_16599 _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X4740 a_21902_11837 a_21463_11471 a_21817_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4741 tdc0.r_ring_ctr10 a_2387_13407 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X4742 a_13698_11989 a_13530_12015 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4743 a_27012_18249 _121_ a_26910_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X4744 a_19267_21263 a_19138_21537 a_18847_21237 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4745 a_19149_16367 tdc1.w_ring_buf5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4746 a_25203_10357 a_25028_10383 a_25382_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4747 tdc1.w_ring_int_norsz16 tdc1.w_ring_norsz15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4748 tdc0.w_ring_norsz21 net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4749 VGND net16 _060_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4750 a_6071_13469 tdc0.r_ring_ctr11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X4751 VPWR tdc1.r_dly_store_ring15 a_25111_20327 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4752 a_17678_20175 _091_ a_17208_20149 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4753 VGND _198_ _051_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R63 VGND net71 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4754 uo_out[2] a_16656_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R64 net59 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4756 a_25520_18903 net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.127 ps=1.1 w=0.42 l=0.15
X4757 tdc0.w_ring_norsz4 tdc0.w_ring_int_norsz4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4758 a_17137_10625 a_16919_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4759 VGND tdc1.w_ring_norsz26 tdc1.w_ring_norsz10 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4761 a_5529_18543 net13 a_5445_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4763 a_11893_10901 a_11675_11305 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X4764 VPWR tdc1.r_dly_store_ring8 a_21768_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
R65 VPWR tt_um_hpretl_tt06_tdc_v2_84.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4765 VGND tdc0.w_ring_int_norsz16 tdc0.w_ring_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4766 VPWR net31 a_11527_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4767 tdc0.w_ring_norsz22 tdc0.w_ring_int_norsz22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4768 tdc1.w_dly_stop3 a_15759_10927 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4769 VGND tdc0.w_ring_norsz30 tdc0.w_ring_int_norsz31 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4770 VGND a_8143_18517 a_8101_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4771 VGND net33 a_16863_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4772 a_10517_13897 tdc0.w_ring_int_norsz25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4773 tdc0.r_dly_store_ring20 a_11915_18267 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4775 a_6557_10901 a_6339_11305 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X4777 VPWR a_10667_10357 a_10654_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4778 a_12207_14013 a_11343_13647 a_11950_13759 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4779 VGND a_30166_18111 a_30124_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
R66 VPWR tdc1.g_ring329.stg01_76.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4781 a_7166_13077 a_6998_13103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4782 _163_ tdc0.r_ring_ctr12 a_2965_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4783 a_25253_15279 a_24915_15511 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X4784 a_15577_16483 _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4786 a_5791_12533 _147_ a_6272_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X4787 VPWR tdc1.w_dly_stop5 a_28915_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4788 a_9781_18543 tdc0.w_ring_int_norsz21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4789 VPWR a_12867_15511 _130_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X4790 a_8841_11471 a_8675_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4791 VGND a_23055_15975 _110_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4793 VGND a_3295_19252 tdc0.w_dly_stop1 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4795 a_19419_10749 _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4796 a_13557_11293 tdc0.r_ring_ctr0 a_13485_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4797 a_12441_10217 a_11251_9845 a_12332_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4798 VGND a_27687_14709 a_27694_15009 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R67 uio_out[2] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4799 VPWR a_7607_20541 a_7775_20443 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4800 a_10957_13897 tdc0.w_ring_norsz25 a_10873_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4801 VPWR tdc0.w_ring_int_norsz10 a_10037_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4802 VPWR a_26031_16885 net41 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4803 a_29265_12559 a_29099_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4804 a_20203_14191 a_19421_14197 a_20119_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4806 tdc1.w_ring_norsz15 tdc1.w_ring_norsz31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4807 a_11582_17023 a_11414_17277 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4808 a_28279_12015 tdc1.r_ring_ctr0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4809 a_23363_12711 tdc1.r_ring_ctr6 a_23537_12587 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4811 a_10129_20175 a_9963_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4812 a_28064_11471 a_26983_11471 a_27717_11713 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X4813 a_1129_12809 a_1099_12744 _001_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X4814 a_12042_19199 a_11874_19453 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4815 a_19820_14569 a_19421_14197 a_19694_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4816 VPWR tdc0.w_ring_norsz14 a_6283_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4817 a_4117_11293 a_4073_10901 a_3951_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4820 a_9206_20719 a_8767_20725 a_9121_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4821 a_27333_20719 net62 a_27249_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R68 net79 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4823 VGND net25 a_24201_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X4824 tdc1.w_ring_buf18 a_21647_20719 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4825 a_9206_16189 a_8767_15823 a_9121_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4826 a_20599_12559 a_20083_12559 a_20504_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4828 VPWR _088_ a_21463_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4829 a_3897_18543 tdc0.w_ring_norsz31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4831 a_22093_21263 tdc1.w_ring_buf17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4832 a_11966_21629 a_11527_21263 a_11881_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4835 a_1099_12744 _158_ a_1485_12809 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4836 a_24835_13335 tdc1.r_ring_ctr4 a_25009_13441 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4839 a_9850_15101 a_9411_14735 a_9765_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X4840 VGND a_22135_14423 _107_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4842 VPWR a_27342_15797 a_27271_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X4843 a_8688_15657 a_8289_15285 a_8562_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4845 _023_ tdc1.r_ring_ctr0 a_28529_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
R69 uio_oe[2] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4847 _040_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4848 a_21361_20719 net15 tdc1.w_ring_norsz18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4849 a_22327_11837 a_21463_11471 a_22070_11583 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4853 VPWR net26 a_8031_13109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4855 a_24677_17821 _064_ a_24589_17821 VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X4858 VGND net17 tdc1.w_ring_norsz28 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4859 a_11763_11445 _146_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X4860 _089_ a_21463_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4861 VPWR a_8895_13103 a_9063_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4863 a_30725_18921 a_30178_18665 a_30378_18820 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4865 a_11747_18365 a_10883_17999 a_11490_18111 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4866 VGND a_11915_15003 a_11873_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4867 VGND a_8895_13103 a_9063_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4868 a_22553_13647 tdc1.r_ring_ctr15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4869 a_20027_11837 a_19163_11471 a_19770_11583 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4871 VGND a_14555_10901 a_14486_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4872 VPWR a_17435_16341 a_17351_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4873 VPWR tdc0.w_ring_norsz15 a_5087_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4875 a_17395_11837 _061_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X4876 a_8577_14985 tdc0.w_ring_norsz11 a_8493_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4877 a_8101_18921 a_7111_18549 a_7975_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
R70 VPWR tt_um_hpretl_tt06_tdc_v2_89.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4878 a_25425_12809 _175_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4879 VGND net29 a_14563_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4881 a_19697_11837 a_19163_11471 a_19602_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4882 tdc1.w_ring_norsz26 tdc1.w_ring_int_norsz26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4883 VPWR _179_ a_23653_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4884 VGND net37 a_29927_16373 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4885 a_19402_16341 a_19234_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4886 a_25297_14569 a_24750_14313 a_24950_14468 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X4888 a_3701_14511 _161_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4889 a_23174_10383 _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X4890 a_15427_12015 a_14563_12021 a_15170_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4892 VGND a_18731_17063 _133_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4893 a_19241_15279 net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X4894 VGND net32 a_16403_16373 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4895 a_29370_15823 a_29055_15975 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X4897 a_7166_15935 a_6998_16189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4898 a_13905_17999 tdc0.w_ring_buf4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4900 VGND a_6503_14013 a_6671_13915 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4901 VPWR a_27687_14709 a_27694_15009 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4902 a_30492_14569 a_30093_14197 a_30366_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X4903 a_15097_12015 a_14563_12021 a_15002_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4904 a_11049_14735 a_10883_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4906 VPWR a_7111_17999 net23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4909 VGND tdc1.w_ring_buf11 a_28425_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X4910 a_19533_19337 tdc1.w_ring_int_norsz8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4911 a_14894_19199 a_14726_19453 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X4913 a_11187_16189 a_10405_15823 a_11103_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4914 a_11322_18365 a_11049_17999 a_11237_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X4915 a_4582_10927 a_3505_10933 a_4420_11305 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4916 a_16276_19087 tdc1.r_dly_store_ring2 a_16055_19414 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X4917 VPWR tdc1.w_ring_buf31 a_27689_20009 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4918 tdc1.w_ring_int_norsz14 net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4919 a_8933_20725 a_8767_20725 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4922 VPWR tdc1.r_dly_store_ctr4 a_23201_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X4924 net21 a_9004_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4925 a_13948_16911 _116_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4926 a_28135_16586 tdc1.w_ring_norsz11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4927 a_12391_21629 a_11527_21263 a_12134_21375 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4929 a_13732_21039 _131_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4931 _055_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4932 a_20717_13897 tdc1.r_dly_store_ctr8 a_20635_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4933 _044_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4934 VPWR a_21223_15101 a_21391_15003 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4935 VGND net19 tdc0.w_ring_norsz15 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4936 a_11950_19605 a_11782_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X4937 tdc0.r_ring_ctr13 a_4595_14709 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X4939 _034_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4940 a_4203_16189 a_3505_15823 a_3946_15935 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X4942 a_12061_21629 a_11527_21263 a_11966_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4943 VPWR a_9931_11445 a_9918_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4944 a_29457_13103 _168_ _024_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4945 tdc0.r_dly_store_ring11 a_9155_15253 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4947 a_14793_11293 _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X4948 tdc0.w_ring_int_norsz24 tdc0.w_ring_norsz23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4949 VPWR a_18383_17076 tdc1.w_ring_buf20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4950 a_16439_15101 a_15575_14735 a_16182_14847 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X4951 a_24725_10383 a_24681_10625 a_24559_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X4952 net20 a_4443_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
R71 VGND net68 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4954 VGND _107_ a_22293_15395 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4955 a_12875_20327 tdc0.r_dly_store_ring22 a_13049_20203 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4956 VPWR a_21164_12559 a_21339_12533 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4957 a_19165_16911 _083_ a_18731_17063 VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4958 VGND a_25571_12319 a_25505_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X4959 VPWR net6 a_25971_18551 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X4961 VPWR a_22311_11989 a_22227_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4962 a_14791_17821 tdc0.r_dly_store_ring4 a_14428_17687 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X4964 _114_ a_12723_17161 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4965 a_20316_18151 _125_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4966 tdc0.w_ring_norsz30 net19 a_6461_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4967 VGND tdc1.w_ring_norsz9 tdc1.w_ring_norsz25 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4969 tdc1.w_ring_buf9 a_20727_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4970 VPWR tdc0.w_dly_stop4 a_3707_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X4971 tdc0.w_ring_buf9 a_14195_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4972 a_27251_13077 a_27095_13345 a_27396_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X4974 VPWR _079_ a_14545_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X4975 a_8113_16073 net39 tdc0.w_ring_int_norsz12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4976 tdc0.w_ring_buf2 a_11067_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4978 tdc1.w_ring_int_norsz16 net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4979 VPWR a_10275_15101 a_10443_15003 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X4980 VGND _197_ _039_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4982 VGND a_24887_15003 a_24845_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X4983 VGND tdc0.w_ring_norsz14 a_6283_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X4984 a_3707_12559 tdc0.r_ring_ctr10 a_3601_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4985 a_22687_17277 a_21905_16911 a_22603_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X4986 a_30005_17455 tdc1.w_ring_buf30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X4987 VPWR a_17987_17429 a_17903_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X4988 VPWR a_5791_12533 _162_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.165 ps=1.33 w=1 l=0.15
X4989 a_17924_17063 _111_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4991 a_21813_18543 a_21279_18549 a_21718_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4993 a_11969_19453 a_11435_19087 a_11874_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4995 a_27182_13103 a_27056_13219 a_26778_13235 VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X4996 VGND tdc1.w_ring_norsz17 tdc1.w_ring_int_norsz18 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4997 a_1297_16367 tdc0.r_ring_ctr15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4998 VPWR a_26627_18543 a_26747_18863 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4999 a_9071_15279 a_8289_15285 a_8987_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5000 a_14917_20719 tdc0.w_ring_buf1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5001 VGND net18 tdc1.w_ring_norsz1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5002 a_2374_14191 a_1297_14197 a_2212_14569 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5003 a_20713_14735 tdc1.w_ring_buf8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5004 a_11049_14735 a_10883_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5005 tdc0.w_ring_int_norsz22 net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5007 VGND a_11103_16189 a_11271_16091 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5008 a_24221_18909 tdc0.r_dly_store_ring30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.103 ps=1 w=0.42 l=0.15
X5009 VPWR net31 a_13551_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5010 tdc0.w_ring_int_norsz3 net39 a_10613_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5011 a_11839_15279 a_10975_15285 a_11582_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5013 VGND a_18751_21415 tdc1.r_dly_store_ring1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5014 VGND a_12594_12671 a_12552_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5015 a_24309_18909 _064_ a_24221_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X5016 a_12134_21375 a_11966_21629 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5017 _194_ a_20911_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X5018 a_22363_10749 _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5019 tdc1.w_ring_int_norsz27 net74 a_26805_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5021 VPWR tdc1.r_dly_store_ring30 a_18877_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X5022 VPWR a_28915_10927 _198_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R72 VGND net75 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5024 VPWR a_12134_21375 a_12061_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5025 a_26686_12147 a_26964_12131 a_26920_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X5026 a_13717_14985 tdc0.r_dly_store_ring16 a_13633_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5027 a_9839_17715 net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X5028 net31 a_16180_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5031 tdc1.w_ring_int_norsz26 tdc1.w_ring_norsz25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5032 VGND a_22615_16599 _105_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X5033 VPWR _071_ a_12989_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5034 VGND a_23907_21237 net35 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5037 VGND tdc1.r_ring_ctr1 a_28977_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5038 VGND tdc0.w_ring_norsz15 a_5087_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5039 a_26755_19863 a_26851_19863 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5041 a_25203_10357 _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5044 VGND net30 a_14195_13109 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5046 VPWR _069_ a_13633_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5049 a_20349_17455 net41 tdc1.w_ring_int_norsz4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5051 VGND a_5694_17023 a_5652_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5052 a_5951_17277 a_5087_16911 a_5694_17023 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5053 VPWR a_24551_11623 _029_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X5055 a_12332_10217 a_11417_9845 a_11985_9813 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5056 VGND _087_ a_20568_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X5057 a_27053_13469 a_26575_13077 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X5058 VPWR a_2571_15797 a_2558_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5059 _071_ a_24275_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5062 VGND net21 tdc0.w_ring_norsz2 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5064 tdc0.w_ring_buf16 a_5363_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5066 VGND net30 a_16127_14197 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5067 a_11414_15279 a_11141_15285 a_11329_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5068 a_24819_17776 _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5069 VPWR ui_in[1] a_29559_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5070 a_22917_19637 a_22751_19637 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5072 _122_ a_27517_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X5073 VGND a_23542_17429 a_23500_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5074 a_6725_13109 a_6559_13109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5075 VPWR a_21886_18517 a_21813_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5077 a_12851_12925 a_11987_12559 a_12594_12671 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5078 VGND net31 a_11343_19637 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5080 a_22457_19087 a_22291_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5081 a_11950_13759 a_11782_14013 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5082 a_10129_20175 a_9963_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5083 a_11540_12393 a_11141_12021 a_11414_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5084 VGND a_10667_10357 a_10601_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5085 a_23542_10901 a_23374_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5086 a_19860_15797 _071_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5087 VGND tdc0.r_ring_ctr2 _144_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5088 a_16937_11471 a_16771_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5089 VGND a_16658_15279 a_16764_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5090 VGND a_22603_17277 a_22771_17179 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5091 VPWR _147_ a_9025_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5092 VPWR net31 a_14287_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5093 tdc1.r_ring_ctr10 a_22995_10357 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X5094 tdc1.w_ring_buf14 a_29743_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5095 VGND tdc1.w_ring_norsz24 a_18979_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5096 a_4621_13481 a_3431_13109 a_4512_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5097 a_15128_20009 a_14729_19637 a_15002_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5099 a_23374_10927 a_23101_10933 a_23289_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5100 a_29785_12381 a_29741_11989 a_29619_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5101 a_6388_14569 a_5989_14197 a_6262_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5102 a_24275_16885 _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.146 ps=1.34 w=0.42 l=0.15
X5103 tdc1.w_ring_norsz2 tdc1.w_ring_norsz18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5107 tdc1.w_ring_buf24 a_18979_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5108 VPWR tdc0.w_ring_buf0 a_9503_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5109 VGND tdc1.w_ring_int_norsz28 tdc1.w_ring_norsz28 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5110 net22 a_6796_17973 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X5112 a_22730_19453 a_22291_19087 a_22645_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5113 tdc0.r_ring_ctr8 a_4595_11231 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X5114 a_22907_12559 _183_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X5115 VGND tdc1.r_ring_ctr13 a_18141_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5116 VGND net16 _063_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5117 net41 a_26031_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5118 tdc0.r_ring_ctr14 a_2571_15797 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X5119 VPWR _197_ _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5120 tdc0.w_ring_norsz20 tdc0.w_ring_int_norsz20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5121 a_17225_14735 tdc0.r_dly_store_ring0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X5122 a_25137_10383 a_23947_10383 a_25028_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5123 VGND _040_ a_4117_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5124 tdc0.r_dly_store_ring6 a_9799_20693 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5127 a_9096_11471 _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5128 _083_ a_16187_19891 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5129 tdc0.w_ring_int_norsz0 net61 a_3897_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5130 a_6841_11471 _147_ a_6769_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5131 a_19142_12015 a_18703_12021 a_19057_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5132 VGND net3 a_12723_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5133 VGND a_2387_13407 a_2321_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5134 tdc1.w_ring_buf27 a_26983_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5135 VPWR tdc1.w_ring_int_norsz31 a_28253_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5137 VPWR a_29519_14165 _170_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5138 VPWR a_20119_14191 a_20287_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5139 a_24087_18775 _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.128 ps=1.03 w=0.42 l=0.15
X5140 VGND _042_ a_1909_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5141 VGND tdc1.w_ring_int_norsz17 tdc1.w_ring_norsz17 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5143 VPWR a_3483_14423 _004_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5145 a_19785_16745 a_18795_16373 a_19659_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5146 a_29057_21428 ui_in[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5147 a_23907_21237 net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X5149 VGND tdc0.w_dly_stop4 a_3707_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5150 a_3601_16911 tdc0.r_ring_ctr15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5151 a_23699_19631 a_22917_19637 a_23615_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5152 a_25049_13889 a_24831_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5153 a_22351_13321 net33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5155 a_6983_10383 a_6633_10383 a_6888_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5157 _075_ a_15451_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5158 a_19835_15279 a_19053_15285 a_19751_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5159 _197_ a_5087_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5160 VGND a_9374_20693 a_9332_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5161 tdc0.w_ring_buf2 a_11067_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5162 _060_ net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5164 _069_ a_14623_16627 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5165 a_18155_17161 _110_ a_18059_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X5167 _121_ a_26747_18863 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X5168 tdc1.w_ring_norsz10 tdc1.w_ring_int_norsz10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5169 a_20813_18543 tdc1.w_ring_norsz25 a_20729_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5170 VPWR _170_ a_26689_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5171 tdc0.w_ring_int_norsz31 net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5173 VGND a_7815_11623 _150_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5174 a_29723_12925 _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5175 VGND a_16187_19891 _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X5176 a_20051_10357 _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5177 VGND a_18383_17076 tdc1.w_ring_buf20 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5179 tdc0.w_ring_norsz17 net20 a_5357_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5180 a_17861_13103 tdc1.r_ring_ctr14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5181 VPWR a_6062_14847 a_5989_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5182 VGND a_11747_18365 a_11915_18267 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5184 VGND a_21463_15823 _089_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5187 _028_ _176_ a_25425_12809 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5188 a_12079_16073 _080_ a_12161_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5189 uo_out[5] a_14372_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X5191 VGND _077_ a_15577_16483 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5192 a_13069_16911 tdc0.r_dly_store_ctr4 a_12723_17161 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5193 VPWR a_14899_10143 a_14886_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5194 a_19529_10625 a_19311_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5195 VGND net8 a_8675_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5196 VPWR a_11547_12827 a_11463_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5197 VPWR a_27871_16885 a_27878_17185 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5199 VPWR tdc1.w_ring_int_norsz6 a_17857_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5201 _003_ _162_ a_1113_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X5202 VPWR a_18021_15797 _109_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5203 tdc0.r_dly_store_ctr12 a_4555_16341 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5204 a_16842_16367 a_16569_16373 a_16757_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
R73 tdc1.g_ring323.stg01_70.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5205 a_28687_21085 a_28467_21097 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X5206 a_7607_20541 a_6909_20175 a_7350_20287 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5207 VGND a_11950_13759 a_11908_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5208 uo_out[7] a_14172_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5209 a_20119_14191 a_19255_14197 a_19862_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5210 _008_ _144_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5211 a_4905_17455 tdc0.w_ring_int_norsz1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5213 a_5161_15823 a_4995_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5214 a_24701_14191 a_24363_14423 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5216 a_29173_12021 a_29007_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5217 a_30423_18365 a_29559_17999 a_30166_18111 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5218 a_9279_21237 net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X5219 a_14560_20425 _142_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X5220 a_24251_19863 tdc1.r_dly_store_ring10 a_24397_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5221 a_27249_20719 net17 tdc1.w_ring_norsz16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5227 a_17500_12335 _185_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5228 a_17286_12559 _062_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5229 _155_ a_5271_12128 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
R74 VPWR tdc1.g_ring116.stg02_62.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5230 VGND net15 tdc1.w_ring_norsz19 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5231 a_17417_12015 tdc1.r_ring_ctr12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X5232 a_18869_12021 a_18703_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5233 a_30093_18365 a_29559_17999 a_29998_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5234 tdc1.w_ring_int_norsz1 net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5235 VGND tdc1.w_ring_norsz27 tdc1.w_ring_int_norsz28 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5236 a_27595_11471 a_27149_11471 a_27499_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5237 a_12897_17455 tdc0.r_dly_store_ctr7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5238 a_6587_14013 a_5805_13647 a_6503_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5241 a_4866_13469 _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5242 _032_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5243 a_21905_10383 a_21739_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5244 a_28529_12335 tdc1.r_ring_ctr1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5245 a_30166_18111 a_29998_18365 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5246 VPWR a_30683_17429 a_30599_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5247 a_10023_10383 a_9577_10383 a_9927_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5248 a_4471_16367 a_3689_16373 a_4387_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5250 a_14865_11293 a_14486_10927 a_14793_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X5252 VGND tdc1.w_ring_norsz23 tdc1.w_ring_norsz7 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5253 a_21633_18543 tdc1.w_ring_buf21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5254 a_7548_10383 a_6467_10383 a_7201_10625 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5255 VGND _056_ a_24725_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5256 a_27722_10927 a_26964_11043 a_27159_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X5257 a_11425_17455 net43 tdc0.w_ring_int_norsz2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5258 a_28289_20719 a_27951_20951 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5260 VGND tdc1.r_dly_store_ring20 a_18337_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5262 a_26778_13235 a_27095_13345 a_27053_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X5263 a_23201_16073 _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5264 a_11517_14191 net39 tdc0.w_ring_int_norsz9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5265 tdc1.w_ring_buf14 a_29743_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5266 tdc0.r_dly_store_ctr5 a_12007_11989 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5267 VGND net28 a_6559_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5268 tdc0.r_dly_store_ring5 a_12467_19355 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5270 tdc0.r_dly_store_ctr5 a_12007_11989 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5271 a_12907_16367 _072_ a_12989_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5272 a_24685_19951 net24 a_24251_19863 VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5273 tdc1.w_ring_norsz21 net14 a_18881_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5274 a_10773_19337 tdc0.w_ring_norsz24 a_10689_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5275 VGND a_17107_12533 a_17041_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5276 VPWR a_27095_13345 a_27056_13219 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5277 VPWR tdc0.w_ring_norsz11 a_8113_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5278 a_18233_18543 net41 tdc1.w_ring_int_norsz6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5279 VPWR tdc1.w_ring_int_norsz18 a_21445_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5280 VPWR tdc1.r_dly_store_ring0 a_20911_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5281 a_26439_14191 _170_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5282 VPWR a_27772_16341 net17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5283 a_27894_14709 a_27694_15009 a_28043_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5284 a_18961_16373 a_18795_16373 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5285 a_13551_15279 _075_ a_13633_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5286 a_20924_14735 a_20525_14735 a_20798_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5287 a_4165_13077 a_3947_13481 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5288 VPWR a_27259_19087 _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5289 a_15128_12393 a_14729_12021 a_15002_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5290 VPWR a_23075_18762 tdc1.w_ring_buf10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5293 _125_ a_20258_16073 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X5294 _023_ a_28279_12015 a_28529_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X5295 VPWR _069_ a_20717_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5296 VPWR tdc1.r_dly_store_ring14 a_19065_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5298 a_26426_17687 tdc1.r_dly_store_ring11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.172 ps=1.46 w=0.42 l=0.15
X5300 a_22898_19199 a_22730_19453 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5302 VGND a_19860_15797 _080_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5303 a_17596_20425 _078_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5304 tdc1.r_dly_store_ring6 a_18723_19605 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5305 a_22558_13380 a_22358_13225 a_22707_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5306 net23 a_7111_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X5308 VGND a_7166_13077 a_7124_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5309 a_24736_12381 _029_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5310 VGND _076_ a_13827_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5313 tdc1.r_dly_store_ring6 a_18723_19605 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5314 VPWR a_30166_18111 a_30093_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5315 VPWR tdc1.w_ring_norsz16 a_25787_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5316 a_25849_15657 a_25302_15401 a_25502_15556 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X5317 VPWR tdc1.w_ring_norsz3 a_20911_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5318 VGND net27 a_8767_20725 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5319 a_30088_12393 a_29007_12021 a_29741_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5321 VGND net14 tdc1.w_ring_norsz20 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5322 a_5767_19453 a_5069_19087 a_5510_19199 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5325 a_8086_17429 a_7918_17455 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5327 a_13161_15823 tdc0.r_dly_store_ctr5 a_12723_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5328 VPWR _034_ a_13879_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5330 VPWR a_7548_10383 a_7723_10357 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5332 VPWR a_25502_15556 a_25431_15657 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5336 VPWR tdc1.w_ring_buf0 a_26615_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5338 net24 a_27403_17973 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5339 VGND _076_ a_13732_21039 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5340 a_7166_13077 a_6998_13103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5341 a_24831_13647 a_24481_13647 a_24736_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5342 a_22178_21629 a_21739_21263 a_22093_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5343 VPWR a_8987_15279 a_9155_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5344 a_9263_17277 a_8565_16911 a_9006_17023 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5347 a_29642_15797 a_29442_16097 a_29791_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5348 a_11153_19337 tdc0.w_ring_norsz8 a_11069_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5349 a_4866_12381 _041_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5350 a_9918_11837 a_8841_11471 a_9756_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5351 a_10954_12925 a_10515_12559 a_10869_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5352 VGND a_8987_15279 a_9155_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5353 VPWR net33 a_21463_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5354 VPWR a_11763_11445 _147_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5356 VPWR net7 a_1131_13109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5358 a_29428_12381 _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5359 _093_ a_13551_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5360 a_7182_20541 a_6909_20175 a_7097_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5361 VGND a_13323_11159 _145_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X5362 a_4512_13481 a_3597_13109 a_4165_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5363 VGND tdc1.w_ring_norsz2 tdc1.w_ring_int_norsz3 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5364 VGND a_2387_14495 tdc0.r_ring_ctr12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5365 a_24113_10383 a_23947_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5366 a_13049_20203 _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X5367 a_9485_18543 tdc0.w_ring_norsz21 a_9401_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5368 a_21339_12533 _063_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5369 _031_ a_25623_11247 a_25861_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5370 a_19860_15797 _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5371 a_13732_21039 _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5372 tdc0.w_ring_norsz0 net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5373 tdc1.r_dly_store_ring26 a_25163_16091 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5374 a_14821_19453 a_14287_19087 a_14726_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5375 a_1843_15645 tdc0.r_ring_ctr14 a_1747_15645 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X5377 a_13344_20693 _134_ a_13732_21039 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5378 VGND tdc1.w_ring_buf29 a_30725_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5381 VGND a_17895_13915 a_17853_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5382 a_22638_14013 a_22199_13647 a_22553_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5383 VGND tdc1.w_ring_norsz1 a_18887_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5384 a_12618_21039 _128_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.117 ps=1.01 w=0.65 l=0.15
X5386 VGND a_19827_16341 a_19785_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5389 a_13671_13103 a_12889_13109 a_13587_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5390 a_19421_17455 tdc1.w_ring_norsz4 a_19337_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5391 a_13633_15279 tdc0.r_dly_store_ring26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5392 a_22255_10383 a_21905_10383 a_22160_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5393 VPWR tdc0.w_ring_norsz19 a_9309_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5394 VPWR _147_ a_7815_11623 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5395 VGND _049_ a_29785_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5396 VGND _104_ a_22615_16599 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X5398 a_16569_16373 a_16403_16373 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5400 VGND net26 a_9411_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5401 VGND tdc1.r_ring_ctr4 a_25297_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X5402 a_30534_15253 a_30366_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5403 a_3505_10933 a_3339_10933 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5405 VPWR a_4595_14709 a_4582_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5406 a_3571_19252 tdc0.w_dly_stop2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5407 VPWR tdc0.r_ring_ctr6 a_6987_12247 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5409 VPWR a_9409_11713 a_9299_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5410 a_1389_16911 a_1223_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5411 VPWR _075_ a_13625_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X5412 a_17047_14735 _089_ a_17225_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5414 a_19862_14165 a_19694_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5415 a_30366_15279 a_30093_15285 a_30281_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
R75 VPWR tt_um_hpretl_tt06_tdc_v2_80.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5417 VGND a_21971_13335 tdc1.r_dly_store_ctr6 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5418 a_16566_14191 a_16127_14197 a_16481_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5419 a_9301_16189 a_8767_15823 a_9206_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5420 VPWR tdc1.w_ring_norsz18 a_20993_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5421 tdc1.r_ring_ctr14 a_17107_12533 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X5422 a_22256_20425 _085_ a_21791_20327 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X5423 tdc1.r_dly_store_ring5 a_19827_16341 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5424 VPWR a_25163_16091 a_25079_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5425 a_2227_15279 tdc0.r_ring_ctr14 _166_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.27 ps=2.54 w=1 l=0.15
X5426 VGND a_28331_20937 a_28338_20841 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5427 a_26755_15975 a_26851_15797 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5428 a_10425_17455 tdc0.w_ring_int_norsz18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5429 VGND a_17987_17429 a_17945_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5430 a_19694_14191 a_19421_14197 a_19609_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5431 tdc1.r_dly_store_ring5 a_19827_16341 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5432 VPWR a_13735_21263 _076_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5433 VPWR a_16727_20951 tdc1.r_dly_store_ring7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5435 _101_ a_13091_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5436 VGND tdc0.w_dly_stop5 a_4443_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X5437 VPWR a_17567_10099 net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X5438 VPWR a_4279_17179 a_4195_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5441 a_14399_11169 net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5442 tdc0.r_dly_store_ring14 a_7775_20443 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5443 VGND a_26755_19863 tdc1.r_dly_store_ring31 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5444 a_25396_13647 a_24315_13647 a_25049_13889 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X5445 a_23289_17455 tdc1.w_ring_buf25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5446 VGND a_24462_14847 a_24420_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5447 tdc0.w_ring_norsz1 net19 a_4989_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5449 a_3946_15935 a_3778_16189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5451 a_27396_13103 a_27182_13103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X5452 VGND net33 a_19255_14197 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5453 a_7245_10383 a_7201_10625 a_7079_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5454 tdc0.r_dly_store_ring27 a_8603_14165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5455 _100_ a_16055_19414 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.113 ps=1.04 w=0.65 l=0.15
X5456 a_13817_14191 tdc0.r_dly_store_ctr2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X5457 VPWR net31 a_14563_20725 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5458 a_2558_16189 a_1481_15823 a_2396_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5459 _627_.X a_29467_15287 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5460 a_2322_15599 tdc0.r_ring_ctr12 _166_ VGND sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.106 ps=0.975 w=0.65 l=0.15
X5461 VGND a_19310_11989 a_19268_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5462 VPWR a_14894_19199 a_14821_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5463 VPWR _170_ a_22711_12533 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X5465 VPWR a_15227_13077 a_15143_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5466 VGND a_27342_19908 a_27271_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5467 VGND tdc0.w_ring_int_norsz14 tdc0.w_ring_norsz14 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5468 a_4595_11231 a_4420_11305 a_4774_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5469 VGND a_23075_18762 tdc1.w_ring_buf10 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5470 VPWR tdc1.r_ring_ctr8 a_23485_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5471 a_4111_17277 a_3413_16911 a_3854_17023 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5472 a_24591_12559 _170_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5473 a_19494_15253 a_19326_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5475 a_24551_11623 a_24694_11517 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X5476 a_16055_19414 tdc0.r_dly_store_ring2 a_16055_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5477 VPWR tdc1.w_ring_norsz29 a_30295_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5478 a_26897_17161 tdc1.w_ring_norsz10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5479 VGND a_19862_14165 a_19820_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5482 a_19721_18543 tdc1.w_ring_norsz24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5484 a_18256_20009 a_17857_19637 a_18130_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5485 a_30366_15279 a_29927_15285 a_30281_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5486 VGND net14 tdc1.w_ring_norsz5 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5487 VPWR a_14555_10901 a_14486_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X5488 VPWR net30 a_16219_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X5489 a_27070_19997 a_26755_19863 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X5490 a_7718_18517 a_7550_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5491 a_24803_15101 a_24021_14735 a_24719_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5493 a_15094_14013 a_14655_13647 a_15009_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5494 a_23264_21237 net35 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5495 a_5342_19453 a_5069_19087 a_5257_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5497 a_25601_18903 net4 a_25520_18903 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X5499 VGND a_15595_11989 a_15553_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5500 a_19728_11471 a_19329_11471 a_19602_11837 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5501 a_29612_13647 _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5502 VPWR a_12375_19605 a_12291_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5503 VGND net23 tdc0.w_ring_norsz9 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5504 VPWR _172_ a_24591_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5505 a_21445_12021 a_21279_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5506 a_12161_15823 tdc0.r_dly_store_ctr13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5507 VPWR _086_ a_22741_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X5508 tdc1.r_dly_store_ctr8 a_20195_11739 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5509 VGND _072_ a_13161_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X5510 a_25509_17571 net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.148 ps=1.34 w=0.42 l=0.15
X5511 a_7645_17461 a_7479_17461 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5512 a_28467_21097 a_28338_20841 a_28047_20951 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5513 a_25892_19951 net6 a_25221_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X5514 tdc1.w_ring_int_norsz9 tdc1.w_ring_norsz8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5515 tdc0.r_dly_store_ring6 a_9799_20693 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5517 VGND a_17435_16341 a_17393_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5518 VGND net15 tdc1.w_ring_norsz3 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5519 a_27491_17063 a_27587_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5520 tdc1.w_ring_int_norsz17 net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5521 a_1755_13103 _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5522 a_10954_12925 a_10681_12559 a_10869_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5523 VPWR net26 a_9411_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5524 VGND net7 a_5823_10933 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5525 a_21445_19637 a_21279_19637 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5527 a_27003_12257 net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5528 VPWR tdc0.r_ring_ctr4 a_8857_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5529 a_24201_15599 tdc1.r_dly_store_ctr7 a_23855_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5530 a_28823_14557 tdc1.r_ring_ctr2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5531 VPWR a_9374_15935 a_9301_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5532 VGND _067_ _072_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5533 a_30534_14165 a_30366_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5534 a_7699_12925 a_7001_12559 a_7442_12671 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5536 _016_ tdc1.r_ring_ctr0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5537 a_7274_12925 a_6835_12559 a_7189_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5538 a_19705_17455 net14 tdc1.w_ring_norsz4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5541 VGND tdc0.r_ring_ctr12 a_863_13897 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5542 VGND tdc1.r_dly_store_ctr9 a_22753_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X5543 VPWR a_25396_13647 a_25571_13621 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
R76 VPWR tdc0.g_ring324.stg01_53.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5545 tdc1.r_ring_ctr11 a_20051_10357 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X5546 _115_ a_12723_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5547 a_30366_14191 a_30093_14197 a_30281_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5548 a_13543_17571 _115_ a_13461_17571 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5549 a_12867_15511 tdc0.r_dly_store_ctr6 a_12993_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X5551 tdc0.r_dly_store_ctr14 a_4371_16091 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5552 a_23799_10927 a_23101_10933 a_23542_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5553 a_18045_19631 tdc1.w_ring_buf6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5554 _170_ a_29519_14165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5555 VPWR tdc1.w_dly_stop5 a_29467_15287 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X5556 a_23374_10927 a_22935_10933 a_23289_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5557 VPWR tdc0.w_ring_norsz13 a_6089_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5559 tdc1.w_ring_norsz17 tdc1.w_ring_norsz1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5560 a_5809_14735 tdc0.w_ring_buf16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5561 a_28135_16586 tdc1.w_ring_norsz11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5562 _075_ a_15451_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5563 a_2658_16911 _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5565 tdc0.r_dly_store_ring24 a_12375_13915 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5566 VPWR a_12507_10143 tdc0.r_ring_ctr0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X5568 a_6983_10383 a_6467_10383 a_6888_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5569 tdc1.r_dly_store_ctr15 a_23231_13915 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5570 a_12425_19087 a_11435_19087 a_12299_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5572 a_7423_19631 a_6725_19637 a_7166_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5573 a_11490_18111 a_11322_18365 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5574 a_2425_15599 tdc0.r_ring_ctr13 a_2322_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X5575 a_18751_21415 a_18847_21237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5576 tdc0.w_ring_norsz20 net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5578 a_3760_11293 _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5579 VGND _092_ a_15117_14741 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5582 a_12092_21263 a_11693_21263 a_11966_21629 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X5585 a_13827_15823 _089_ a_14005_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5586 a_1481_15823 a_1315_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5587 a_14899_10143 _033_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5588 VGND a_9647_15253 net26 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5589 VGND a_16187_19891 _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5590 a_15078_10205 _033_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5592 VPWR net12 a_11425_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5593 a_20729_18543 tdc1.w_ring_int_norsz9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5594 VPWR a_29791_18775 tdc1.r_dly_store_ring29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5595 tdc1.w_ring_norsz14 tdc1.w_ring_int_norsz14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5596 VPWR a_4687_12319 a_4674_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5597 VPWR net11 a_11517_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5598 _192_ a_17047_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5599 tdc0.w_ring_buf9 a_14195_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5601 a_26689_14191 tdc1.r_ring_ctr4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R77 VPWR tdc1.g_ring318.stg01_65.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5602 tdc0.w_ring_norsz27 tdc0.w_ring_int_norsz27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5603 a_25441_19631 net6 _087_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.153 ps=1.3 w=1 l=0.15
X5604 VPWR a_6904_11305 a_7079_11231 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5606 a_5357_17455 tdc0.w_ring_norsz1 a_5273_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5607 tdc0.r_dly_store_ring15 a_5935_19355 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5608 VPWR a_22820_10383 a_22995_10357 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5611 VPWR tdc1.w_ring_buf4 a_16097_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X5612 a_3413_16911 a_3247_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5613 _089_ a_21463_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5614 a_13817_14511 tdc0.r_dly_store_ctr10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5615 a_4909_18249 tdc0.w_ring_norsz0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5616 VGND net30 a_16219_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5617 VPWR tdc1.w_dly_stop1 a_15575_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5619 VGND tdc0.w_ring_int_norsz12 tdc0.w_ring_norsz12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5620 a_15259_16885 a_15543_16885 a_15478_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X5621 VPWR a_4387_16367 a_4555_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5622 a_13195_15279 tdc0.r_dly_store_ctr14 a_12993_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5623 VPWR a_4371_16091 a_4287_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
R78 uio_out[5] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5624 a_23264_21237 net35 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5625 a_24673_12559 tdc1.r_ring_ctr6 a_24591_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5626 a_19216_10383 _018_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
R79 tdc1.g_ring331.stg01_78.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5629 a_17857_19337 tdc1.w_ring_norsz22 a_17773_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5631 VGND a_4387_16367 a_4555_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5633 a_27182_13103 a_27095_13345 a_26778_13235 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X5635 a_8933_15823 a_8767_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5636 tdc1.w_ring_norsz11 net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5637 a_15715_17674 tdc1.w_ring_norsz4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5638 net16 a_17567_10099 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5639 VGND tdc0.w_ring_norsz10 tdc0.w_ring_int_norsz11 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5640 VPWR a_25049_11989 a_24939_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5641 VPWR a_14172_20149 uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5642 a_27149_11471 a_26983_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5645 tdc1.w_dly_stop5 a_16587_10927 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5646 a_4774_14735 _045_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5647 VPWR a_17647_18762 tdc1.w_ring_buf22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X5648 VGND a_28047_21237 net43 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5649 VGND net26 a_4995_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5650 a_19326_15279 a_19053_15285 a_19241_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5652 VPWR _177_ a_22199_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5653 a_17647_18762 tdc1.w_ring_norsz22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5654 a_9577_10383 a_9411_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5656 a_27607_11837 a_26983_11471 a_27499_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5657 VPWR net9 a_29007_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5658 VPWR _067_ a_27351_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5659 a_24397_19631 net24 a_24251_19863 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X5661 a_17044_17161 _100_ a_16656_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5662 a_9631_20719 a_8767_20725 a_9374_20693 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5663 VGND a_1551_15253 _165_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X5664 a_29883_21428 ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5665 VPWR _057_ a_27304_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X5667 a_19605_13103 tdc1.r_ring_ctr15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5668 _072_ a_24635_17973 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5669 a_22227_18543 a_21445_18549 a_22143_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5672 a_20695_12559 a_20249_12559 a_20599_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5673 a_18961_10383 a_18795_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5677 VPWR a_23967_10901 a_23883_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5678 a_9953_14191 net23 tdc0.w_ring_norsz10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5679 a_21729_16687 tdc1.r_dly_store_ring19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5680 a_5529_16189 a_4995_15823 a_5434_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5681 tdc0.w_ring_norsz7 net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5682 a_6837_17455 tdc0.w_ring_int_norsz29 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5683 a_16155_15975 tdc0.r_dly_store_ring25 a_16301_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5684 a_16182_14847 a_16014_15101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5685 a_14641_19087 tdc0.w_ring_buf2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5686 a_24995_16189 a_24297_15823 a_24738_15935 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5687 a_5261_12559 _156_ _161_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5688 tdc0.r_dly_store_ctr11 a_6855_14165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5689 a_1552_14557 _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5690 VGND a_25839_16341 net25 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5694 a_11877_14013 a_11343_13647 a_11782_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5695 a_4387_16367 a_3523_16373 a_4130_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5696 a_26893_20719 tdc1.w_ring_int_norsz16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5697 _106_ a_21647_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5698 VGND net5 a_25892_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5699 tdc1.w_ring_norsz7 tdc1.w_ring_int_norsz7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5700 VGND net38 a_29099_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X5702 VGND a_28279_12015 _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X5704 a_3686_17277 a_3247_16911 a_3601_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5705 VGND _008_ a_15118_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X5707 a_4057_16367 a_3523_16373 a_3962_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5709 a_13717_17999 a_13551_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5710 VPWR a_14123_11989 a_14039_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5711 VPWR a_11839_12015 a_12007_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5712 VGND ui_in[1] a_29559_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5714 a_7277_18549 a_7111_18549 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5715 VGND a_12299_19453 a_12467_19355 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5716 a_23259_18164 tdc1.w_ring_norsz25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5718 a_17192_11471 _020_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5719 VGND a_11839_12015 a_12007_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5720 VPWR net35 a_22199_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5721 VGND net34 a_22291_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5722 a_7274_12925 a_7001_12559 a_7189_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5723 a_10689_19337 net22 tdc0.w_ring_norsz8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5724 _030_ _179_ a_23653_10159 VGND sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X5725 a_7925_14191 tdc0.w_ring_buf27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5726 a_26111_20938 tdc1.w_ring_norsz16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5727 tdc0.w_ring_buf16 a_5363_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5728 VGND a_24467_16599 _096_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5729 _084_ net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5730 VPWR _154_ a_5791_12533 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X5731 a_2750_15823 _046_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5732 a_24275_16885 a_24631_16891 a_24589_16917 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5733 VPWR net34 a_18795_16373 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5734 tdc0.w_ring_buf17 a_4811_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5735 VGND a_12375_19605 a_12333_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5736 a_15271_14985 _093_ a_15199_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5737 a_12762_20719 _127_ a_12448_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.28 ps=1.56 w=1 l=0.15
X5738 a_16269_19414 tdc0.r_dly_store_ring2 a_16055_19414 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.193 ps=1.34 w=0.42 l=0.15
X5739 a_13625_18543 tdc0.r_dly_store_ring5 a_13541_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5741 a_15027_15823 _108_ a_15196_16073 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5742 VGND a_26667_21237 net5 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X5744 a_6035_17277 a_5253_16911 a_5951_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5745 a_9409_11713 a_9191_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5747 _103_ a_13827_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5750 VGND tdc0.w_ring_norsz7 tdc0.w_ring_int_norsz8 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5751 a_7423_19631 a_6559_19637 a_7166_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5752 a_23489_15823 _075_ a_23055_15975 VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5753 VPWR tdc1.w_ring_int_norsz29 a_28713_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5754 VPWR tdc1.w_ring_norsz23 a_20533_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5755 VPWR net29 a_12723_13109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5757 a_24433_13441 _170_ a_24347_13441 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5759 a_21997_11837 a_21463_11471 a_21902_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5761 a_25093_12381 a_25049_11989 a_24927_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5763 VGND _076_ a_16276_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
X5764 a_30791_16367 a_30093_16373 a_30534_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5765 VGND a_5875_11623 _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X5766 a_1552_14557 _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X5767 tdc0.r_dly_store_ring0 a_16607_15003 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5768 VPWR a_15750_16885 a_15679_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5769 net3 a_28415_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5770 a_7093_19631 a_6559_19637 a_6998_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5771 VPWR a_13587_13103 a_13755_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5773 VPWR net34 a_16955_17461 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5776 a_21633_12015 tdc1.r_ring_ctr11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5777 VGND a_13587_13103 a_13755_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5778 VGND a_8086_17429 a_8044_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5780 a_21905_21263 a_21739_21263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5781 a_24131_19337 _072_ a_24213_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5782 tdc1.w_ring_int_norsz20 net67 a_20089_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5784 tdc1.r_dly_store_ring3 a_22771_17179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5785 a_6998_19631 a_6559_19637 a_6913_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X5786 tdc0.r_ring_ctr15 a_2479_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X5787 VGND tdc0.w_ring_int_norsz9 tdc0.w_ring_norsz9 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5788 tdc1.w_ring_buf27 a_26983_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5789 a_4357_17455 tdc0.w_ring_norsz16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5790 VGND a_11582_11989 a_11540_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5791 a_16569_10383 a_16403_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5792 tdc0.w_ring_norsz23 net22 a_9773_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5793 VPWR tdc1.w_ring_int_norsz23 a_17489_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5795 a_11069_19337 tdc0.w_ring_int_norsz24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5797 a_24570_16189 a_24297_15823 a_24485_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5798 VPWR _172_ a_24347_13441 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5799 a_25932_12533 tdc1.w_ring_buf0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X5800 _159_ a_3431_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X5801 a_2953_10927 tdc0.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5803 VPWR a_24950_14468 a_24879_14569 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X5804 net14 a_18243_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5805 VGND a_16734_14165 a_16692_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5806 a_27135_15797 net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5807 a_3686_17277 a_3413_16911 a_3601_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5808 tdc1.w_ring_int_norsz15 net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5810 VGND net7 a_3431_13109 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5811 a_22569_14511 _080_ a_22135_14423 VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5812 a_15185_13481 a_14195_13109 a_15059_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5813 a_25861_11247 _180_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5814 a_12507_10143 _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5815 VGND tdc1.w_ring_norsz11 tdc1.w_ring_int_norsz12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5816 VGND net20 _046_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5817 a_22825_19453 a_22291_19087 a_22730_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5818 VGND a_12851_12925 a_13019_12827 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5819 a_14802_13077 a_14634_13103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5820 a_14729_19637 a_14563_19637 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5821 a_21886_19605 a_21718_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5822 tdc1.w_ring_int_norsz11 net41 a_26897_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5825 uo_out[3] a_15196_16073 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5826 tdc1.w_ring_int_norsz25 net72 a_19721_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5827 VGND a_17647_18762 tdc1.w_ring_buf22 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5828 a_27093_16189 a_26755_15975 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X5830 a_13732_21039 _134_ a_13344_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5831 a_11417_9845 a_11251_9845 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5832 a_20525_14735 a_20359_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5835 VPWR a_29925_13889 a_29815_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X5836 a_8895_13103 a_8031_13109 a_8638_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5837 tdc1.r_dly_store_ring2 a_15595_19605 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5838 a_27717_11713 a_27499_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X5839 a_14634_13103 a_14361_13109 a_14549_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5840 a_17647_18762 tdc1.w_ring_norsz22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5842 a_17562_17429 a_17394_17455 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5843 a_21353_10633 tdc1.r_ring_ctr10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5845 tdc0.r_dly_store_ring5 a_12467_19355 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5846 a_25287_18517 a_25643_18775 a_25601_18903 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5847 a_22255_10383 a_21739_10383 a_22160_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5848 tdc1.w_ring_buf13 a_29375_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X5851 a_13587_13103 a_12723_13109 a_13330_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5852 VGND _156_ a_3707_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X5853 uo_out[0] a_17804_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5854 VPWR a_29427_20693 net38 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5857 VPWR tdc0.r_ring_ctr9 a_2743_12711 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X5858 a_8565_13103 a_8031_13109 a_8470_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5859 tdc1.r_dly_store_ctr7 a_24887_15003 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5860 a_30378_18820 a_30178_18665 a_30527_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X5862 a_13265_19631 net3 a_13183_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5863 a_9466_12671 a_9298_12925 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5864 VGND a_5951_17277 a_6119_17179 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5865 a_13257_13103 a_12723_13109 a_13162_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5866 VGND tdc0.w_ring_norsz1 a_5455_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5868 a_17862_10927 _186_ a_17559_11159 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X5870 a_4329_15823 a_3339_15823 a_4203_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5871 VPWR a_7166_19605 a_7093_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5872 VGND a_30534_15253 a_30492_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5873 a_11782_19631 a_11509_19637 a_11697_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5874 a_28043_15511 a_28139_15511 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5876 a_29818_20541 a_29571_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5877 a_17777_11247 _187_ a_17559_11159 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5878 a_6503_14013 a_5805_13647 a_6246_13759 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X5879 VPWR a_22343_15975 _082_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
R80 uio_out[7] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5881 a_29925_13889 a_29707_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X5882 VPWR a_19131_21237 a_19138_21537 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5883 VPWR tdc1.w_ring_int_norsz0 a_26597_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5884 VPWR a_19659_16367 a_19827_16341 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X5885 VGND _162_ a_3788_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5887 a_10911_20541 a_10129_20175 a_10827_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5888 VGND a_26755_15975 tdc1.r_dly_store_ring27 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5889 a_5445_18543 net19 tdc0.w_ring_norsz31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5890 a_12889_18543 tdc0.r_dly_store_ring20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5893 _191_ a_13551_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X5894 tdc0.w_ring_norsz16 net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5895 a_7091_10749 _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X5896 VGND a_19659_16367 a_19827_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5898 a_10189_10383 a_10145_10625 a_10023_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X5899 a_10137_18543 net40 tdc0.w_ring_int_norsz5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5900 a_19141_14735 tdc1.r_dly_store_ctr6 a_18703_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5902 a_12805_16073 _118_ a_12723_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5903 VPWR a_14399_11169 a_14360_11043 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5905 a_8105_14191 a_7571_14197 a_8010_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5907 VGND tdc0.r_ring_ctr10 a_1317_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5908 VGND _145_ _008_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5909 VGND a_15196_16073 uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5910 a_9006_17023 a_8838_17277 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5911 VGND _162_ a_2425_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X5913 VGND a_30791_14191 a_30959_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5916 a_26721_11293 a_26686_11059 a_26483_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X5918 VPWR a_22898_19199 a_22825_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5920 a_23021_18249 tdc1.w_ring_norsz10 a_22937_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5921 VPWR net20 _042_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5922 VGND a_15163_17063 tdc1.r_dly_store_ring4 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5926 a_16014_15101 a_15741_14735 a_15929_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5929 tdc0.w_ring_norsz14 tdc0.w_ring_norsz30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5930 a_25382_10383 _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X5932 VPWR a_25287_18517 _068_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5933 VGND net7 a_3431_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5934 a_1647_13481 a_1297_13109 a_1552_13469 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5935 tdc0.w_ring_norsz22 net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5936 VGND a_26483_11989 tdc1.r_ring_ctr6 VGND sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X5937 VGND a_29642_15797 a_29571_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X5938 a_7091_10749 a_6467_10383 a_6983_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5939 a_9374_15935 a_9206_16189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5940 _108_ a_22293_15395 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X5941 VGND a_7591_16091 a_7549_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5942 a_30093_16373 a_29927_16373 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5943 VPWR net31 a_9963_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5946 tdc0.w_ring_norsz25 net23 a_10601_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5949 VPWR a_8638_13077 a_8565_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X5950 a_20525_14735 a_20359_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5951 a_15170_20693 a_15002_20719 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X5952 a_24719_15101 a_23855_14735 a_24462_14847 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X5953 a_24745_12559 _170_ a_24673_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X5955 _092_ a_14366_15599 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5957 VGND a_15319_19355 a_15277_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5959 VPWR a_7775_20443 a_7691_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X5960 tdc1.w_ring_norsz16 net17 a_26977_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5961 a_12447_14191 _080_ a_12529_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5963 a_24389_15101 a_23855_14735 a_24294_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X5964 VGND a_14158_18111 a_14116_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X5965 a_25221_19605 net6 a_25892_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5966 a_5349_15823 tdc0.r_ring_ctr13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X5967 tdc0.w_ring_buf17 a_4811_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5968 a_29435_20149 net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5969 _074_ a_26754_19133 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X5971 a_19651_12015 a_18869_12021 a_19567_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5972 tdc1.w_ring_norsz22 tdc1.w_ring_norsz6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5973 a_11873_17999 a_10883_17999 a_11747_18365 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5974 a_27489_13469 _052_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X5975 a_22653_20175 _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.102 ps=0.965 w=0.65 l=0.15
X5976 a_8857_10633 _147_ a_8775_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5979 a_23003_12559 _177_ a_22907_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X5980 a_9585_14191 net23 tdc0.w_ring_norsz26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R81 tdc1.g_ring321.stg01_68.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5981 a_2413_12335 _156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5982 a_24462_14847 a_24294_15101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X5986 VGND a_25203_10357 a_25137_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X5987 a_22638_14013 a_22365_13647 a_22553_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X5988 a_17490_20719 a_17243_21097 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X5989 a_23109_12559 _172_ a_23003_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X5990 _066_ a_24822_19133 a_25085_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5991 a_26735_15101 a_25953_14735 a_26651_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X5992 a_20153_11471 a_19163_11471 a_20027_11837 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X5994 a_23289_10927 tdc1.r_ring_ctr10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X5995 a_12447_14191 _080_ a_12529_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5996 a_17903_16599 tdc1.r_dly_store_ring28 a_18049_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X5997 VGND _103_ a_15027_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5998 VGND tdc1.w_ring_norsz3 a_20911_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X5999 VPWR a_8086_17429 a_8013_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6001 tdc1.r_ring_ctr13 a_18027_11445 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6002 a_11103_16189 a_10405_15823 a_10846_15935 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6003 tdc0.r_dly_store_ring28 a_9431_17179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6004 a_12901_18863 tdc0.r_dly_store_ring12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6006 VPWR a_8178_14165 a_8105_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6007 a_20911_15823 _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X6008 VPWR tdc1.r_ring_ctr4 a_24835_13335 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6009 a_1647_14569 a_1131_14197 a_1552_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6010 a_7507_16189 a_6725_15823 a_7423_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6011 VPWR a_23542_17429 a_23469_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6012 VGND _079_ a_14081_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6013 VGND a_13735_21263 _076_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6014 VGND a_12207_14013 a_12375_13915 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6015 a_6246_13759 a_6078_14013 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6016 VGND a_15904_11445 _624_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6017 a_23193_20725 a_23027_20725 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6018 a_11141_15285 a_10975_15285 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6019 VPWR tdc1.r_ring_ctr12 a_16861_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6021 VGND net35 a_22199_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6023 VGND net5 a_25971_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X6024 net8 a_9503_12015 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X6025 VPWR a_30959_15253 a_30875_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6026 VPWR _087_ a_20911_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X6027 VPWR net7 a_1315_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6028 net26 a_9647_15253 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
R82 net72 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6031 tdc1.w_ring_buf13 a_29375_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6033 VPWR net36 a_24131_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6035 VPWR a_2623_12335 _015_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X6037 a_14081_12393 a_13091_12021 a_13955_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6039 VGND tdc0.w_ring_norsz12 a_7479_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6041 a_19216_10383 _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6042 a_22469_16073 _080_ a_22671_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6043 a_13698_11989 a_13530_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6045 a_7079_11231 _039_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6046 a_9769_20425 net52 tdc0.w_ring_int_norsz23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6047 tdc0.w_ring_norsz16 tdc0.w_ring_int_norsz16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6049 a_2212_13481 a_1131_13109 a_1865_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6050 VPWR net27 a_3247_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6051 a_18785_14985 _133_ a_18703_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6052 tdc0.w_ring_int_norsz28 tdc0.w_ring_norsz27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6053 tdc0.w_ring_buf12 a_7479_17999 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6054 a_16861_9839 a_16831_9813 _019_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X6055 VPWR a_2743_12711 _158_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X6056 VGND a_19751_15279 a_19919_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6057 a_20993_20719 net66 tdc1.w_ring_int_norsz19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6058 a_19329_11471 a_19163_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6059 VPWR a_9431_17179 a_9347_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6060 VPWR a_13879_10901 tdc0.r_ring_ctr2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X6061 VGND tdc1.r_ring_ctr3 _171_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6062 a_12993_15279 _071_ a_13195_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R83 tdc0.g_ring321.stg01_50.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6064 a_13530_12015 a_13257_12021 a_13445_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6065 VGND a_14428_17687 _117_ VGND sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X6066 VPWR a_19395_17076 tdc1.w_ring_buf5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6067 a_19261_19337 tdc1.w_ring_norsz7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6068 a_20230_10383 _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6069 a_29791_18775 a_29887_18775 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6070 VPWR net28 a_8767_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6071 VGND tdc1.w_ring_norsz27 tdc1.w_ring_norsz11 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6073 VGND a_11490_14847 a_11448_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6074 VGND _069_ a_21993_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6075 tdc0.w_ring_int_norsz11 net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6076 a_16565_14735 a_15575_14735 a_16439_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6077 a_20258_16073 tdc1.r_dly_store_ctr13 a_20175_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6078 VPWR a_12507_10143 a_12494_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6080 net43 a_28047_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6083 VGND a_12559_21531 a_12517_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6084 a_14357_11293 a_13879_10901 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X6085 a_22603_17277 a_21905_16911 a_22346_17023 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6086 a_3571_19252 tdc0.w_dly_stop2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6087 a_17314_20996 a_17107_20937 a_17490_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6088 VGND net3 a_13735_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6090 a_14917_19631 tdc1.w_ring_buf2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6091 a_22005_11247 _179_ _184_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6094 _015_ _157_ a_2953_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X6095 a_30534_12559 _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6096 a_16656_16885 _089_ a_17044_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6097 a_21327_10071 tdc1.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6098 VGND _055_ a_25093_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6099 a_3513_12559 tdc0.r_ring_ctr8 a_3431_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X6100 a_17243_21097 a_17107_20937 a_16823_20951 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6102 VPWR a_5935_19355 a_5851_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6103 a_5875_11623 a_6018_11517 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X6104 a_15094_14013 a_14821_13647 a_15009_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6105 tdc0.w_ring_int_norsz30 net59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6106 a_24939_14013 _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6107 a_22281_14191 _080_ a_22135_14423 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X6108 VGND a_14623_16627 _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X6109 tdc0.r_ring_ctr11 a_4687_13407 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6111 a_13732_21039 _132_ a_13344_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X6112 VPWR _068_ a_24213_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6114 a_6339_11305 a_5823_10933 a_6244_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6115 VGND _067_ a_26785_17687 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X6116 VGND net9 a_18795_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6117 a_11831_15101 a_11049_14735 a_11747_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6118 a_22645_19087 tdc1.w_ring_buf10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6119 a_22937_20175 _075_ a_22527_20327 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X6120 VGND _122_ a_26581_18145 VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X6122 VGND _124_ a_20316_18151 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6123 VGND tdc0.w_ring_norsz23 tdc0.w_ring_norsz7 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6124 a_17945_17833 a_16955_17461 a_17819_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6126 a_28537_13647 tdc1.r_ring_ctr1 a_28455_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X6127 a_30258_17429 a_30090_17455 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6128 tdc1.w_ring_norsz13 net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
R84 net77 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6131 a_1647_13481 a_1131_13109 a_1552_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6132 VGND a_6687_14191 a_6855_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6133 net25 a_25839_16341 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6135 VGND _069_ a_12425_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6136 VGND a_20027_11837 a_20195_11739 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6137 net11 a_11435_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6139 VGND a_12007_15253 a_11965_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6142 a_17192_11471 _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6143 _174_ tdc1.r_ring_ctr4 a_24030_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X6144 net39 a_9839_17715 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X6145 VGND _110_ a_17924_17063 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6146 a_11937_11293 a_11893_10901 a_11771_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6147 VPWR a_6987_12247 _154_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X6148 VPWR a_30959_14165 a_30875_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6149 _058_ net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6150 VGND net7 a_1223_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6151 VGND _105_ a_22293_15395 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6152 VGND tdc1.w_ring_norsz29 a_30295_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6153 VPWR a_17159_18517 a_17075_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6154 tdc1.r_ring_ctr8 a_25203_10357 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X6157 a_21971_13335 a_22067_13335 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6158 VPWR a_11747_18365 a_11915_18267 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6160 a_11080_12559 a_10681_12559 a_10954_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6161 a_28737_12809 _170_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6164 VPWR a_23264_21237 net34 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6165 a_17593_10383 a_16403_10383 a_17484_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6167 VGND a_6487_15003 a_6445_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6171 a_27135_19849 net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6172 a_5602_15935 a_5434_16189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6173 tdc1.w_ring_int_norsz11 tdc1.w_ring_norsz10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6175 a_25009_13441 tdc1.r_ring_ctr5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X6176 a_17520_17833 a_17121_17461 a_17394_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6177 a_1736_15823 _005_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6179 a_11893_10901 a_11675_11305 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6181 net5 a_26667_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6183 VGND _079_ a_13989_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X6184 VGND _072_ a_13669_19115 VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X6185 a_13633_14985 _190_ a_13551_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6186 VPWR a_16825_15797 _077_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6188 a_25287_18517 a_25643_18775 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6189 a_18298_19605 a_18130_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6190 tdc0.w_ring_int_norsz8 net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6191 a_22143_19631 a_21445_19637 a_21886_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6194 a_19402_16341 a_19234_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6195 VGND tdc1.w_ring_int_norsz1 tdc1.w_ring_norsz1 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6196 a_14005_15823 tdc0.r_dly_store_ring3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6198 VGND net9 a_16771_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6201 VPWR net26 a_3339_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6202 VPWR tdc1.w_ring_norsz21 a_18509_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
R85 uio_out[4] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6204 a_16367_12559 a_15851_12559 a_16272_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6205 VGND a_23211_14735 net33 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6206 VGND a_16439_15101 a_16607_15003 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6207 VGND net7 a_3339_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6210 a_19234_16367 a_18961_16373 a_19149_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6211 a_21844_18921 a_21445_18549 a_21718_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6214 VPWR a_16219_11471 _625_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6216 a_24950_14468 a_24750_14313 a_25099_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6218 VPWR a_28915_10927 _198_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6219 VPWR _197_ _038_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6222 a_9765_14735 tdc0.w_ring_buf10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6223 VPWR net35 a_22751_19637 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6224 VGND net6 a_25971_18551 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6228 VGND net26 a_6559_13109 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6229 a_17489_19631 tdc1.w_ring_norsz7 a_17405_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6231 VGND net31 a_9963_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6233 a_28139_15511 a_28430_15401 a_28381_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6234 a_17857_19637 a_17691_19637 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6235 a_22711_12533 _172_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X6236 a_13989_14735 tdc0.r_dly_store_ctr0 a_13551_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6237 VPWR tdc0.r_ring_ctr8 a_2785_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6238 VGND a_29791_20938 tdc1.w_ring_buf15 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6239 VGND _197_ _032_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6240 uo_out[3] a_15196_16073 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6242 VGND a_26031_16885 net41 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6244 VGND a_10570_20287 a_10528_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6245 VGND tdc1.w_dly_stop1 a_15575_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6246 _059_ net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6248 tdc0.r_ring_ctr7 a_7079_11231 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6249 VGND _191_ a_17638_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6250 a_12537_21039 _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.189 ps=1.88 w=0.65 l=0.15
X6251 a_27491_15823 a_27271_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6252 a_29435_20149 net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6253 VGND _198_ _057_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6254 a_18141_11247 tdc1.r_ring_ctr12 _186_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6255 a_19659_16367 a_18961_16373 a_19402_16341 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6258 a_8596_13481 a_8197_13109 a_8470_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6259 VGND net32 a_16162_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X6260 a_13611_20327 _075_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6261 a_19234_16367 a_18795_16373 a_19149_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6263 a_30281_15279 tdc1.r_ring_ctr2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6264 net39 a_9839_17715 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X6265 VPWR tdc1.r_ring_ctr10 a_21185_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6266 VGND tdc1.w_ring_buf16 a_25849_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6267 VPWR a_12299_19453 a_12467_19355 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6271 a_13288_13481 a_12889_13109 a_13162_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6272 tdc0.w_ring_norsz11 tdc0.w_ring_norsz27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6273 VPWR tdc0.w_dly_stop1 a_2971_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6274 VGND a_17804_15279 uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6276 net38 a_29427_20693 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6277 a_13257_12021 a_13091_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6279 VGND a_24719_15101 a_24887_15003 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6280 a_14366_15599 tdc0.r_dly_store_ring18 a_14280_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X6282 VPWR a_17567_10099 net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6283 tdc0.w_ring_buf24 a_11159_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6284 _073_ a_12907_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6285 uo_out[1] a_17208_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6286 VPWR tdc0.r_ring_ctr10 a_5875_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X6287 tdc0.r_dly_store_ctr15 a_4279_17179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6290 VGND a_19395_17076 tdc1.w_ring_buf5 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6291 a_15715_17674 tdc1.w_ring_norsz4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6292 a_29055_20327 a_29151_20149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6293 a_10413_17161 net21 tdc0.w_ring_norsz3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6295 a_9389_16911 a_8399_16911 a_9263_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6296 a_27159_11989 a_27003_12257 a_27304_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X6297 a_6998_13103 a_6725_13109 a_6913_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6299 a_20169_11247 tdc1.r_ring_ctr11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6300 VPWR a_7867_12827 a_7783_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6301 a_4674_13103 a_3597_13109 a_4512_13481 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6302 VPWR tdc1.w_ring_norsz23 a_21923_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6303 VPWR _079_ a_12889_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6304 _169_ a_28823_14557 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X6305 VPWR a_28043_15511 tdc1.r_dly_store_ctr1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6306 a_20258_16073 _080_ a_20258_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X6307 a_29883_21428 ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6309 tdc1.r_ring_ctr3 a_30355_12533 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X6310 VGND a_30591_18267 a_30549_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6312 VPWR _147_ a_5791_12533 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0746 ps=0.775 w=0.42 l=0.15
X6313 _054_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6314 VPWR tdc0.r_ring_ctr12 a_3703_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X6315 a_22741_16367 tdc1.r_dly_store_ring3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X6316 a_25839_16341 _066_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6317 a_26597_20719 tdc1.w_ring_norsz16 a_26513_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6318 a_18639_19631 a_17857_19637 a_18555_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6320 VPWR net7 a_3339_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6321 VGND a_4443_18543 net20 VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6322 a_10827_20541 a_9963_20175 a_10570_20287 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6324 a_12723_18543 net24 a_12901_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X6325 a_7201_10625 a_6983_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6326 a_22707_13469 a_22487_13481 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6327 a_27090_12015 a_26964_12131 a_26686_12147 VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X6328 tdc1.r_dly_store_ctr5 a_26819_15003 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6329 VGND net19 tdc0.w_ring_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6330 tdc1.w_ring_buf16 a_25787_20719 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6332 a_18509_20719 net41 tdc1.w_ring_int_norsz7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6333 VPWR a_14032_16911 uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6334 VPWR a_27003_11169 a_26964_11043 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6335 _119_ a_12723_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6336 a_1949_15645 tdc0.r_ring_ctr13 a_1843_15645 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X6337 a_27607_11837 _048_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6338 VPWR a_19567_12015 a_19735_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6339 a_10497_20541 a_9963_20175 a_10402_20541 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6340 a_12415_11231 _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6341 a_1317_12559 _158_ _001_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.25 ps=1.42 w=0.65 l=0.15
X6342 VGND a_19567_12015 a_19735_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6344 a_28227_16911 a_28007_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6345 a_23358_19605 a_23190_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6346 a_7918_17455 a_7479_17461 a_7833_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6347 VGND net63 tdc1.w_ring_int_norsz16 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6348 VPWR a_19529_10625 a_19419_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6349 a_20625_20719 net15 tdc1.w_ring_norsz2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6350 VPWR tdc1.w_ring_int_norsz24 a_19973_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6351 a_29989_20175 a_29435_20149 a_29642_20149 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X6352 a_8987_15279 a_8123_15285 a_8730_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6353 a_29571_20175 a_29442_20449 a_29151_20149 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6354 VGND a_16656_16885 uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X6355 VPWR a_16932_12559 a_17107_12533 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6356 VGND tdc0.w_ring_norsz20 tdc0.w_ring_norsz4 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6358 tdc1.w_ring_norsz10 net15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6359 VPWR tdc1.w_ring_norsz28 a_29743_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6360 _011_ _150_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6361 a_23190_19631 a_22917_19637 a_23105_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6362 a_21768_14191 _075_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X6363 _068_ a_25287_18517 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6364 VPWR tdc1.w_ring_norsz9 a_20727_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6365 VGND net9 a_21739_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6367 a_8657_15279 a_8123_15285 a_8562_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6369 a_18014_11837 a_16937_11471 a_17852_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6370 VGND a_21463_15823 _089_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6371 VGND a_23323_19355 a_23281_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6372 _178_ a_22199_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6374 VGND net33 a_23855_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6375 a_18961_16373 a_18795_16373 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6377 a_17946_13103 a_17507_13109 a_17861_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6378 a_9865_18543 tdc0.w_ring_norsz5 a_9781_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6379 VPWR tdc1.w_ring_buf11 a_28425_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6380 tdc1.w_ring_int_norsz8 net41 a_19261_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6382 a_30281_14191 tdc1.r_ring_ctr3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6383 a_30641_17833 a_29651_17461 a_30515_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6384 a_13621_19951 tdc0.r_dly_store_ring31 a_13183_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6385 a_14852_19087 a_14453_19087 a_14726_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6387 a_12529_14191 tdc0.r_dly_store_ctr8 a_12447_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6388 net39 a_9839_17715 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6389 tdc1.w_ring_int_norsz31 net78 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6390 a_11675_11305 a_11159_10933 a_11580_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6391 a_22603_21629 a_21739_21263 a_22346_21375 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6392 a_20433_16911 a_20267_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6393 VPWR _008_ a_15118_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X6395 a_29913_17999 tdc1.w_ring_buf13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6398 VPWR a_29435_20149 a_29442_20449 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6400 VGND tdc1.w_ring_int_norsz15 tdc1.w_ring_norsz15 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6401 a_19567_12015 a_18703_12021 a_19310_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6402 _162_ a_5791_12533 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X6404 VPWR tdc0.w_ring_norsz21 a_9033_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6405 a_24131_16483 _096_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X6406 a_22143_12015 a_21445_12021 a_21886_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6407 VGND _037_ a_9453_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6408 VGND tdc1.r_ring_ctr1 a_28279_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6409 VGND a_28538_20996 a_28467_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X6410 VPWR a_17903_16599 _111_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X6412 a_27689_15823 a_27142_16097 a_27342_15797 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6413 a_22273_21629 a_21739_21263 a_22178_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6415 VGND _102_ a_15027_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6417 a_19237_12015 a_18703_12021 a_19142_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6418 a_21886_11989 a_21718_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6419 _025_ _170_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6421 a_14461_14985 _101_ a_14379_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6422 a_22343_15975 _081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X6423 a_8757_19337 net40 tdc0.w_ring_int_norsz7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6424 a_19751_15279 a_19053_15285 a_19494_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6425 a_18847_21237 a_19138_21537 a_19089_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6426 a_28266_21085 a_27951_20951 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X6427 a_22028_11471 a_21629_11471 a_21902_11837 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6428 VPWR net3 _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6429 a_18021_15797 _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X6430 a_4237_16911 a_3247_16911 a_4111_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6431 tdc0.r_dly_store_ctr1 a_15595_11989 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6432 a_21586_14191 _195_ a_21337_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X6434 a_14415_18365 a_13551_17999 a_14158_18111 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6436 _069_ a_14623_16627 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X6437 a_17484_10383 a_16569_10383 a_17137_10625 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6438 a_16097_16911 a_15550_17185 a_15750_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X6439 VPWR a_17505_11713 a_17395_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6440 tdc0.r_dly_store_ring26 a_11915_15003 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6442 tdc0.w_ring_buf28 a_7571_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6443 VPWR net34 a_23027_20725 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6444 VPWR net29 a_10975_15285 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6445 VPWR _079_ a_18869_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6446 uo_out[3] a_15196_16073 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6447 a_14085_18365 a_13551_17999 a_13990_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6448 VPWR _197_ _040_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6449 a_21445_20719 tdc1.w_ring_norsz2 a_21361_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6450 a_8197_13109 a_8031_13109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6451 VPWR tdc1.w_ring_norsz13 a_29089_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6452 a_6904_11305 a_5823_10933 a_6557_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6453 a_22820_10383 a_21739_10383 a_22473_10625 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6454 a_4069_13647 _161_ a_3851_13621 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6458 a_14158_18111 a_13990_18365 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6459 tdc0.r_dly_store_ctr9 a_9063_13077 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6460 VGND tdc0.w_dly_stop1 a_2971_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6461 a_24213_19337 tdc1.r_dly_store_ring31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6462 VGND a_14899_10143 tdc0.r_ring_ctr1 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6463 a_29925_13889 a_29707_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6464 a_17513_19337 tdc1.w_ring_norsz22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6466 a_25571_12319 a_25396_12393 a_25750_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6467 a_24463_10383 a_24113_10383 a_24368_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6469 a_16734_18517 a_16566_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
R86 VGND net73 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6470 tdc0.r_dly_store_ctr9 a_9063_13077 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6471 VPWR a_9891_12827 a_9807_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6472 a_26575_13077 a_26778_13235 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X6474 a_14817_14735 tdc0.r_dly_store_ctr3 a_14379_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6475 VPWR _090_ a_17596_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X6476 tdc0.r_dly_store_ctr2 a_13755_13077 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6477 a_26226_15101 a_25953_14735 a_26141_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6478 _134_ a_18703_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
R87 tdc1.g_ring324.stg01_71.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6479 VPWR tdc0.w_ring_norsz20 a_10331_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R88 VPWR tdc0.g_ring330.stg01_59.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6481 VPWR a_26483_10901 tdc1.r_ring_ctr9 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X6482 VPWR a_10492_10383 a_10667_10357 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6483 VPWR tdc1.r_ring_ctr0 a_28731_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X6485 a_20706_17277 a_20267_16911 a_20621_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
R89 uio_oe[4] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6486 a_16566_18543 a_16293_18549 a_16481_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6487 tdc1.w_ring_norsz24 tdc1.w_ring_norsz8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6489 VPWR a_28239_11445 a_28226_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6490 VPWR a_30180_12559 a_30355_12533 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6491 VPWR net33 a_23855_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6494 VPWR a_5602_15935 a_5529_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6495 a_23055_15975 tdc1.r_dly_store_ctr4 a_23201_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X6496 a_22346_21375 a_22178_21629 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6497 VGND a_25971_18551 _067_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X6499 a_9332_21097 a_8933_20725 a_9206_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
R90 net76 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6500 VPWR a_8143_18517 a_8059_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6501 a_16569_16373 a_16403_16373 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6502 VPWR a_22346_21375 a_22273_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6504 a_9332_15823 a_8933_15823 a_9206_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6505 VPWR _156_ a_2953_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6506 tdc0.r_dly_store_ctr10 a_6671_13915 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6508 tdc0.w_ring_int_norsz16 net39 a_4909_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6509 a_21065_15823 _086_ a_20993_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X6510 VPWR tdc0.r_ring_ctr0 _000_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6512 a_17596_20425 _090_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X6513 a_7549_20009 a_6559_19637 a_7423_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6515 a_9976_14735 a_9577_14735 a_9850_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6516 VGND a_29519_14165 _170_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6517 VGND _197_ _041_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6518 a_6273_13469 tdc0.r_ring_ctr9 a_6167_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X6519 VGND a_25381_17429 _086_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.176 ps=1.84 w=0.65 l=0.15
X6520 a_16823_20951 a_17114_20841 a_17065_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X6521 VPWR a_4595_11231 a_4582_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6522 tdc1.r_dly_store_ring25 a_23967_17429 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6524 _187_ a_17586_12335 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X6525 a_13637_18863 tdc0.r_dly_store_ring5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6527 tdc1.w_ring_int_norsz3 net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6528 a_11325_10933 a_11159_10933 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6529 tdc1.r_dly_store_ring25 a_23967_17429 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6531 tdc0.w_ring_buf19 a_10515_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6532 a_13445_12015 tdc0.r_ring_ctr3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6533 a_11747_15101 a_10883_14735 a_11490_14847 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6534 a_22806_13759 a_22638_14013 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6535 a_12475_21629 a_11693_21263 a_12391_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6537 VPWR a_14158_18111 a_14085_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6538 _148_ tdc0.r_ring_ctr3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6539 a_1739_16911 a_1223_16911 a_1644_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6541 VGND _131_ a_13732_21039 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6543 VPWR a_29057_21428 net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6544 VPWR _198_ _055_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6545 a_24227_16483 _097_ a_24131_16483 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6546 a_16566_18543 a_16127_18549 a_16481_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6547 a_22135_14423 tdc1.r_dly_store_ctr3 a_22281_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X6549 a_2743_12711 tdc0.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6550 VPWR tdc0.w_ring_norsz24 a_10229_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6551 tdc0.r_ring_ctr3 a_12415_11231 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6552 _183_ a_20819_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X6553 a_15679_16911 a_15550_17185 a_15259_16885 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X6554 a_2304_16911 a_1223_16911 a_1957_17153 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6555 a_24131_18249 _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
R91 net52 VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6556 a_21223_15101 a_20359_14735 a_20966_14847 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6557 VGND net77 tdc1.w_ring_int_norsz30 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6558 a_27346_17687 a_27815_17429 a_27759_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X6559 VPWR a_14899_10143 tdc0.r_ring_ctr1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6560 a_13809_9295 tdc0.r_ring_ctr1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6562 VPWR tdc1.w_ring_norsz17 a_22005_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6563 VGND net53 tdc0.w_ring_int_norsz24 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6564 a_17924_17063 _109_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X6565 VPWR tdc1.r_dly_store_ring5 a_20175_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X6566 a_14623_16627 _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X6567 VPWR tdc0.w_ring_norsz30 a_6457_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6570 a_7124_20009 a_6725_19637 a_6998_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6571 a_25505_13647 a_24315_13647 a_25396_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6572 a_22293_15395 _106_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6573 VGND a_22351_13321 a_22358_13225 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6574 VGND tdc1.w_ring_buf7 a_17661_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X6578 tdc0.w_ring_buf6 a_8675_20175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6579 a_25028_10383 a_23947_10383 a_24681_10625 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X6581 a_20966_14847 a_20798_15101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6582 a_19053_15285 a_18887_15285 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6583 _048_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6584 VGND tdc1.w_ring_norsz28 a_29743_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6585 tdc0.w_ring_norsz13 tdc0.w_ring_int_norsz13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6588 a_11322_15101 a_11049_14735 a_11237_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6589 VPWR a_15170_20693 a_15097_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6590 VPWR net16 _062_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6591 a_6177_14191 tdc0.r_ring_ctr11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6592 tdc0.r_dly_store_ring10 a_10443_15003 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6593 a_10667_10357 a_10492_10383 a_10846_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6595 tdc0.r_ring_ctr5 a_9931_11445 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X6596 _120_ a_13459_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X6598 a_18801_17455 tdc1.w_ring_norsz20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6599 a_18051_12015 tdc1.r_ring_ctr13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.153 ps=1.3 w=1 l=0.15
X6601 tdc0.w_ring_norsz4 net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6602 a_9121_20719 tdc0.w_ring_buf6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6603 VPWR a_22473_10625 a_22363_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6604 a_3855_14735 a_3339_14735 a_3760_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6606 a_26686_12147 a_27003_12257 a_26961_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X6607 VPWR tdc0.w_ring_norsz7 a_11057_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6608 a_26651_15101 a_25953_14735 a_26394_14847 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6609 VGND a_9839_17715 net39 VGND sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X6610 a_13669_19115 tdc0.r_dly_store_ring23 a_13583_19115 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6611 _174_ tdc1.r_ring_ctr5 a_23947_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6612 tdc1.w_ring_norsz26 net15 a_23021_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6613 VPWR a_21331_10901 _182_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X6614 tdc0.r_dly_store_ring9 a_15687_13915 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6615 a_20361_18543 tdc1.w_ring_int_norsz25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6618 VGND a_6607_11623 _152_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X6619 a_22346_17023 a_22178_17277 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6620 a_29642_15797 a_29435_15797 a_29818_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X6621 tdc1.w_ring_norsz1 tdc1.w_ring_norsz17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6622 VPWR a_2387_14495 a_2374_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6623 VPWR tdc0.w_ring_int_norsz15 a_5529_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6625 tdc0.r_dly_store_ring3 a_11271_16091 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6626 tdc0.w_ring_buf27 a_7295_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6627 tdc0.r_dly_store_ring22 a_10995_20443 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6628 a_10018_14847 a_9850_15101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6629 VPWR net27 a_8399_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6631 VPWR a_2304_16911 a_2479_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6633 VGND a_11547_12827 a_11505_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6634 tdc0.w_ring_buf8 a_15483_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6635 net33 a_23211_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6636 a_18751_21415 a_18847_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6639 VGND a_8435_14191 a_8603_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6640 a_29571_15823 a_29435_15797 a_29151_15797 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6641 a_3601_16911 tdc0.r_ring_ctr15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6643 _049_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6645 VPWR tdc1.w_ring_norsz14 a_28445_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6646 VGND a_3485_15253 _164_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X6648 a_2387_13407 a_2212_13481 a_2566_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6649 VGND _069_ a_13437_14511 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X6650 tdc0.w_ring_norsz18 net21 a_10509_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6651 _625_.X a_16219_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X6652 _198_ a_28915_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6653 a_21633_18543 tdc1.w_ring_buf21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6656 VGND a_6062_14847 a_6020_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6657 VGND a_16180_21237 net31 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6659 VPWR tdc1.r_ring_ctr10 a_21331_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X6660 VGND net73 tdc1.w_ring_int_norsz26 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6664 VPWR a_14799_11445 net29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6665 a_22711_12533 _183_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X6668 a_11533_10633 _147_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6669 a_19529_10625 a_19311_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6670 VPWR a_25028_10383 a_25203_10357 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6671 VPWR _197_ _037_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6672 VGND tdc0.w_ring_norsz20 a_10331_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6673 VGND a_18371_13103 a_18539_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6674 a_27814_13103 a_27056_13219 a_27251_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X6675 VGND a_23231_13915 a_23189_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6676 a_28047_21237 net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6678 VPWR net27 a_4903_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6680 VPWR a_15687_13915 a_15603_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6681 tdc0.w_ring_buf28 a_7571_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6682 a_29741_11989 a_29523_12393 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6684 VPWR _198_ _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6685 a_24508_16917 _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.127 ps=1.1 w=0.42 l=0.15
X6686 a_6607_11623 tdc0.r_ring_ctr6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6687 a_23381_20719 tdc1.w_ring_buf18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6688 VGND a_23967_10901 a_23925_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6689 _078_ a_15577_16483 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X6690 VPWR a_20027_11837 a_20195_11739 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6691 VPWR a_24275_16885 _071_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X6693 a_14366_15599 _076_ a_14197_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X6694 a_24462_14847 a_24294_15101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6695 VGND a_9631_20719 a_9799_20693 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6696 VPWR a_11271_16091 a_11187_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6697 VGND a_27491_17063 tdc1.r_dly_store_ring11 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6698 a_19521_18249 net41 tdc1.w_ring_int_norsz5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6699 VPWR a_17659_10357 a_17646_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6700 VGND tdc0.w_ring_norsz9 tdc0.w_ring_norsz25 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6701 a_19211_19850 tdc1.w_ring_norsz6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6702 a_25953_10927 tdc1.r_ring_ctr9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X6703 a_6403_15101 a_5621_14735 a_6319_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6705 VGND a_29435_20149 a_29442_20449 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6706 a_20874_17023 a_20706_17277 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6708 VPWR _057_ a_26483_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6709 a_4774_11293 _040_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X6710 a_1831_15823 a_1315_15823 a_1736_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6711 a_4585_17674 tdc0.w_ring_norsz0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6712 a_12935_12925 a_12153_12559 a_12851_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6713 a_1957_17153 a_1739_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6714 a_11509_19637 a_11343_19637 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6715 a_14833_10217 a_13643_9845 a_14724_10217 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6716 a_30917_16745 a_29927_16373 a_30791_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6717 a_12299_19453 a_11601_19087 a_12042_19199 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6718 a_11839_12015 a_10975_12021 a_11582_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6719 a_863_13897 _162_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6721 VPWR a_24995_16189 a_25163_16091 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6722 a_7097_20175 tdc0.w_ring_buf14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6723 a_22351_10383 a_21905_10383 a_22255_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6724 VGND net23 tdc0.w_ring_norsz11 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6726 a_8385_13103 tdc0.r_ring_ctr9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6727 a_29435_15797 net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6729 VGND a_21886_19605 a_21844_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6730 a_13077_13103 tdc0.r_ring_ctr2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6731 VGND a_13611_20327 _127_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X6732 VGND a_13559_9545 _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X6733 VPWR a_4111_17277 a_4279_17179 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6735 a_23101_10933 a_22935_10933 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6736 VPWR a_29055_20327 tdc1.r_dly_store_ring14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6737 VGND tdc1.w_ring_int_norsz3 tdc1.w_ring_norsz3 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6738 a_27159_10901 a_26964_11043 a_27469_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X6739 a_18371_13103 a_17507_13109 a_18114_13077 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6740 VGND a_4595_11231 tdc0.r_ring_ctr8 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6741 VGND _064_ a_24635_17973 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6742 a_7577_11721 tdc0.r_ring_ctr6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6743 a_18049_16687 _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X6745 VPWR net10 a_23947_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6746 VPWR net35 a_21279_18549 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6748 _197_ a_5087_11471 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6749 a_22748_16687 _087_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X6750 VPWR tdc1.w_ring_int_norsz4 a_19789_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6751 a_9927_10383 a_9577_10383 a_9832_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6753 a_18041_13103 a_17507_13109 a_17946_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6755 a_25513_16687 _068_ a_25103_16599 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X6757 a_22855_20425 tdc1.r_dly_store_ring9 a_22653_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6758 tdc1.r_ring_ctr12 a_17659_10357 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X6759 VGND net9 a_26983_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6760 VGND net16 _061_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6761 a_14081_14511 tdc0.r_dly_store_ctr2 a_13735_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6762 VPWR a_22143_18543 a_22311_18517 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6764 VGND a_9963_19631 net40 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6766 a_28630_15556 a_28430_15401 a_28779_15645 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6767 VGND a_17010_16341 a_16968_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6768 a_17505_11713 a_17287_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6769 VGND a_22143_18543 a_22311_18517 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6770 VPWR a_29833_12801 a_29723_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X6771 a_10570_20287 a_10402_20541 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6772 a_11414_12015 a_11141_12021 a_11329_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6773 VPWR tdc0.w_ring_int_norsz2 a_11141_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6775 VGND net8 a_9411_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6777 net11 a_11435_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6778 a_4073_14977 a_3855_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6779 a_29081_16367 tdc1.w_ring_norsz12 a_28997_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6780 a_15543_16885 net32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6781 VGND _088_ a_21463_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6782 VPWR a_22771_17179 a_22687_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6784 _063_ net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6787 _053_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6788 a_11417_9845 a_11251_9845 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6789 a_7815_11623 _149_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X6790 VPWR a_5087_11471 _197_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6791 a_11965_15657 a_10975_15285 a_11839_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6792 a_26667_21237 ui_in[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6793 a_26755_15975 a_26851_15797 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6794 VGND _183_ a_22005_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6796 _140_ a_24131_19337 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6797 a_15501_17277 a_15163_17063 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6798 VPWR a_19827_16341 a_19743_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6799 a_17107_12533 _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6800 tdc1.w_ring_norsz9 net15 a_20813_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6801 tdc1.w_ring_int_norsz23 net70 a_17513_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6803 a_30090_17455 a_29651_17461 a_30005_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6804 a_14642_20175 _143_ a_14172_20149 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6805 a_14159_10217 a_13809_9845 a_14064_10205 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6806 tdc0.w_ring_norsz27 net23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6807 a_25441_19631 net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X6808 VPWR tdc0.w_ring_norsz15 a_4903_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6810 a_6629_13647 a_5639_13647 a_6503_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6811 _089_ a_21463_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6812 tdc1.w_ring_int_norsz29 tdc1.w_ring_norsz28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6813 a_27555_17775 tdc1.r_dly_store_ctr5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.126 ps=1.11 w=0.42 l=0.15
X6815 a_22615_16599 _084_ a_23084_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6816 a_22553_13647 tdc1.r_ring_ctr15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6817 a_15163_17063 a_15259_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6818 a_27304_12015 a_27090_12015 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X6819 VGND net34 a_18795_16373 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6820 VGND a_8912_21237 net27 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6821 a_20599_12559 a_20249_12559 a_20504_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6822 a_22856_19087 a_22457_19087 a_22730_19453 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6823 _087_ net6 a_25441_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X6824 a_24481_12021 a_24315_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6825 a_27871_16885 net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6827 a_22143_18543 a_21279_18549 a_21886_18517 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X6832 a_3897_19337 net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6833 a_8013_17455 a_7479_17461 a_7918_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X6834 a_15719_21237 net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X6835 _015_ a_2623_12335 a_2861_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X6836 VPWR net35 a_20267_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6837 VPWR a_14172_20149 uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6838 a_29815_14013 _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6840 a_4989_17455 tdc0.w_ring_norsz17 a_4905_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6841 a_7718_18517 a_7550_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X6843 a_19268_12393 a_18869_12021 a_19142_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X6845 VGND _087_ a_21065_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6846 a_27829_17277 a_27491_17063 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X6847 _056_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6849 VPWR a_18114_13077 a_18041_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X6850 a_6633_10383 a_6467_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6852 VGND tdc1.w_ring_norsz18 a_21647_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6853 a_12993_15279 _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X6854 tdc0.r_ring_ctr0 a_12507_10143 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6855 a_15929_14735 net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6856 a_1927_15823 a_1481_15823 a_1831_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6857 a_12723_17161 _069_ a_12805_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X6858 a_30507_18365 a_29725_17999 a_30423_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X6859 a_5257_19087 tdc0.w_ring_buf15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6860 a_7550_18543 a_7277_18549 a_7465_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X6861 a_30527_18909 a_30307_18921 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X6863 a_25396_13647 a_24481_13647 a_25049_13889 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6864 a_7733_20175 a_6743_20175 a_7607_20541 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6865 VGND net34 a_16955_17461 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6866 a_6769_11471 _149_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X6867 a_27491_17063 a_27587_16885 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X6868 VGND tdc1.w_ring_norsz0 tdc1.w_ring_int_norsz1 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6869 VGND a_27679_21237 net42 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6870 VGND a_30263_12319 a_30197_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X6871 tdc0.w_ring_buf27 a_7295_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6872 VGND net31 a_13551_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6873 _188_ a_17691_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X6875 a_12425_15823 tdc0.r_dly_store_ring29 a_12079_16073 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6877 net6 a_25879_21263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6879 a_10869_12559 tdc0.r_ring_ctr4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X6880 a_1743_14569 a_1297_14197 a_1647_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6881 a_22160_20175 a_21934_20221 a_21791_20327 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6882 a_1909_13469 a_1865_13077 a_1743_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X6883 VPWR tdc1.w_ring_norsz24 a_18979_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6884 VPWR net30 a_16481_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X6885 tdc0.w_dly_stop4 a_3247_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6887 VGND a_11747_15101 a_11915_15003 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6888 a_23996_16599 _098_ a_24227_16483 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6889 VPWR net9 a_20083_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6890 a_19211_19850 tdc1.w_ring_norsz6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6891 VPWR a_4203_16189 a_4371_16091 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6893 a_24589_17821 tdc1.r_dly_store_ring25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.103 ps=1 w=0.42 l=0.15
X6895 VGND a_7591_13077 a_7549_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6896 VGND a_17562_17429 a_17520_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6897 tdc1.w_ring_buf24 a_18979_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6899 a_16175_20938 net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6901 VGND a_10995_20443 a_10953_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6902 VGND a_7718_18517 a_7676_18921 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X6903 a_14461_14985 _083_ a_14545_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6904 a_13541_18543 _076_ a_13459_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6905 a_7301_19337 tdc0.w_ring_norsz14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6906 tdc0.w_ring_buf21 a_8767_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X6910 VGND net34 a_21739_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6911 a_24463_10383 a_23947_10383 a_24368_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6912 tdc0.r_ring_ctr1 a_14899_10143 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X6913 a_29365_16367 net75 tdc1.w_ring_int_norsz28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6915 VPWR tdc0.r_ring_ctr9 a_3431_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X6916 _167_ tdc1.r_ring_ctr1 a_28814_13423 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X6918 _167_ tdc1.r_ring_ctr2 a_28731_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6919 a_14267_9839 a_13643_9845 a_14159_10217 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6920 a_3701_14511 _164_ a_3483_14423 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6921 a_7975_18543 a_7277_18549 a_7718_18517 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6923 a_27251_13077 a_27056_13219 a_27561_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X6924 VGND tdc0.w_ring_norsz20 tdc0.w_ring_int_norsz21 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6926 VPWR tdc0.w_ring_int_norsz8 a_10773_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6927 a_27095_13345 net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6930 a_10667_10357 _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6931 VGND net14 tdc1.w_ring_norsz24 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6933 a_14453_19087 a_14287_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6934 a_28226_11837 a_27149_11471 a_28064_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6935 VGND tdc1.r_ring_ctr4 a_26439_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6936 _114_ a_12723_17161 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X6937 a_22473_10625 a_22255_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X6938 tdc1.w_ring_int_norsz21 net68 a_18801_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6939 VGND tdc1.w_ring_norsz14 tdc1.w_ring_norsz30 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6940 VGND tdc0.w_ring_norsz4 a_12355_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6941 VPWR a_17208_20149 uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6942 a_11229_15823 a_10239_15823 a_11103_16189 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X6944 _067_ a_25971_18551 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6945 _009_ _147_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6946 tdc0.w_ring_int_norsz12 net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6947 VPWR tdc1.w_ring_int_norsz19 a_20617_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6948 VPWR tdc1.r_ring_ctr6 a_22905_13481 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X6949 a_28070_15101 a_27823_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X6950 VPWR a_23783_19605 a_23699_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X6951 net16 a_17567_10099 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R92 VGND net60 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6952 a_15059_13103 a_14361_13109 a_14802_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6953 VGND tdc1.w_ring_norsz23 a_21923_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X6954 VPWR _078_ a_17596_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6955 VPWR a_30171_18761 a_30178_18665 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6956 VGND net35 a_21279_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6957 a_29998_18365 a_29559_17999 a_29913_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X6959 a_21629_11471 a_21463_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6960 a_17596_20425 _091_ a_17208_20149 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6961 _170_ a_29519_14165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6962 a_24347_13441 _170_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X6963 a_30307_18921 a_30171_18761 a_29887_18775 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X6965 _041_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6967 VPWR a_23799_17455 a_23967_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6968 uo_out[6] a_13344_20693 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6969 a_21337_14165 _193_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X6970 VPWR a_28135_16586 tdc1.w_ring_buf11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X6973 a_6340_11721 _152_ a_5875_11623 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X6974 a_27090_12015 a_27003_12257 a_26686_12147 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X6975 VGND a_23799_17455 a_23967_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6977 a_6435_11305 a_5989_10933 a_6339_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6978 a_6059_11989 _155_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
R93 VGND net55 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X6979 VGND a_30959_16341 a_30917_16745 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6980 a_13551_14735 _083_ a_13729_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X6981 tdc1.w_ring_int_norsz12 net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6983 VPWR net32 a_14563_19637 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X6985 VGND tdc0.w_ring_int_norsz11 tdc0.w_ring_norsz11 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6986 a_11582_15253 a_11414_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X6988 a_3852_13469 _002_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X6989 tdc0.r_dly_store_ring11 a_9155_15253 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6991 a_1743_13481 a_1297_13109 a_1647_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6992 tdc0.w_ring_buf26 a_9227_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6993 VGND net35 a_20359_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6994 a_27346_17687 a_27705_17687 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X6995 VPWR _065_ a_24131_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X6996 tdc0.w_ring_norsz24 net22 a_11153_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6997 VPWR a_15427_19631 a_15595_19605 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X6998 VGND a_9799_16091 a_9757_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X6999 _190_ a_12447_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X7000 a_14917_20719 tdc0.w_ring_buf1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7001 VPWR a_24451_18864 a_24087_18775 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X7002 a_20825_20425 tdc1.w_ring_norsz1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7003 tdc1.w_ring_int_norsz30 tdc1.w_ring_norsz29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7004 a_1297_13109 a_1131_13109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7005 VPWR tdc1.r_dly_store_ctr12 a_18239_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X7006 VGND a_15427_19631 a_15595_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7007 VGND a_13344_20693 uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7008 a_20111_11837 a_19329_11471 a_20027_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7009 _095_ a_15117_14741 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X7010 a_12207_14013 a_11509_13647 a_11950_13759 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7014 VGND tdc1.w_ring_norsz9 a_20727_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7015 VPWR tdc0.w_ring_norsz9 a_14195_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7016 a_28241_14735 a_27687_14709 a_27894_14709 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7018 VPWR tdc0.w_ring_int_norsz5 a_9485_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7020 VGND a_20966_14847 a_20924_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7021 a_22729_16911 a_21739_16911 a_22603_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7023 VGND _198_ _054_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7024 VPWR tdc0.w_ring_norsz2 a_11067_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7025 VPWR tdc1.w_ring_norsz4 a_19521_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7027 a_30093_16373 a_29927_16373 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7030 a_23201_16073 _075_ a_23055_15975 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X7031 _071_ a_24275_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7033 a_11767_10217 a_11417_9845 a_11672_10205 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7035 VPWR a_25971_17999 _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7037 a_10035_10749 _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7038 VGND _054_ a_26721_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X7039 a_22905_13481 a_22351_13321 a_22558_13380 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7040 a_27894_14709 a_27687_14709 a_28070_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7042 a_25285_20203 net24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X7043 tdc0.r_dly_store_ctr6 a_9891_12827 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7044 VGND a_21791_20327 _090_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X7045 _135_ a_13583_19115 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X7046 a_21561_10205 tdc1.r_ring_ctr9 a_21489_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7048 VPWR a_6671_13915 a_6587_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7049 VGND tdc1.w_ring_norsz31 tdc1.w_ring_int_norsz0 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7050 VPWR a_28239_11445 tdc1.r_ring_ctr0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7051 VPWR tdc1.w_ring_int_norsz20 a_19421_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7052 a_21009_18249 tdc1.w_ring_norsz9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7053 VGND _067_ a_27351_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7055 a_11693_21263 a_11527_21263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
R94 tdc0.g_ring316.stg01_45.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7057 a_13265_19631 net24 a_13349_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7059 a_7189_12559 tdc0.r_ring_ctr7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7060 VPWR a_15519_14013 a_15687_13915 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7061 a_9577_14735 a_9411_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7062 VPWR _065_ a_27705_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.134 ps=1.48 w=0.42 l=0.15
X7063 _102_ a_14379_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X7064 a_27127_16885 tdc1.w_dly_stop5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X7065 a_5173_18543 tdc0.w_ring_norsz16 a_5089_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7066 VPWR tdc0.r_dly_store_ring9 a_17043_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X7067 VGND a_11582_17023 a_11540_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7068 a_11839_17277 a_10975_16911 a_11582_17023 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7069 tdc0.r_ring_ctr9 a_4687_12319 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7070 a_9715_16189 a_8933_15823 a_9631_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7071 tdc0.w_dly_stop4 a_3247_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7072 a_5529_19631 tdc0.w_ring_norsz31 a_5445_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7073 _153_ _150_ a_7577_11721 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7074 a_28047_20951 a_28338_20841 a_28289_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7075 VPWR _052_ a_27396_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X7076 a_25502_15556 a_25302_15401 a_25651_15645 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7077 VPWR tdc0.r_ring_ctr0 a_13809_9545 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7078 a_2479_16885 _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7079 a_22304_21263 a_21905_21263 a_22178_21629 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7080 VPWR a_18027_11445 a_18014_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7081 a_16463_12559 a_16017_12559 a_16367_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7082 VGND tdc1.r_dly_store_ring26 a_25513_16687 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X7084 a_29151_15797 a_29442_16097 a_29393_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X7085 a_24213_19087 tdc1.r_dly_store_ring23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7086 a_21327_10071 _179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7088 a_24939_12015 a_24315_12021 a_24831_12393 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7090 VPWR _065_ a_27517_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X7091 a_6447_10927 _039_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7092 tdc0.r_ring_ctr14 a_2571_15797 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X7093 a_28331_20937 net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7095 VGND net19 tdc0.w_ring_norsz14 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7096 tdc0.w_ring_buf21 a_8767_18543 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7097 a_14082_11059 a_14360_11043 a_14316_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X7098 a_10509_17455 tdc0.w_ring_norsz2 a_10425_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7099 a_13814_20719 _132_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X7101 _000_ tdc0.r_ring_ctr0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7102 VGND net8 a_13643_9845 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7103 VGND tdc1.w_ring_norsz11 tdc1.w_ring_norsz27 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7104 a_16727_20951 a_16823_20951 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7105 a_15451_20149 net24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X7107 tdc1.w_ring_norsz25 net15 a_20445_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7108 VPWR tdc1.w_ring_norsz15 a_27709_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7110 a_11141_15285 a_10975_15285 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7112 net29 a_14799_11445 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7113 a_12805_16073 _083_ a_12889_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7114 a_11747_18365 a_11049_17999 a_11490_18111 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7115 a_4621_18249 tdc0.w_ring_norsz0 a_4537_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7116 tdc0.r_ring_ctr4 a_10667_10357 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X7120 _037_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7121 VPWR net35 a_20359_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7122 VPWR _087_ a_21311_15617 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7124 tdc1.w_ring_int_norsz13 tdc1.w_ring_norsz12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7126 VGND _119_ a_14195_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.172 ps=1.83 w=0.65 l=0.15
X7127 VPWR _064_ a_26747_18863 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X7128 _052_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7129 a_22764_13647 a_22365_13647 a_22638_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7130 a_7833_17455 tdc0.w_ring_buf12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7131 VPWR _147_ a_6607_11623 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X7132 VGND a_21337_14165 _196_ VGND sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X7133 VPWR tdc0.w_ring_norsz16 a_5363_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7134 a_20993_15823 tdc1.r_dly_store_ring0 a_20911_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7137 a_20027_11837 a_19329_11471 a_19770_11583 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7138 a_11414_17277 a_11141_16911 a_11329_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7141 a_24455_17687 tdc1.r_dly_store_ring25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.141 ps=1.33 w=0.42 l=0.15
X7143 VPWR a_1865_13077 a_1755_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X7144 a_17646_10749 a_16569_10383 a_17484_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7145 tdc0.w_ring_norsz25 tdc0.w_ring_int_norsz25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7146 a_22269_20009 a_21279_19637 a_22143_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7147 VGND net14 tdc1.w_ring_norsz22 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7148 a_22363_10749 a_21739_10383 a_22255_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7149 a_6913_13103 tdc0.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7150 a_26839_17775 a_26785_17687 a_26739_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X7151 VPWR a_6430_14165 a_6357_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7152 a_6319_15101 a_5455_14735 a_6062_14847 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7153 a_29101_18249 tdc1.w_ring_int_norsz13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7155 a_8044_17833 a_7645_17461 a_7918_17455 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7156 a_22734_13103 a_22487_13481 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7157 tdc1.w_ring_norsz5 tdc1.w_ring_norsz21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7158 a_11875_9839 a_11251_9845 a_11767_10217 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7159 a_26483_10901 a_26686_11059 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X7161 a_20801_17277 a_20267_16911 a_20706_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7162 VPWR tdc1.w_ring_norsz14 a_29743_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7163 a_25505_12393 a_24315_12021 a_25396_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7164 VGND a_23211_12015 _179_ VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7167 a_3703_15279 tdc0.r_ring_ctr13 a_3485_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7168 a_16607_20502 tdc1.r_dly_store_ring1 a_16535_20502 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X7169 VPWR a_29435_15797 a_29442_16097 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7170 a_9647_15253 net28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X7172 tdc0.w_ring_int_norsz16 net45 a_3897_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7173 tdc0.w_ring_norsz9 tdc0.w_ring_norsz25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7175 a_9309_17455 net49 tdc0.w_ring_int_norsz20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7176 a_17302_14013 a_17029_13647 a_17217_13647 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7179 _088_ a_21311_15617 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X7181 a_16692_14569 a_16293_14197 a_16566_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7182 a_6062_14847 a_5894_15101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7184 VGND net41 tdc1.w_ring_int_norsz9 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7185 VGND a_30258_17429 a_30216_17833 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7187 a_26394_14847 a_26226_15101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7188 tdc1.w_ring_norsz3 tdc1.w_ring_norsz19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7190 VGND tdc1.w_ring_norsz16 tdc1.w_ring_int_norsz17 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7192 VGND a_18021_15797 _109_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7193 a_5989_10933 a_5823_10933 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7194 a_18072_13481 a_17673_13109 a_17946_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7195 a_9577_14735 a_9411_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7196 _624_.X a_15904_11445 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7197 a_5526_17277 a_5253_16911 a_5441_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7198 a_22005_20719 net65 tdc1.w_ring_int_norsz18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7199 a_15645_13647 a_14655_13647 a_15519_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7200 VPWR tdc0.w_ring_int_norsz26 a_9669_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7201 VPWR a_27135_15797 a_27142_16097 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7203 VGND tdc1.r_ring_ctr0 _016_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7204 VPWR net20 a_5087_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7205 a_19789_17455 tdc1.w_ring_norsz20 a_19705_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7206 VGND net9 a_20083_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7207 a_14158_18111 a_13990_18365 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7211 a_9865_11471 a_8675_11471 a_9756_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7212 a_1847_17277 _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7215 VPWR tdc1.w_ring_norsz27 a_26983_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7216 _061_ net16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7217 a_23937_15599 tdc1.r_dly_store_ctr15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7218 a_4130_16341 a_3962_16367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7220 VGND a_29057_21428 net4 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7221 a_12426_12925 a_12153_12559 a_12341_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7222 a_24485_15823 tdc1.w_ring_buf26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7223 a_27404_11471 _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X7224 a_20819_11471 tdc1.r_ring_ctr10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X7225 a_16439_15101 a_15741_14735 a_16182_14847 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7227 tdc0.w_ring_buf19 a_10515_15279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
R95 uio_oe[0] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7228 a_16014_15101 a_15575_14735 a_15929_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7229 a_9113_15657 a_8123_15285 a_8987_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7230 _039_ _197_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7231 VPWR a_17924_17063 _112_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X7232 VPWR a_15543_16885 a_15550_17185 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7234 VGND tdc0.w_ring_norsz2 a_11067_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7236 VGND tdc1.r_dly_store_ring29 a_27793_18909 VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X7238 VGND a_2656_18517 _626_.X VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X7239 VGND a_22070_11583 a_22028_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7240 VGND net33 a_19163_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7241 a_26426_17687 a_26895_17429 a_26839_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.15
X7242 VGND net22 tdc0.w_ring_norsz12 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7243 a_27093_19631 a_26755_19863 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X7244 VGND tdc0.w_ring_norsz5 tdc0.w_ring_int_norsz6 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7245 a_28425_16911 a_27878_17185 a_28078_16885 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7247 a_30492_15657 a_30093_15285 a_30366_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7248 VPWR a_26755_15975 tdc1.r_dly_store_ring27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7250 a_27823_14735 a_27694_15009 a_27403_14709 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7251 VGND a_14372_18543 uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0894 ps=0.925 w=0.65 l=0.15
X7252 tdc0.w_ring_int_norsz15 net39 a_7301_19337 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7253 a_29833_12801 a_29615_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X7254 VGND a_29791_18775 tdc1.r_dly_store_ring29 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7255 tdc1.w_ring_norsz11 tdc1.w_ring_int_norsz11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7256 VPWR a_29642_20149 a_29571_20175 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7258 a_22558_13380 a_22351_13321 a_22734_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7259 a_2571_15797 _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7260 a_15220_13647 a_14821_13647 a_15094_14013 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7261 VPWR tdc1.w_ring_norsz27 a_29365_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7262 VGND tdc1.w_ring_norsz30 tdc1.w_ring_norsz14 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7264 tdc0.w_ring_int_norsz4 net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7265 a_9213_12559 tdc0.r_ring_ctr6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7266 a_3851_13621 _161_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X7267 tdc0.w_ring_buf6 a_8675_20175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7268 VGND a_19770_11583 a_19728_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7269 a_14172_20149 _143_ a_14642_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7271 VPWR a_20874_17023 a_20801_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
R96 VPWR tt_um_hpretl_tt06_tdc_v2_92.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7275 VGND tdc0.w_ring_norsz11 tdc0.w_ring_norsz27 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7276 VPWR net5 a_25441_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7277 a_15151_19453 a_14287_19087 a_14894_19199 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7279 a_17819_17455 a_17121_17461 a_17562_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7280 a_18785_14985 _080_ a_18869_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7281 a_23201_15823 _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X7282 VPWR a_15163_17063 tdc1.r_dly_store_ring4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7283 a_11329_12015 tdc0.r_ring_ctr5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7284 tdc0.r_dly_store_ctr12 a_4555_16341 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7285 a_12867_15511 _129_ a_13195_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7287 VPWR net10 a_24315_12021 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7288 a_19437_13103 _188_ a_19355_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7289 a_7400_12559 a_7001_12559 a_7274_12925 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7291 a_2861_12335 _157_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7292 a_23855_15279 _071_ a_23937_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7294 a_13559_9545 tdc0.r_ring_ctr0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7295 a_11771_11305 a_11325_10933 a_11675_11305 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7296 a_7182_20541 a_6743_20175 a_7097_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7297 VGND a_16587_10927 tdc1.w_dly_stop5 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7298 VGND net7 a_3339_10933 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7299 VGND tdc1.r_ring_ctr13 a_17586_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X7300 VGND tdc0.w_ring_norsz7 a_11251_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7301 VPWR net29 a_10239_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7305 a_15553_21097 a_14563_20725 a_15427_20719 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7306 VPWR net7 a_6467_10383 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7307 a_23500_11305 a_23101_10933 a_23374_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7309 a_11490_14847 a_11322_15101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
R97 VGND net66 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7311 a_24546_20327 _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X7312 a_16656_16885 _100_ a_17044_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7313 a_17309_17455 tdc1.w_ring_buf22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7315 VPWR a_29099_19631 net37 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7316 VPWR _188_ a_19605_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7317 VGND a_24635_17973 _072_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7318 tdc0.w_ring_buf23 a_11067_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7319 a_22281_14511 _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X7321 VGND a_12134_21375 a_12092_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7322 net42 a_27679_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7324 a_23634_20693 a_23466_20719 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7325 a_20717_13647 tdc1.r_dly_store_ctr8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7326 a_12161_16073 tdc0.r_dly_store_ring29 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7327 a_6725_19637 a_6559_19637 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7328 a_6089_18543 net39 tdc0.w_ring_int_norsz14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7331 a_30381_13647 a_29191_13647 a_30272_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7332 a_28599_15797 net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X7333 a_21813_19631 a_21279_19637 a_21718_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7335 a_10681_12559 a_10515_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7336 VPWR a_9263_17277 a_9431_17179 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7337 VGND _160_ a_5261_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7339 a_20245_14569 a_19255_14197 a_20119_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7340 tdc0.r_dly_store_ring31 a_7591_19605 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7341 a_16481_18543 tdc0.w_ring_buf30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7343 a_26977_20719 tdc1.w_ring_norsz0 a_26893_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7344 a_16842_16367 a_16403_16373 a_16757_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7345 tdc1.w_ring_int_norsz2 net41 a_20825_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7346 tdc0.w_ring_int_norsz3 tdc0.w_ring_norsz2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7347 tdc0.r_dly_store_ring31 a_7591_19605 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7348 a_29523_12393 a_29007_12021 a_29428_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7349 VGND tdc1.w_ring_norsz14 a_29743_19631 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7350 VGND _067_ _074_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7351 _176_ tdc1.r_ring_ctr6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7353 a_8638_13077 a_8470_13103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7354 a_29725_17999 a_29559_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7355 VPWR net36 a_29927_14197 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7356 VPWR a_4512_12393 a_4687_12319 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7357 VPWR a_27251_13077 a_27182_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X7358 a_22269_12393 a_21279_12021 a_22143_12015 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7359 VGND a_20316_18151 _126_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X7360 VGND a_27159_10901 a_27090_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X7362 a_18939_20327 _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X7363 a_13330_13077 a_13162_13103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7364 _189_ tdc1.r_ring_ctr14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.176 ps=1.84 w=0.65 l=0.15
X7365 a_12897_17775 tdc0.r_dly_store_ctr15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7366 a_22365_13647 a_22199_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7367 VGND _079_ a_14817_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X7368 tdc0.w_ring_int_norsz21 net50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7369 a_29055_20327 a_29151_20149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7370 a_22457_19087 a_22291_19087 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7371 VPWR tdc0.r_ring_ctr1 a_13603_11445 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X7372 VPWR net34 a_21739_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7373 a_25049_11989 a_24831_12393 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X7374 VGND _113_ a_13461_17571 VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7375 VGND a_13735_21263 _076_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7376 a_12207_19631 a_11509_19637 a_11950_19605 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7377 VGND net31 a_14287_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7378 a_19877_15657 a_18887_15285 a_19751_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7379 tdc1.w_ring_norsz30 tdc1.w_ring_int_norsz30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7380 a_24835_13335 tdc1.r_ring_ctr5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X7381 _136_ a_12815_17455 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7382 a_4585_17674 tdc0.w_ring_norsz0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7383 a_21327_10071 tdc1.r_ring_ctr8 a_21561_10205 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7384 a_3693_15823 tdc0.r_ring_ctr14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7385 a_13541_18543 _089_ a_13625_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7389 a_17314_20996 a_17114_20841 a_17463_21085 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7390 a_20617_19631 tdc1.w_ring_norsz3 a_20533_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7391 a_11783_10927 _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7393 a_5069_19087 a_4903_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
R98 VGND net78 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7394 VPWR tdc0.w_ring_norsz10 a_8849_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7396 VGND tdc0.w_ring_norsz13 tdc0.w_ring_norsz29 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7398 a_7507_19631 a_6725_19637 a_7423_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7399 VPWR a_4443_18543 net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7402 VGND a_6059_11989 _156_ VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X7403 a_17208_20149 _089_ a_17596_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7405 a_12889_13109 a_12723_13109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7407 a_13437_14511 tdc0.r_dly_store_ring27 a_13091_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7410 tdc1.w_ring_norsz7 net14 a_17133_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7411 VPWR a_21886_19605 a_21813_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7413 VPWR _156_ a_3431_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X7415 a_5342_19453 a_4903_19087 a_5257_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7417 VPWR a_25111_20327 _139_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X7418 VGND _061_ a_17549_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7419 a_17804_15279 _196_ a_17638_15599 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X7420 a_3812_16911 a_3413_16911 a_3686_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7422 VPWR a_6503_14013 a_6671_13915 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7423 a_1835_16911 a_1389_16911 a_1739_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
R99 tdc0.g_ring116.stg02_44.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7427 _057_ _198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7428 a_25396_12393 a_24481_12021 a_25049_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7430 a_27397_11293 _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X7431 VPWR a_9631_16189 a_9799_16091 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7432 a_17470_13759 a_17302_14013 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7434 a_26961_11293 a_26483_10901 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X7435 VGND tdc1.w_ring_buf14 a_29989_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7436 VGND a_17727_14013 a_17895_13915 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7437 a_9693_13897 tdc0.w_ring_norsz25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7438 tdc0.r_dly_store_ring18 a_12007_17179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7439 VGND a_18243_17999 net14 VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X7440 a_27689_20009 a_27135_19849 a_27342_19908 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7442 VGND net20 _044_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7443 a_27271_20009 a_27142_19753 a_26851_19863 VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X7445 a_3597_13109 a_3431_13109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7447 VGND a_25571_13621 a_25505_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X7448 a_16831_9813 _185_ a_17217_9839 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7449 a_19487_21263 a_19267_21263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.09 w=0.42 l=0.15
X7450 a_13634_10383 tdc0.r_ring_ctr0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X7451 tdc0.r_dly_store_ring27 a_8603_14165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7452 tdc0.r_dly_store_ctr0 a_13019_12827 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7453 a_17638_15599 _196_ a_17804_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7454 VGND tdc0.w_ring_norsz15 a_4903_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7455 a_18877_17161 _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X7456 a_22527_20327 _084_ a_22855_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7457 a_6070_12559 _160_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.175 ps=1.26 w=0.42 l=0.15
X7458 a_14032_16911 _089_ a_13861_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7460 VGND a_2387_14495 a_2321_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X7462 a_12989_16367 tdc0.r_dly_store_ctr9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X7463 a_4513_16745 a_3523_16373 a_4387_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7464 VPWR a_12467_19355 a_12383_19453 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7465 a_8979_13103 a_8197_13109 a_8895_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7466 _064_ a_25971_17999 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X7468 a_9756_11471 a_8841_11471 a_9409_11713 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7469 VGND _044_ a_1909_14557 VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7470 a_24589_16917 _065_ a_24508_16917 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X7471 a_9931_11445 a_9756_11471 a_10110_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7473 VPWR _181_ a_21353_10633 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7475 a_10846_15935 a_10678_16189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7478 a_15199_14985 _094_ a_15117_14741 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7480 tdc1.w_ring_int_norsz0 net79 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7481 VGND a_17804_15279 uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7482 a_15170_20693 a_15002_20719 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7483 a_6339_11305 a_5989_10933 a_6244_11293 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7484 tdc1.r_ring_ctr0 a_28239_11445 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X7485 a_25861_11247 tdc1.r_ring_ctr9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7486 a_3951_14735 a_3505_14735 a_3855_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7487 VGND net31 a_11527_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7488 a_25251_19951 a_25221_19605 _087_ VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7490 a_29151_20149 a_29435_20149 a_29370_20175 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X7491 VPWR a_3571_19252 tdc0.w_dly_stop3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7492 _046_ net20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7493 tdc0.w_ring_buf23 a_11067_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7494 a_13349_19631 tdc0.r_dly_store_ring15 a_13265_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7495 VPWR a_17159_14165 a_17075_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7496 uo_out[4] a_14032_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7497 a_27070_15823 a_26755_15975 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7498 tdc0.r_dly_store_ring17 a_6119_17179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7499 VGND net4 a_27259_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X7500 VPWR tdc0.w_ring_int_norsz3 a_10497_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7501 a_5089_18543 tdc0.w_ring_int_norsz0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7503 _151_ tdc0.r_ring_ctr4 a_8850_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X7504 a_20893_15101 a_20359_14735 a_20798_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7505 VPWR a_24059_20693 a_23975_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7506 _091_ a_16607_20502 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X7508 tdc1.w_dly_stop4 a_16311_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7509 VPWR a_12007_15253 a_11923_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7511 VGND net22 tdc0.w_ring_norsz28 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7512 VPWR a_21131_17277 a_21299_17179 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7514 VGND tdc1.w_dly_stop2 a_15759_10927 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7515 a_8427_17455 a_7645_17461 a_8343_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7516 a_22473_10625 a_22255_10383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7518 net6 a_25879_21263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7519 a_19862_14165 a_19694_14191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7520 a_18298_19605 a_18130_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7524 a_14316_10927 a_13879_10901 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7525 a_30515_17455 a_29817_17461 a_30258_17429 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7526 a_8519_14191 a_7737_14197 a_8435_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7527 tdc1.w_ring_norsz27 tdc1.w_ring_int_norsz27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7529 a_20089_17455 tdc1.w_ring_norsz19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7531 VPWR a_14032_16911 uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7532 a_27403_17973 _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X7533 VGND a_27871_16885 a_27878_17185 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7534 a_23883_17455 a_23101_17461 a_23799_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7535 VGND a_14583_18267 a_14541_17999 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7539 VGND a_27135_19849 a_27142_19753 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7540 VGND net29 a_10975_15285 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7541 VGND a_22558_13380 a_22487_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0989 ps=0.995 w=0.64 l=0.15
X7542 a_12889_16073 tdc0.r_dly_store_ring21 a_12805_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7543 a_18130_19631 a_17857_19637 a_18045_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7546 a_1099_12744 tdc0.r_ring_ctr10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7547 VGND a_4404_19061 net19 VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X7548 a_29998_18365 a_29725_17999 a_29913_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7550 tdc1.r_dly_store_ctr3 a_30959_14165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7551 a_21311_15617 _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7552 VPWR _198_ _056_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7553 VPWR tdc1.w_ring_int_norsz2 a_20709_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7554 a_22286_13469 a_21971_13335 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X7555 a_15163_17063 a_15259_16885 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7556 a_26777_14735 a_25787_14735 a_26651_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7559 VGND a_22771_21531 a_22729_21263 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7560 a_3597_12021 a_3431_12021 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7561 VGND net26 a_5455_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7562 a_6913_19631 tdc0.w_ring_buf31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7563 tdc0.w_ring_buf13 a_6927_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7564 a_30725_18921 a_30171_18761 a_30378_18820 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7565 VGND tdc1.r_ring_ctr0 a_28241_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X7566 a_20451_18249 _084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.148 ps=1.34 w=0.42 l=0.15
X7568 VPWR a_16187_19891 _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7569 a_2227_15279 tdc0.r_ring_ctr13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.153 ps=1.3 w=1 l=0.15
X7570 a_29173_17161 tdc1.w_ring_norsz28 a_29089_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7571 _179_ a_23211_12015 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X7572 VPWR a_24251_19863 _097_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7573 VGND tdc0.r_ring_ctr5 _151_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7574 VPWR _147_ a_5271_12128 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7575 _131_ a_12618_21039 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.265 ps=2.53 w=1 l=0.15
X7576 a_7079_10383 a_6633_10383 a_6983_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7577 VGND a_20287_14165 a_20245_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7578 a_2321_14569 a_1131_14197 a_2212_14569 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
R100 VPWR tdc1.g_ring325.stg01_72.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7580 VPWR a_15427_12015 a_15595_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7581 a_22093_16911 tdc1.w_ring_buf3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7582 a_25705_11247 _180_ a_25623_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X7585 VGND net20 _043_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7587 a_30272_13647 a_29357_13647 a_29925_13889 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7588 VGND a_15427_12015 a_15595_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7589 VPWR a_20966_14847 a_20893_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7590 VPWR _065_ a_25551_17545 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.118 ps=1.4 w=0.42 l=0.15
X7591 a_8853_19631 tdc0.w_ring_norsz6 a_8769_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7592 a_21633_19631 tdc1.w_ring_buf9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7593 tdc1.w_ring_buf1 a_18887_20719 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7594 VGND tdc1.w_ring_int_norsz22 tdc1.w_ring_norsz22 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7595 tdc0.r_dly_store_ctr6 a_9891_12827 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7597 VPWR tdc1.r_dly_store_ring28 a_18049_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X7598 a_27815_17429 _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.0588 ps=0.7 w=0.42 l=0.15
X7599 VGND tdc1.w_ring_norsz5 tdc1.w_ring_norsz21 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7600 a_27722_10927 a_27003_11169 a_27159_10901 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X7601 _094_ a_13735_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X7602 VGND tdc0.w_ring_norsz4 tdc0.w_ring_int_norsz5 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7603 tdc0.w_ring_buf7 a_11251_20719 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7604 a_14267_9839 _033_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7605 a_9669_14191 tdc0.w_ring_norsz10 a_9585_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7606 _157_ tdc0.r_ring_ctr8 a_2413_12335 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7607 a_4595_14709 _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7608 a_10681_12559 a_10515_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7609 VGND a_22311_11989 a_22269_12393 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7611 a_14887_17494 tdc1.r_dly_store_ring4 a_14428_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X7612 a_11601_19087 a_11435_19087 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7613 a_4165_11989 a_3947_12393 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7616 a_27404_11471 _016_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7617 a_9191_11471 a_8841_11471 a_9096_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7618 tdc1.w_ring_buf12 a_28271_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7619 a_1957_17153 a_1739_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7620 a_5425_12381 _149_ a_5353_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X7622 a_14428_17687 tdc1.r_dly_store_ring4 a_14570_17821 VGND sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7623 a_20504_12559 _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X7625 VPWR a_29467_15287 _627_.X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7626 VGND a_28135_16586 tdc1.w_ring_buf11 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7628 VGND a_19919_15253 a_19877_15657 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7629 a_16656_16885 _100_ a_17126_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7630 a_25221_19605 net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7631 VPWR a_24835_13335 _172_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X7632 VPWR _197_ _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7633 VGND a_18939_20327 _132_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X7634 tdc1.w_dly_stop5 a_16587_10927 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X7635 a_11874_19453 a_11435_19087 a_11789_19087 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7636 VGND net21 tdc0.w_ring_norsz6 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7637 VGND _152_ _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7638 a_11122_12671 a_10954_12925 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7639 a_1755_13103 a_1131_13109 a_1647_13481 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7640 a_29707_13647 a_29191_13647 a_29612_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7641 _626_.X a_2656_18517 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7642 a_22365_13647 a_22199_13647 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7644 VGND a_21391_15003 a_21349_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7645 tdc0.w_ring_int_norsz6 net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7646 a_30355_12533 _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7647 VGND a_9503_12015 net8 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7649 a_3431_12559 tdc0.r_ring_ctr8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X7650 net9 a_25932_12533 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7651 a_30171_18761 net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7652 VGND tdc0.r_dly_store_ring25 a_16589_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X7653 a_7166_15935 a_6998_16189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7655 a_6167_13469 tdc0.r_ring_ctr10 a_6071_13469 VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X7656 VGND tdc0.w_ring_norsz9 a_14195_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7657 a_21164_12559 a_20083_12559 a_20817_12801 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7658 tdc1.w_ring_norsz8 net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7659 a_24297_15823 a_24131_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7660 a_9965_19337 tdc0.w_ring_int_norsz7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7661 a_23155_19453 a_22291_19087 a_22898_19199 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7662 VGND net34 a_17691_19637 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7663 VPWR a_24681_10625 a_24571_10749 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X7665 VGND _026_ a_27814_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X7666 a_22671_16073 tdc1.r_dly_store_ctr9 a_22469_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7667 a_11873_14735 a_10883_14735 a_11747_15101 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7668 tdc1.r_dly_store_ring0 a_19919_15253 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7670 a_19053_15285 a_18887_15285 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7671 VPWR net26 a_5455_14735 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7673 VPWR _064_ a_24631_16891 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7675 a_18869_14985 tdc1.r_dly_store_ctr14 a_18785_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7676 tdc1.r_dly_store_ring0 a_19919_15253 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7677 VGND net57 tdc0.w_ring_int_norsz28 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7679 a_14994_20175 _142_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X7680 a_25750_12381 _055_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7683 VPWR a_15715_17674 tdc1.w_ring_buf4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7684 VPWR _108_ a_15196_16073 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X7685 VPWR a_25049_13889 a_24939_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X7687 a_19602_11837 a_19329_11471 a_19517_11471 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7690 VGND net8 a_11159_10933 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7691 VGND a_10443_15003 a_10401_14735 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7692 VPWR a_17010_16341 a_16937_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7693 VGND _069_ a_20981_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
R101 VPWR tt_um_hpretl_tt06_tdc_v2_81.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7694 VGND a_14415_18365 a_14583_18267 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7695 VPWR a_15595_19605 a_15511_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7696 VPWR tdc0.r_ring_ctr1 a_13641_9545 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7699 a_26031_16885 net43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X7700 a_2321_13481 a_1131_13109 a_2212_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7701 a_8477_15279 tdc0.w_ring_buf11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7702 VPWR a_17484_10383 a_17659_10357 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7705 VGND net29 a_13091_12021 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7706 a_22070_11583 a_21902_11837 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7707 VPWR _069_ a_12529_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7708 a_11141_12021 a_10975_12021 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7709 VPWR a_29883_21428 net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7711 a_3963_15101 _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7712 a_29181_13103 _168_ _171_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7713 VGND tdc0.w_ring_int_norsz10 tdc0.w_ring_norsz10 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7714 net37 a_29099_19631 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X7715 VPWR a_22595_14887 _195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7716 VGND tdc0.w_ring_norsz29 tdc0.w_ring_int_norsz30 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7717 a_22135_14423 tdc1.r_dly_store_ctr11 a_22281_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7720 VPWR tdc0.w_ring_norsz18 a_10699_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7721 VGND tdc1.w_ring_buf0 a_26615_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X7722 a_17044_17161 _095_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7723 a_19770_11583 a_19602_11837 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7724 VPWR a_17895_13915 a_17811_14013 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7725 VPWR tdc0.r_ring_ctr12 a_1551_15253 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X7726 VGND net25 a_13161_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X7727 VPWR _067_ a_27346_17687 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X7728 a_20817_12801 a_20599_12559 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X7729 a_29519_14165 _169_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X7730 tdc0.r_dly_store_ring29 a_7591_16091 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7733 a_12851_12925 a_12153_12559 a_12594_12671 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7734 a_21993_16687 tdc1.r_dly_store_ring27 a_21647_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7736 tdc0.w_ring_buf18 a_10699_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7737 VPWR a_22527_20327 _085_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X7738 VPWR net29 a_10515_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7739 VGND a_7867_12827 a_7825_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7740 a_14486_10927 a_14360_11043 a_14082_11059 VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X7742 net16 a_17567_10099 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7743 a_24570_16189 a_24131_15823 a_24485_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7745 a_27469_11293 a_27090_10927 a_27397_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X7746 a_28806_15279 a_28559_15657 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7748 VGND a_21299_17179 a_21257_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7749 tdc0.r_ring_ctr6 a_7723_10357 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7750 a_30534_16341 a_30366_16367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7752 tdc0.w_ring_int_norsz26 net55 a_9693_13897 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7755 a_4073_14977 a_3855_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7757 VGND a_23259_18164 tdc1.w_ring_buf25 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7758 VGND a_30791_15279 a_30959_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7759 a_1389_16911 a_1223_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7760 a_11675_11305 a_11325_10933 a_11580_11293 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7762 VGND a_30263_12319 tdc1.r_ring_ctr1 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7763 a_4687_12319 _041_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7764 a_30366_16367 a_30093_16373 a_30281_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7765 VPWR a_26111_20938 tdc1.w_ring_buf16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7766 VGND a_25203_10357 tdc1.r_ring_ctr8 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7767 a_26833_18863 a_26431_18543 a_26747_18863 VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X7768 VGND tdc0.w_ring_norsz16 a_5363_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7769 a_9206_20719 a_8933_20725 a_9121_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7770 a_30281_14191 tdc1.r_ring_ctr3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7771 tdc0.r_dly_store_ring20 a_11915_18267 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7773 a_5951_17277 a_5253_16911 a_5694_17023 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7774 VGND a_29055_20327 tdc1.r_dly_store_ring14 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7775 a_27814_13103 a_27095_13345 a_27251_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X7776 VPWR a_22558_13380 a_22487_13481 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7777 VPWR tdc0.w_ring_norsz17 a_4811_16911 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
R102 tdc1.g_ring327.stg01_74.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7778 VPWR ui_in[5] a_25879_21263 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7779 a_9298_12925 a_8859_12559 a_9213_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7780 a_6077_16911 a_5087_16911 a_5951_17277 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7781 a_9931_11445 _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7782 VPWR tdc0.w_ring_int_norsz19 a_10129_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7783 tdc0.w_ring_norsz13 net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7784 a_13461_17571 _114_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7785 a_2656_18517 net19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X7786 VGND net11 tdc0.w_ring_int_norsz9 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7787 a_27689_20009 a_27142_19753 a_27342_19908 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0683 ps=0.745 w=0.42 l=0.15
X7788 VPWR net28 a_8123_15285 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7790 a_14729_20725 a_14563_20725 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7791 VGND net41 tdc1.w_ring_int_norsz11 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7792 a_8753_16911 tdc0.w_ring_buf28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7794 VPWR a_7591_16091 a_7507_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7795 _143_ a_14583_21590 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.158 ps=1.39 w=1 l=0.15
X7796 a_13344_20693 _131_ a_14166_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7797 a_24673_21513 net18 tdc1.w_ring_norsz17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7798 a_23358_19605 a_23190_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7800 VPWR a_27342_19908 a_27271_20009 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.08 w=0.75 l=0.15
X7801 a_6607_11623 _149_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X7802 a_11874_19453 a_11601_19087 a_11789_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7803 a_10846_10383 _036_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7804 VPWR tdc1.w_ring_norsz11 a_29641_16367 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7805 a_16824_10383 _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X7806 VPWR tdc1.r_ring_ctr12 a_18051_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.162 ps=1.33 w=1 l=0.15
X7807 a_16734_14165 a_16566_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7808 a_24736_13647 _027_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X7809 VPWR a_17562_17429 a_17489_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7811 a_17659_10357 a_17484_10383 a_17838_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X7812 VGND net40 tdc0.w_ring_int_norsz1 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7813 _156_ a_6059_11989 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7814 VGND _185_ a_16831_9813 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7815 net30 a_16162_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7816 VGND net35 a_21279_18549 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7817 a_21215_17277 a_20433_16911 a_21131_17277 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7818 a_16937_11471 a_16771_11471 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7820 VPWR tdc1.r_ring_ctr7 a_25016_11721 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X7821 a_16475_12925 _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7823 a_16566_14191 a_16293_14197 a_16481_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7824 a_3505_15823 a_3339_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7825 a_3505_14735 a_3339_14735 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7826 a_23634_20693 a_23466_20719 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7827 a_11582_15253 a_11414_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7828 a_30366_16367 a_29927_16373 a_30281_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7829 _035_ _197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7830 a_17181_10383 a_17137_10625 a_17015_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X7832 VGND tdc1.w_ring_norsz27 a_26983_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7833 a_18731_17063 tdc1.r_dly_store_ring22 a_18877_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7834 a_6244_11293 _013_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X7835 tdc1.w_ring_buf12 a_28271_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7836 a_28630_15556 a_28423_15497 a_28806_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X7837 a_23466_20719 a_23193_20725 a_23381_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7838 VGND a_22343_15975 _082_ VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X7840 tdc0.w_ring_int_norsz27 net56 a_7669_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7841 VGND a_14802_13077 a_14760_13481 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7842 VPWR net4 a_27259_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X7843 a_2049_16065 a_1831_15823 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X7845 tdc1.w_ring_norsz31 tdc1.w_ring_norsz15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7846 VGND a_21103_10633 _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7847 a_2566_13469 _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7849 a_28559_15657 a_28423_15497 a_28139_15511 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7850 a_27517_18543 _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X7851 VGND a_11839_17277 a_12007_17179 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7852 a_6062_14847 a_5894_15101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7853 a_2212_14569 a_1297_14197 a_1865_14165 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7854 VGND _118_ a_12723_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7855 VPWR a_17559_11159 _020_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X7856 a_14634_13103 a_14195_13109 a_14549_13103 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7857 a_26739_17775 _065_ a_26635_17775 VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X7858 _044_ net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7859 a_14857_17753 _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7861 VGND a_2703_10927 _014_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7862 a_12594_12671 a_12426_12925 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X7863 a_24765_20719 net18 tdc1.w_ring_norsz1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7866 VPWR a_13603_11445 _146_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X7867 VGND net26 a_8031_13109 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7868 a_4055_12015 _041_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X7869 _051_ _198_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7870 VGND a_11950_19605 a_11908_20009 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7871 VGND a_14857_17753 a_14791_17821 VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7872 a_12240_11305 a_11159_10933 a_11893_10901 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X7873 VGND a_17659_10357 tdc1.r_ring_ctr12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7875 VPWR a_26575_13077 tdc1.r_ring_ctr4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X7876 a_17638_15599 _192_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7877 VGND _173_ _027_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7878 VPWR tdc1.w_ring_norsz13 a_29375_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7879 VGND net47 tdc0.w_ring_int_norsz18 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7880 VPWR tdc0.w_ring_norsz30 a_6651_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7881 VPWR tdc0.r_dly_store_ring14 a_13611_20327 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7884 a_27679_21237 net43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X7885 a_19310_11989 a_19142_12015 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X7886 tdc1.r_ring_ctr15 a_21339_12533 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7887 a_21813_12015 a_21279_12021 a_21718_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7889 a_11839_15279 a_11141_15285 a_11582_15253 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7890 net40 a_9963_19631 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X7891 _028_ _175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7893 a_11414_15279 a_10975_15285 a_11329_15279 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7894 a_1865_13077 a_1647_13481 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X7896 VGND tdc1.r_ring_ctr9 a_25705_11247 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X7897 VPWR a_25571_12319 a_25558_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7898 a_3778_16189 a_3339_15823 a_3693_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7899 a_11141_17455 tdc0.w_ring_norsz18 a_11057_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7901 VPWR a_27717_11713 a_27607_11837 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X7902 a_10497_17161 tdc0.w_ring_norsz19 a_10413_17161 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7903 a_1481_15823 a_1315_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7904 a_25297_14569 a_24743_14409 a_24950_14468 VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X7905 VGND a_28043_15511 tdc1.r_dly_store_ctr1 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7906 a_23259_18164 tdc1.w_ring_norsz25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7907 a_18417_12809 _189_ _021_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7908 VPWR a_4687_13407 a_4674_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7909 VGND a_22711_12533 _185_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X7910 VPWR a_14857_17753 a_14887_17494 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7911 VPWR tdc1.w_ring_norsz2 a_20441_20425 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7912 VGND net8 a_11251_9845 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7915 VGND _154_ a_5425_12381 VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7916 a_18509_18543 net69 tdc1.w_ring_int_norsz22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7917 a_6078_14013 a_5639_13647 a_5993_13647 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7919 a_25103_16599 _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X7920 a_19514_21629 a_19267_21263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X7922 uo_out[0] a_17804_15279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X7923 a_3413_16911 a_3247_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7924 a_28415_21237 ui_in[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X7926 a_3505_14735 a_3339_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7927 a_14994_20175 _138_ a_14172_20149 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7928 a_15009_13647 tdc0.w_ring_buf9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7929 VPWR a_11103_16189 a_11271_16091 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7930 VPWR net33 a_18887_15285 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7932 a_11329_15279 tdc0.w_ring_buf19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7935 a_9298_12925 a_9025_12559 a_9213_12559 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X7936 uo_out[4] a_14032_16911 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7937 a_23799_17455 a_22935_17461 a_23542_17429 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X7938 tdc0.r_dly_store_ring16 a_6487_15003 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7939 _062_ net16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
R103 tdc1.g_ring320.stg01_67.HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
X7940 a_27003_11169 net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7943 VPWR a_12240_11305 a_12415_11231 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7944 VGND a_23363_12711 _177_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X7945 a_8933_15823 a_8767_15823 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7946 VGND tdc0.w_ring_norsz18 a_10699_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7947 a_22469_16073 _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.157 ps=1.32 w=1 l=0.15
X7948 a_3877_16367 tdc0.r_ring_ctr12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7950 _176_ _173_ a_25149_12809 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7953 net27 a_8912_21237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7954 a_14372_18543 _120_ a_14278_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X7955 a_23469_17455 a_22935_17461 a_23374_17455 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X7956 a_27342_15797 a_27142_16097 a_27491_15823 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X7958 a_27823_14735 a_27687_14709 a_27403_14709 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X7959 tdc0.w_ring_buf18 a_10699_16911 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7960 a_20709_20719 tdc1.w_ring_norsz18 a_20625_20719 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7962 a_19360_16745 a_18961_16373 a_19234_16367 VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7964 a_2212_13481 a_1297_13109 a_1865_13077 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7966 a_6177_14191 tdc0.r_ring_ctr11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X7967 a_23289_10927 tdc1.r_ring_ctr10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7968 tdc0.r_ring_ctr8 a_4595_11231 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X7969 a_10037_14191 tdc0.w_ring_norsz26 a_9953_14191 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7970 VPWR tdc1.r_ring_ctr13 _186_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7971 VGND _151_ _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7972 tdc0.w_ring_buf10 a_9135_14735 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X7973 VGND net18 tdc1.w_ring_norsz15 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7974 VPWR a_16187_19891 _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7975 a_21905_10383 a_21739_10383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7978 a_22227_19631 a_21445_19637 a_22143_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7979 _168_ a_28455_13647 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X7981 a_23537_12587 tdc1.r_ring_ctr7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X7982 VPWR a_27159_10901 a_27090_10927 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X7983 VPWR a_21886_11989 a_21813_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X7984 a_8561_14569 a_7571_14197 a_8435_14191 VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7986 a_29089_17161 net17 tdc1.w_ring_norsz12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7987 a_27722_12015 a_26964_12131 a_27159_11989 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X7988 _066_ _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X7989 tdc0.r_dly_store_ctr0 a_13019_12827 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7990 a_22753_15823 _080_ a_22343_15975 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X7992 VPWR _065_ a_26431_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X7993 tdc0.w_ring_norsz21 net21 a_9865_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7994 VPWR _076_ a_14329_21590 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.118 ps=1.4 w=0.42 l=0.15
X7995 a_5943_16189 a_5161_15823 a_5859_16189 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7996 VGND tdc0.w_ring_norsz17 a_4811_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X7997 VPWR a_15451_20149 _075_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7998 tdc1.r_ring_ctr2 a_30447_13621 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7999 VPWR a_27491_17063 tdc1.r_dly_store_ring11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8000 VPWR a_14623_16627 _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X8002 a_30166_18111 a_29998_18365 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X8003 VGND tdc1.w_ring_norsz30 tdc1.w_ring_int_norsz31 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8004 a_22687_21629 a_21905_21263 a_22603_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8006 VPWR tdc0.w_ring_int_norsz16 a_4241_18543 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8007 VPWR a_22603_17277 a_22771_17179 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8008 a_8769_19631 tdc0.w_ring_int_norsz22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8009 tdc1.w_ring_buf21 a_19071_18543 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8010 a_3778_16189 a_3505_15823 a_3693_15823 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8011 a_14082_11059 a_14399_11169 a_14357_11293 VGND sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X8012 VPWR a_16155_15975 _070_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X8014 VPWR a_11122_12671 a_11049_12925 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X8015 VGND a_30171_18761 a_30178_18665 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8019 tdc1.w_ring_norsz21 tdc1.w_ring_int_norsz21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8020 a_19338_21237 a_19131_21237 a_19514_21629 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0767 ps=0.785 w=0.42 l=0.15
X8022 a_20316_18151 _125_ a_20547_18249 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X8023 a_9191_11471 a_8675_11471 a_9096_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8024 VGND net29 a_10515_12559 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8025 a_20258_15823 tdc1.r_dly_store_ctr13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X8026 VGND _076_ a_14329_21590 VGND sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.109 ps=1.36 w=0.42 l=0.15
X8027 VPWR net31 a_11435_19087 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8028 VPWR tdc1.r_ring_ctr3 a_29181_13103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8029 a_15002_19631 a_14729_19637 a_14917_19631 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X8030 VGND a_9279_21237 net28 VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X8031 VGND a_15170_20693 a_15128_21097 VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8032 VGND _171_ _025_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8033 VGND a_9931_11445 a_9865_11471 VGND sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X8034 a_14545_14985 tdc0.r_dly_store_ring19 a_14461_14985 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8035 a_19267_21263 a_19131_21237 a_18847_21237 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X8036 a_28078_16885 a_27878_17185 a_28227_16911 VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X8037 VPWR net27 a_3523_16373 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8038 a_16017_12559 a_15851_12559 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8039 VPWR a_27951_20951 tdc1.r_dly_store_ring15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8040 a_17126_16911 _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X8041 a_14499_18365 a_13717_17999 a_14415_18365 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X8043 a_28361_12015 tdc1.r_ring_ctr0 a_28279_12015 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8044 a_5989_15101 a_5455_14735 a_5894_15101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X8045 tdc0.w_ring_buf24 a_11159_14191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X8046 VPWR tdc0.w_ring_norsz1 a_5455_17999 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X8047 a_30106_18909 a_29791_18775 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X8048 tdc1.w_ring_norsz29 tdc1.w_ring_norsz13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8049 a_17217_13647 tdc1.r_ring_ctr12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X8050 a_21337_14165 _195_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X8051 VGND tdc1.w_ring_norsz13 a_29375_18543 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X8052 a_24251_19863 tdc1.r_dly_store_ring18 a_24397_19951 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X8053 VPWR a_6687_14191 a_6855_14165 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8055 VGND net33 a_22935_10933 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8056 VPWR net25 a_23937_15279 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8057 a_13955_12015 a_13257_12021 a_13698_11989 VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X8058 a_16757_16367 tdc1.w_ring_buf20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X8059 VGND tdc1.w_ring_norsz24 tdc1.w_ring_norsz8 VGND sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8060 a_19985_10383 a_18795_10383 a_19876_10383 VGND sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X8063 _147_ a_11763_11445 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 ena VGND 0.0979f
C1 clk VGND 0.0979f
C2 rst_n VGND 0.0979f
C3 ui_in[6] VGND 0.0979f
C4 ui_in[7] VGND 0.0979f
C5 uio_in[0] VGND 0.0979f
C6 uio_in[1] VGND 0.0979f
C7 uio_in[2] VGND 0.0979f
C8 uio_in[3] VGND 0.0979f
C9 uio_in[4] VGND 0.0979f
C10 uio_in[5] VGND 0.0979f
C11 uio_in[6] VGND 0.0979f
C12 uio_in[7] VGND 0.0979f
C13 uo_out[0] VGND 3.65f
C14 uo_out[3] VGND 3.35f
C15 uo_out[2] VGND 2.88f
C16 uo_out[4] VGND 2.73f
C17 uo_out[5] VGND 1.98f
C18 uo_out[1] VGND 1.57f
C19 uo_out[7] VGND 2.13f
C20 uo_out[6] VGND 1.28f
C21 uio_out[0] VGND 1.23f
C22 ui_in[0] VGND 1.05f
C23 ui_in[1] VGND 1.17f
C24 ui_in[3] VGND 1.64f
C25 ui_in[2] VGND 1.05f
C26 ui_in[4] VGND 0.928f
C27 ui_in[5] VGND 0.87f
C28 uio_out[1] VGND 0.967f
C29 uio_out[2] VGND 0.967f
C30 uio_out[3] VGND 0.967f
C31 uio_out[4] VGND 0.989f
C32 uio_out[5] VGND 0.969f
C33 uio_out[6] VGND 0.967f
C34 uio_out[7] VGND 0.967f
C35 uio_oe[0] VGND 0.967f
C36 uio_oe[1] VGND 0.967f
C37 uio_oe[2] VGND 1.05f
C38 uio_oe[3] VGND 0.967f
C39 uio_oe[4] VGND 1.03f
C40 uio_oe[5] VGND 0.967f
C41 uio_oe[6] VGND 0.967f
C42 uio_oe[7] VGND 0.967f
C43 VPWR VGND 2.88p
C44 a_13809_9545 VGND 0.219f
C45 a_13559_9545 VGND 0.684f
C46 a_23653_9839 VGND 0.219f
C47 a_16861_9839 VGND 0.219f
C48 a_14267_9839 VGND 0.168f
C49 a_14064_10205 VGND 0.259f
C50 a_11875_9839 VGND 0.168f
C51 a_11672_10205 VGND 0.259f
C52 a_23403_9839 VGND 0.684f
C53 a_21327_10071 VGND 0.619f
C54 a_17567_10099 VGND 1.2f
C55 a_16831_9813 VGND 0.684f
C56 a_14724_10217 VGND 0.736f
C57 a_14899_10143 VGND 1.13f
C58 a_14159_10217 VGND 0.714f
C59 _033_ VGND 1.64f
C60 a_14377_9813 VGND 0.653f
C61 a_13809_9845 VGND 1.57f
C62 _007_ VGND 1.24f
C63 a_13643_9845 VGND 1.92f
C64 a_12332_10217 VGND 0.736f
C65 a_12507_10143 VGND 1.54f
C66 a_11767_10217 VGND 0.714f
C67 _032_ VGND 1.8f
C68 a_11985_9813 VGND 0.653f
C69 a_11417_9845 VGND 1.57f
C70 _000_ VGND 1.28f
C71 a_11251_9845 VGND 1.92f
C72 a_24571_10749 VGND 0.168f
C73 a_24368_10383 VGND 0.259f
C74 a_25028_10383 VGND 0.736f
C75 a_25203_10357 VGND 1.13f
C76 a_24463_10383 VGND 0.714f
C77 _056_ VGND 1.64f
C78 a_24681_10625 VGND 0.653f
C79 a_24113_10383 VGND 1.57f
C80 _030_ VGND 1.34f
C81 a_23947_10383 VGND 1.92f
C82 a_22363_10749 VGND 0.168f
C83 a_22160_10383 VGND 0.259f
C84 a_22820_10383 VGND 0.736f
C85 a_22995_10357 VGND 0.971f
C86 a_22255_10383 VGND 0.714f
C87 _058_ VGND 1.66f
C88 a_22473_10625 VGND 0.653f
C89 a_21905_10383 VGND 1.57f
C90 a_21739_10383 VGND 1.92f
C91 _017_ VGND 1.08f
C92 a_21353_10633 VGND 0.219f
C93 a_19419_10749 VGND 0.168f
C94 a_19216_10383 VGND 0.259f
C95 a_21103_10633 VGND 0.684f
C96 _181_ VGND 1.16f
C97 a_19876_10383 VGND 0.736f
C98 a_20051_10357 VGND 0.971f
C99 a_19311_10383 VGND 0.714f
C100 _059_ VGND 1.61f
C101 a_19529_10625 VGND 0.653f
C102 a_18961_10383 VGND 1.57f
C103 a_18795_10383 VGND 1.92f
C104 a_17027_10749 VGND 0.168f
C105 a_16824_10383 VGND 0.259f
C106 a_17484_10383 VGND 0.736f
C107 a_17659_10357 VGND 1.13f
C108 a_16919_10383 VGND 0.714f
C109 _060_ VGND 1.64f
C110 a_17137_10625 VGND 0.653f
C111 a_16569_10383 VGND 1.57f
C112 _019_ VGND 1.26f
C113 a_16403_10383 VGND 1.92f
C114 a_13551_10633 VGND 0.238f
C115 a_10035_10749 VGND 0.168f
C116 a_9832_10383 VGND 0.259f
C117 _144_ VGND 0.674f
C118 a_10492_10383 VGND 0.736f
C119 a_10667_10357 VGND 0.971f
C120 a_9927_10383 VGND 0.714f
C121 _036_ VGND 1.66f
C122 a_10145_10625 VGND 0.653f
C123 a_9577_10383 VGND 1.57f
C124 a_9411_10383 VGND 1.92f
C125 _010_ VGND 1.08f
C126 a_9025_10633 VGND 0.219f
C127 a_7091_10749 VGND 0.168f
C128 a_6888_10383 VGND 0.259f
C129 a_8775_10633 VGND 0.684f
C130 a_7548_10383 VGND 0.736f
C131 a_7723_10357 VGND 0.971f
C132 a_6983_10383 VGND 0.714f
C133 _038_ VGND 1.64f
C134 a_7201_10625 VGND 0.653f
C135 a_6633_10383 VGND 1.57f
C136 a_6467_10383 VGND 1.92f
C137 a_27304_10927 VGND 0.168f
C138 a_27722_10927 VGND 0.259f
C139 a_25861_11247 VGND 0.211f
C140 a_23289_10927 VGND 0.23f
C141 a_20169_11247 VGND 0.171f
C142 _018_ VGND 1.43f
C143 a_17777_11247 VGND 0.171f
C144 a_14700_10927 VGND 0.168f
C145 a_15118_10927 VGND 0.259f
C146 _148_ VGND 1.56f
C147 a_11783_10927 VGND 0.168f
C148 a_8767_10927 VGND 0.238f
C149 a_11580_11293 VGND 0.259f
C150 _012_ VGND 1.59f
C151 a_6447_10927 VGND 0.168f
C152 a_6244_11293 VGND 0.259f
C153 a_3963_10927 VGND 0.168f
C154 a_2953_10927 VGND 0.219f
C155 a_3760_11293 VGND 0.259f
C156 a_28915_10927 VGND 0.988f
C157 _031_ VGND 1.63f
C158 a_27090_10927 VGND 0.653f
C159 a_27159_10901 VGND 0.714f
C160 a_26964_11043 VGND 1.57f
C161 a_27003_11169 VGND 1.92f
C162 _057_ VGND 1.68f
C163 a_26686_11059 VGND 0.736f
C164 a_26483_10901 VGND 0.971f
C165 a_25623_11247 VGND 0.706f
C166 _180_ VGND 1.1f
C167 a_23799_10927 VGND 0.609f
C168 a_23967_10901 VGND 0.817f
C169 a_23374_10927 VGND 0.626f
C170 a_23542_10901 VGND 0.581f
C171 a_23101_10933 VGND 1.43f
C172 a_22935_10933 VGND 1.81f
C173 a_21331_10901 VGND 0.729f
C174 _182_ VGND 1.05f
C175 a_19951_11159 VGND 0.546f
C176 _184_ VGND 2.63f
C177 _186_ VGND 0.782f
C178 a_17559_11159 VGND 0.546f
C179 a_16587_10927 VGND 0.698f
C180 tdc1.w_dly_stop4 VGND 0.688f
C181 a_16311_10927 VGND 0.524f
C182 tdc1.w_dly_stop3 VGND 0.8f
C183 a_15759_10927 VGND 0.524f
C184 _008_ VGND 1.57f
C185 a_14486_10927 VGND 0.653f
C186 a_14555_10901 VGND 0.714f
C187 a_14360_11043 VGND 1.57f
C188 a_14399_11169 VGND 1.92f
C189 _034_ VGND 1.68f
C190 a_14082_11059 VGND 0.736f
C191 a_13879_10901 VGND 0.971f
C192 a_13323_11159 VGND 0.619f
C193 _145_ VGND 1.55f
C194 a_12240_11305 VGND 0.736f
C195 a_12415_11231 VGND 0.971f
C196 a_11675_11305 VGND 0.714f
C197 _035_ VGND 1.82f
C198 a_11893_10901 VGND 0.653f
C199 a_11325_10933 VGND 1.57f
C200 _009_ VGND 1.19f
C201 a_11159_10933 VGND 1.92f
C202 a_6904_11305 VGND 0.736f
C203 a_7079_11231 VGND 0.971f
C204 a_6339_11305 VGND 0.714f
C205 _039_ VGND 2.09f
C206 a_6557_10901 VGND 0.653f
C207 a_5989_10933 VGND 1.57f
C208 a_5823_10933 VGND 1.92f
C209 a_4420_11305 VGND 0.736f
C210 a_4595_11231 VGND 1.13f
C211 a_3855_11305 VGND 0.714f
C212 _040_ VGND 1.64f
C213 a_4073_10901 VGND 0.653f
C214 a_3505_10933 VGND 1.57f
C215 _014_ VGND 1.1f
C216 a_3339_10933 VGND 1.92f
C217 a_2703_10927 VGND 0.684f
C218 a_24920_11471 VGND 0.205f
C219 a_27607_11837 VGND 0.168f
C220 a_27404_11471 VGND 0.259f
C221 a_28064_11471 VGND 0.736f
C222 a_28239_11445 VGND 1.13f
C223 a_27499_11471 VGND 0.714f
C224 _048_ VGND 1.66f
C225 a_27717_11713 VGND 0.653f
C226 a_27149_11471 VGND 1.57f
C227 a_26983_11471 VGND 1.92f
C228 _016_ VGND 1.04f
C229 a_21817_11471 VGND 0.23f
C230 a_24694_11517 VGND 0.443f
C231 a_24551_11623 VGND 0.65f
C232 a_22327_11837 VGND 0.609f
C233 a_22495_11739 VGND 0.817f
C234 a_21902_11837 VGND 0.626f
C235 a_22070_11583 VGND 0.581f
C236 a_21629_11471 VGND 1.43f
C237 a_21463_11471 VGND 1.81f
C238 a_19517_11471 VGND 0.23f
C239 a_20819_11471 VGND 0.729f
C240 tdc1.r_ring_ctr10 VGND 3.95f
C241 tdc1.r_ring_ctr9 VGND 5.97f
C242 a_20027_11837 VGND 0.609f
C243 a_20195_11739 VGND 0.817f
C244 a_19602_11837 VGND 0.626f
C245 a_19770_11583 VGND 0.581f
C246 a_19329_11471 VGND 1.43f
C247 tdc1.r_ring_ctr8 VGND 6.84f
C248 a_19163_11471 VGND 1.81f
C249 a_17395_11837 VGND 0.168f
C250 a_17192_11471 VGND 0.259f
C251 a_17852_11471 VGND 0.736f
C252 a_18027_11445 VGND 0.971f
C253 a_17287_11471 VGND 0.714f
C254 _061_ VGND 1.64f
C255 a_17505_11713 VGND 0.653f
C256 a_16937_11471 VGND 1.57f
C257 _020_ VGND 1.24f
C258 a_16771_11471 VGND 1.92f
C259 _625_.X VGND 0.226f
C260 a_16219_11471 VGND 0.648f
C261 _624_.X VGND 0.226f
C262 tdc1.w_dly_stop2 VGND 0.834f
C263 a_9299_11837 VGND 0.168f
C264 a_9096_11471 VGND 0.259f
C265 a_15904_11445 VGND 0.648f
C266 a_15575_11471 VGND 0.524f
C267 tdc1.w_dly_stop1 VGND 0.683f
C268 a_15299_11471 VGND 0.524f
C269 a_14799_11445 VGND 0.698f
C270 a_13603_11445 VGND 0.729f
C271 _146_ VGND 1.29f
C272 a_11763_11445 VGND 0.698f
C273 a_9756_11471 VGND 0.736f
C274 a_9931_11445 VGND 0.971f
C275 a_9191_11471 VGND 0.714f
C276 _037_ VGND 1.6f
C277 a_9409_11713 VGND 0.653f
C278 a_8841_11471 VGND 1.57f
C279 a_8675_11471 VGND 1.92f
C280 _011_ VGND 1.07f
C281 _153_ VGND 0.863f
C282 a_6244_11471 VGND 0.205f
C283 _013_ VGND 1.16f
C284 _151_ VGND 0.958f
C285 a_7815_11623 VGND 0.56f
C286 _150_ VGND 1.22f
C287 a_6607_11623 VGND 0.619f
C288 _152_ VGND 1.82f
C289 a_6018_11517 VGND 0.443f
C290 a_5875_11623 VGND 0.65f
C291 a_5087_11471 VGND 0.988f
C292 _197_ VGND 12.5f
C293 a_29631_12015 VGND 0.168f
C294 a_28529_12015 VGND 0.219f
C295 a_27304_12015 VGND 0.168f
C296 a_29428_12381 VGND 0.259f
C297 a_27722_12015 VGND 0.259f
C298 a_24939_12015 VGND 0.168f
C299 a_24736_12381 VGND 0.259f
C300 _179_ VGND 6.48f
C301 a_21633_12015 VGND 0.23f
C302 a_18051_12015 VGND 0.184f
C303 a_17417_12015 VGND 0.253f
C304 a_19057_12015 VGND 0.23f
C305 _187_ VGND 1.19f
C306 a_14917_12015 VGND 0.23f
C307 a_13445_12015 VGND 0.23f
C308 a_11329_12015 VGND 0.23f
C309 a_4055_12015 VGND 0.168f
C310 a_3852_12381 VGND 0.259f
C311 a_2861_12335 VGND 0.211f
C312 a_30088_12393 VGND 0.736f
C313 a_30263_12319 VGND 1.13f
C314 a_29523_12393 VGND 0.714f
C315 _049_ VGND 1.74f
C316 a_29741_11989 VGND 0.653f
C317 a_29173_12021 VGND 1.57f
C318 _023_ VGND 1.14f
C319 a_29007_12021 VGND 1.92f
C320 a_28279_12015 VGND 0.684f
C321 a_27090_12015 VGND 0.653f
C322 a_27159_11989 VGND 0.714f
C323 a_26964_12131 VGND 1.57f
C324 a_27003_12257 VGND 1.92f
C325 a_26686_12147 VGND 0.736f
C326 a_26483_11989 VGND 0.971f
C327 a_25396_12393 VGND 0.736f
C328 a_25571_12319 VGND 0.971f
C329 a_24831_12393 VGND 0.714f
C330 _055_ VGND 1.74f
C331 a_25049_11989 VGND 0.653f
C332 a_24481_12021 VGND 1.57f
C333 _029_ VGND 1.11f
C334 a_24315_12021 VGND 1.92f
C335 a_23211_12015 VGND 0.698f
C336 a_22143_12015 VGND 0.609f
C337 a_22311_11989 VGND 0.817f
C338 a_21718_12015 VGND 0.626f
C339 a_21886_11989 VGND 0.581f
C340 a_21445_12021 VGND 1.43f
C341 tdc1.r_ring_ctr11 VGND 2.79f
C342 a_21279_12021 VGND 1.81f
C343 a_19567_12015 VGND 0.609f
C344 a_19735_11989 VGND 0.817f
C345 a_19142_12015 VGND 0.626f
C346 a_19310_11989 VGND 0.581f
C347 a_18869_12021 VGND 1.43f
C348 a_18703_12021 VGND 1.81f
C349 a_17586_12335 VGND 0.55f
C350 a_15427_12015 VGND 0.609f
C351 a_15595_11989 VGND 0.817f
C352 a_15002_12015 VGND 0.626f
C353 a_15170_11989 VGND 0.581f
C354 a_14729_12021 VGND 1.43f
C355 tdc0.r_ring_ctr1 VGND 5.19f
C356 a_14563_12021 VGND 1.81f
C357 a_13955_12015 VGND 0.609f
C358 a_14123_11989 VGND 0.817f
C359 a_13530_12015 VGND 0.626f
C360 a_13698_11989 VGND 0.581f
C361 a_13257_12021 VGND 1.43f
C362 tdc0.r_ring_ctr3 VGND 2.57f
C363 a_13091_12021 VGND 1.81f
C364 a_11839_12015 VGND 0.609f
C365 a_12007_11989 VGND 0.817f
C366 a_11414_12015 VGND 0.626f
C367 a_11582_11989 VGND 0.581f
C368 a_11141_12021 VGND 1.43f
C369 tdc0.r_ring_ctr5 VGND 3.34f
C370 a_10975_12021 VGND 1.81f
C371 a_9503_12015 VGND 0.698f
C372 a_9103_12247 VGND 0.56f
C373 a_6987_12247 VGND 0.56f
C374 _155_ VGND 0.842f
C375 a_6059_11989 VGND 0.698f
C376 a_5271_12128 VGND 0.619f
C377 a_4512_12393 VGND 0.736f
C378 a_4687_12319 VGND 0.971f
C379 a_3947_12393 VGND 0.714f
C380 _041_ VGND 1.74f
C381 a_4165_11989 VGND 0.653f
C382 a_3597_12021 VGND 1.57f
C383 _015_ VGND 1.13f
C384 a_3431_12021 VGND 1.92f
C385 a_2623_12335 VGND 0.706f
C386 _157_ VGND 1.06f
C387 a_29723_12925 VGND 0.168f
C388 a_29520_12559 VGND 0.259f
C389 a_30180_12559 VGND 0.736f
C390 a_30355_12533 VGND 0.971f
C391 a_29615_12559 VGND 0.714f
C392 _051_ VGND 1.6f
C393 a_29833_12801 VGND 0.653f
C394 a_29265_12559 VGND 1.57f
C395 a_29099_12559 VGND 1.92f
C396 _025_ VGND 1.15f
C397 _054_ VGND 1.65f
C398 _028_ VGND 2.27f
C399 _178_ VGND 1.1f
C400 a_20707_12925 VGND 0.168f
C401 a_20504_12559 VGND 0.259f
C402 a_25932_12533 VGND 0.648f
C403 _176_ VGND 0.764f
C404 _175_ VGND 1.48f
C405 a_24591_12559 VGND 0.619f
C406 a_23363_12711 VGND 0.56f
C407 _177_ VGND 1.53f
C408 _183_ VGND 2.57f
C409 a_22711_12533 VGND 0.729f
C410 a_22199_12559 VGND 0.619f
C411 a_21164_12559 VGND 0.736f
C412 a_21339_12533 VGND 0.971f
C413 a_20599_12559 VGND 0.714f
C414 a_20817_12801 VGND 0.653f
C415 a_20249_12559 VGND 1.57f
C416 a_20083_12559 VGND 1.92f
C417 a_16475_12925 VGND 0.168f
C418 a_16272_12559 VGND 0.259f
C419 _189_ VGND 0.93f
C420 a_17691_12559 VGND 0.729f
C421 _185_ VGND 5.63f
C422 tdc1.r_ring_ctr13 VGND 3.84f
C423 a_16932_12559 VGND 0.736f
C424 a_17107_12533 VGND 0.971f
C425 a_16367_12559 VGND 0.714f
C426 _062_ VGND 1.66f
C427 a_16585_12801 VGND 0.653f
C428 a_16017_12559 VGND 1.57f
C429 _021_ VGND 1.84f
C430 a_15851_12559 VGND 1.92f
C431 a_12341_12559 VGND 0.23f
C432 a_12851_12925 VGND 0.609f
C433 a_13019_12827 VGND 0.817f
C434 a_12426_12925 VGND 0.626f
C435 a_12594_12671 VGND 0.581f
C436 a_12153_12559 VGND 1.43f
C437 tdc0.r_ring_ctr0 VGND 6.29f
C438 a_11987_12559 VGND 1.81f
C439 a_10869_12559 VGND 0.23f
C440 a_11379_12925 VGND 0.609f
C441 a_11547_12827 VGND 0.817f
C442 a_10954_12925 VGND 0.626f
C443 a_11122_12671 VGND 0.581f
C444 a_10681_12559 VGND 1.43f
C445 tdc0.r_ring_ctr4 VGND 4.66f
C446 a_10515_12559 VGND 1.81f
C447 a_9213_12559 VGND 0.23f
C448 a_9723_12925 VGND 0.609f
C449 a_9891_12827 VGND 0.817f
C450 a_9298_12925 VGND 0.626f
C451 a_9466_12671 VGND 0.581f
C452 a_9025_12559 VGND 1.43f
C453 tdc0.r_ring_ctr6 VGND 4.06f
C454 a_8859_12559 VGND 1.81f
C455 a_7189_12559 VGND 0.23f
C456 a_7699_12925 VGND 0.609f
C457 a_7867_12827 VGND 0.817f
C458 a_7274_12925 VGND 0.626f
C459 a_7442_12671 VGND 0.581f
C460 a_7001_12559 VGND 1.43f
C461 tdc0.r_ring_ctr7 VGND 2.7f
C462 a_6835_12559 VGND 1.81f
C463 a_1129_12809 VGND 0.219f
C464 _147_ VGND 7.79f
C465 _149_ VGND 4.59f
C466 _154_ VGND 2.02f
C467 a_5791_12533 VGND 0.887f
C468 a_3431_12559 VGND 0.729f
C469 _156_ VGND 5.68f
C470 a_2743_12711 VGND 0.619f
C471 _158_ VGND 1.39f
C472 a_1099_12744 VGND 0.684f
C473 a_28731_13103 VGND 0.238f
C474 a_27396_13103 VGND 0.168f
C475 _171_ VGND 1.05f
C476 a_27814_13103 VGND 0.259f
C477 _172_ VGND 3.54f
C478 a_22905_13481 VGND 0.23f
C479 a_19605_13103 VGND 0.219f
C480 _063_ VGND 1.71f
C481 _022_ VGND 1.37f
C482 a_17861_13103 VGND 0.23f
C483 a_14549_13103 VGND 0.23f
C484 a_13077_13103 VGND 0.23f
C485 a_8385_13103 VGND 0.23f
C486 a_6913_13103 VGND 0.23f
C487 _160_ VGND 1.5f
C488 a_4055_13103 VGND 0.168f
C489 a_3852_13469 VGND 0.259f
C490 a_1755_13103 VGND 0.168f
C491 a_1552_13469 VGND 0.259f
C492 _167_ VGND 0.872f
C493 a_27182_13103 VGND 0.653f
C494 a_27251_13077 VGND 0.714f
C495 a_27056_13219 VGND 1.57f
C496 a_27095_13345 VGND 1.92f
C497 _052_ VGND 1.82f
C498 a_26778_13235 VGND 0.736f
C499 a_26575_13077 VGND 0.971f
C500 _198_ VGND 11.7f
C501 _173_ VGND 1.61f
C502 a_24835_13335 VGND 0.56f
C503 a_24347_13441 VGND 0.56f
C504 tdc1.r_ring_ctr6 VGND 3.9f
C505 a_22487_13481 VGND 0.581f
C506 a_22558_13380 VGND 0.626f
C507 a_22358_13225 VGND 1.43f
C508 a_22351_13321 VGND 1.81f
C509 a_22067_13335 VGND 0.609f
C510 a_21971_13335 VGND 0.817f
C511 a_19355_13103 VGND 0.684f
C512 _188_ VGND 2f
C513 a_18371_13103 VGND 0.609f
C514 a_18539_13077 VGND 0.817f
C515 a_17946_13103 VGND 0.626f
C516 a_18114_13077 VGND 0.581f
C517 a_17673_13109 VGND 1.43f
C518 tdc1.r_ring_ctr14 VGND 2.25f
C519 a_17507_13109 VGND 1.81f
C520 a_15059_13103 VGND 0.609f
C521 a_15227_13077 VGND 0.817f
C522 a_14634_13103 VGND 0.626f
C523 a_14802_13077 VGND 0.581f
C524 a_14361_13109 VGND 1.43f
C525 tdc0.w_ring_buf25 VGND 2.08f
C526 a_14195_13109 VGND 1.81f
C527 a_13587_13103 VGND 0.609f
C528 a_13755_13077 VGND 0.817f
C529 a_13162_13103 VGND 0.626f
C530 a_13330_13077 VGND 0.581f
C531 a_12889_13109 VGND 1.43f
C532 tdc0.r_ring_ctr2 VGND 3.6f
C533 a_12723_13109 VGND 1.81f
C534 a_11067_13103 VGND 0.524f
C535 a_8895_13103 VGND 0.609f
C536 a_9063_13077 VGND 0.817f
C537 a_8470_13103 VGND 0.626f
C538 a_8638_13077 VGND 0.581f
C539 a_8197_13109 VGND 1.43f
C540 a_8031_13109 VGND 1.81f
C541 a_7423_13103 VGND 0.609f
C542 a_7591_13077 VGND 0.817f
C543 a_6998_13103 VGND 0.626f
C544 a_7166_13077 VGND 0.581f
C545 a_6725_13109 VGND 1.43f
C546 a_6559_13109 VGND 1.81f
C547 tdc0.r_ring_ctr8 VGND 6.51f
C548 tdc0.r_ring_ctr9 VGND 5.93f
C549 a_5875_13077 VGND 0.729f
C550 a_4512_13481 VGND 0.736f
C551 a_4687_13407 VGND 0.971f
C552 a_3947_13481 VGND 0.714f
C553 _043_ VGND 1.82f
C554 a_4165_13077 VGND 0.653f
C555 a_3597_13109 VGND 1.57f
C556 a_3431_13109 VGND 1.92f
C557 a_2212_13481 VGND 0.736f
C558 a_2387_13407 VGND 0.971f
C559 a_1647_13481 VGND 0.714f
C560 _042_ VGND 1.6f
C561 a_1865_13077 VGND 0.653f
C562 a_1297_13109 VGND 1.57f
C563 _001_ VGND 1.35f
C564 a_1131_13109 VGND 1.92f
C565 a_29815_14013 VGND 0.168f
C566 a_29612_13647 VGND 0.259f
C567 a_30272_13647 VGND 0.736f
C568 a_30447_13621 VGND 0.971f
C569 a_29707_13647 VGND 0.714f
C570 _050_ VGND 1.66f
C571 a_29925_13889 VGND 0.653f
C572 a_29357_13647 VGND 1.57f
C573 _024_ VGND 1.08f
C574 a_29191_13647 VGND 1.92f
C575 _168_ VGND 1.43f
C576 a_24939_14013 VGND 0.168f
C577 a_24736_13647 VGND 0.259f
C578 a_28455_13647 VGND 0.619f
C579 a_26615_13647 VGND 0.698f
C580 a_25396_13647 VGND 0.736f
C581 a_25571_13621 VGND 0.971f
C582 a_24831_13647 VGND 0.714f
C583 _053_ VGND 1.61f
C584 a_25049_13889 VGND 0.653f
C585 a_24481_13647 VGND 1.57f
C586 _027_ VGND 1.46f
C587 a_24315_13647 VGND 1.92f
C588 net10 VGND 9.17f
C589 _174_ VGND 1.37f
C590 a_23947_13897 VGND 0.238f
C591 a_22553_13647 VGND 0.23f
C592 a_23063_14013 VGND 0.609f
C593 a_23231_13915 VGND 0.817f
C594 a_22638_14013 VGND 0.626f
C595 a_22806_13759 VGND 0.581f
C596 a_22365_13647 VGND 1.43f
C597 tdc1.r_ring_ctr15 VGND 2.94f
C598 a_22199_13647 VGND 1.81f
C599 a_20717_13897 VGND 0.206f
C600 a_17217_13647 VGND 0.23f
C601 a_20635_13897 VGND 0.804f
C602 tdc1.r_dly_store_ctr8 VGND 1.45f
C603 a_17727_14013 VGND 0.609f
C604 a_17895_13915 VGND 0.817f
C605 a_17302_14013 VGND 0.626f
C606 a_17470_13759 VGND 0.581f
C607 a_17029_13647 VGND 1.43f
C608 tdc1.r_ring_ctr12 VGND 5.25f
C609 a_16863_13647 VGND 1.81f
C610 a_15009_13647 VGND 0.23f
C611 a_15519_14013 VGND 0.609f
C612 a_15687_13915 VGND 0.817f
C613 a_15094_14013 VGND 0.626f
C614 a_15262_13759 VGND 0.581f
C615 a_14821_13647 VGND 1.43f
C616 a_14655_13647 VGND 1.81f
C617 tdc0.w_ring_buf9 VGND 0.984f
C618 a_11697_13647 VGND 0.23f
C619 a_14195_13647 VGND 0.524f
C620 a_12207_14013 VGND 0.609f
C621 a_12375_13915 VGND 0.817f
C622 a_11782_14013 VGND 0.626f
C623 a_11950_13759 VGND 0.581f
C624 a_11509_13647 VGND 1.43f
C625 a_11343_13647 VGND 1.81f
C626 tdc0.w_ring_int_norsz25 VGND 0.722f
C627 net54 VGND 0.822f
C628 tdc0.g_ring325.stg01_54.HI VGND 0.415f
C629 tdc0.g_ring327.stg01_56.HI VGND 0.415f
C630 tdc0.w_ring_norsz25 VGND 2.58f
C631 a_4069_13647 VGND 0.171f
C632 a_5993_13647 VGND 0.23f
C633 a_6503_14013 VGND 0.609f
C634 a_6671_13915 VGND 0.817f
C635 a_6078_14013 VGND 0.626f
C636 a_6246_13759 VGND 0.581f
C637 a_5805_13647 VGND 1.43f
C638 tdc0.r_ring_ctr10 VGND 4.82f
C639 a_5639_13647 VGND 1.81f
C640 _002_ VGND 1.09f
C641 a_1113_13897 VGND 0.219f
C642 _159_ VGND 1.15f
C643 a_3851_13621 VGND 0.546f
C644 a_863_13897 VGND 0.684f
C645 a_26689_14191 VGND 0.219f
C646 a_30281_14191 VGND 0.23f
C647 _026_ VGND 1.77f
C648 a_25297_14569 VGND 0.23f
C649 a_22281_14191 VGND 0.206f
C650 a_21768_14191 VGND 0.259f
C651 tdc1.r_dly_store_ring24 VGND 0.969f
C652 a_19609_14191 VGND 0.23f
C653 a_13817_14191 VGND 0.206f
C654 a_13173_14191 VGND 0.206f
C655 a_12529_14191 VGND 0.206f
C656 a_16481_14191 VGND 0.23f
C657 tdc0.w_ring_int_norsz9 VGND 1.08f
C658 tdc0.w_ring_buf24 VGND 1.08f
C659 a_30791_14191 VGND 0.609f
C660 a_30959_14165 VGND 0.817f
C661 a_30366_14191 VGND 0.626f
C662 a_30534_14165 VGND 0.581f
C663 a_30093_14197 VGND 1.43f
C664 a_29927_14197 VGND 1.81f
C665 _169_ VGND 0.702f
C666 a_29519_14165 VGND 0.698f
C667 a_28823_14557 VGND 0.729f
C668 tdc1.r_ring_ctr3 VGND 3.29f
C669 a_26439_14191 VGND 0.684f
C670 _170_ VGND 8.64f
C671 tdc1.r_ring_ctr4 VGND 4.39f
C672 a_24879_14569 VGND 0.581f
C673 a_24950_14468 VGND 0.626f
C674 a_24750_14313 VGND 1.43f
C675 a_24743_14409 VGND 1.81f
C676 a_24459_14423 VGND 0.609f
C677 a_24363_14423 VGND 0.817f
C678 tdc1.r_dly_store_ctr11 VGND 1.43f
C679 tdc1.r_dly_store_ctr3 VGND 4.38f
C680 a_22135_14423 VGND 0.804f
C681 _193_ VGND 1.04f
C682 a_21337_14165 VGND 0.672f
C683 a_20119_14191 VGND 0.609f
C684 a_20287_14165 VGND 0.817f
C685 a_19694_14191 VGND 0.626f
C686 a_19862_14165 VGND 0.581f
C687 a_19421_14197 VGND 1.43f
C688 tdc1.w_ring_buf24 VGND 0.872f
C689 a_19255_14197 VGND 1.81f
C690 a_18979_14191 VGND 0.524f
C691 a_16991_14191 VGND 0.609f
C692 a_17159_14165 VGND 0.817f
C693 a_16566_14191 VGND 0.626f
C694 a_16734_14165 VGND 0.581f
C695 a_16293_14197 VGND 1.43f
C696 tdc0.w_ring_buf8 VGND 1.03f
C697 a_16127_14197 VGND 1.81f
C698 a_15483_14191 VGND 0.524f
C699 a_13735_14191 VGND 0.804f
C700 tdc0.r_dly_store_ctr2 VGND 1.09f
C701 tdc0.r_dly_store_ctr10 VGND 4.06f
C702 a_13091_14191 VGND 0.804f
C703 a_12447_14191 VGND 0.804f
C704 tdc0.r_dly_store_ring24 VGND 0.833f
C705 tdc0.r_dly_store_ctr8 VGND 3.14f
C706 a_11159_14191 VGND 0.524f
C707 tdc0.w_ring_norsz9 VGND 3.5f
C708 tdc0.g_ring326.stg01_55.HI VGND 0.415f
C709 net55 VGND 1.26f
C710 tdc0.r_dly_store_ring27 VGND 2.59f
C711 a_7925_14191 VGND 0.23f
C712 tdc0.r_dly_store_ctr11 VGND 3.31f
C713 a_6177_14191 VGND 0.23f
C714 a_3701_14511 VGND 0.171f
C715 a_1755_14191 VGND 0.168f
C716 a_1552_14557 VGND 0.259f
C717 tdc0.w_ring_int_norsz10 VGND 0.839f
C718 tdc0.w_ring_int_norsz26 VGND 0.878f
C719 a_9227_14191 VGND 0.524f
C720 a_8435_14191 VGND 0.609f
C721 a_8603_14165 VGND 0.817f
C722 a_8010_14191 VGND 0.626f
C723 a_8178_14165 VGND 0.581f
C724 a_7737_14197 VGND 1.43f
C725 a_7571_14197 VGND 1.81f
C726 a_6687_14191 VGND 0.609f
C727 a_6855_14165 VGND 0.817f
C728 a_6262_14191 VGND 0.626f
C729 a_6430_14165 VGND 0.581f
C730 a_5989_14197 VGND 1.43f
C731 tdc0.r_ring_ctr11 VGND 2.87f
C732 a_5823_14197 VGND 1.81f
C733 _161_ VGND 2.35f
C734 a_3483_14423 VGND 0.546f
C735 a_2212_14569 VGND 0.736f
C736 a_2387_14495 VGND 1.13f
C737 a_1647_14569 VGND 0.714f
C738 _044_ VGND 1.64f
C739 a_1865_14165 VGND 0.653f
C740 a_1297_14197 VGND 1.57f
C741 _003_ VGND 1.15f
C742 a_1131_14197 VGND 1.92f
C743 a_28241_14735 VGND 0.23f
C744 a_26141_14735 VGND 0.23f
C745 tdc1.r_ring_ctr0 VGND 5.92f
C746 a_27823_14735 VGND 0.581f
C747 a_27894_14709 VGND 0.626f
C748 a_27687_14709 VGND 1.81f
C749 a_27694_15009 VGND 1.43f
C750 a_27403_14709 VGND 0.609f
C751 a_27307_14887 VGND 0.817f
C752 a_26651_15101 VGND 0.609f
C753 a_26819_15003 VGND 0.817f
C754 a_26226_15101 VGND 0.626f
C755 a_26394_14847 VGND 0.581f
C756 a_25953_14735 VGND 1.43f
C757 tdc1.r_ring_ctr5 VGND 3.27f
C758 a_25787_14735 VGND 1.81f
C759 a_24209_14735 VGND 0.23f
C760 a_24719_15101 VGND 0.609f
C761 a_24887_15003 VGND 0.817f
C762 a_24294_15101 VGND 0.626f
C763 a_24462_14847 VGND 0.581f
C764 a_24021_14735 VGND 1.43f
C765 tdc1.r_ring_ctr7 VGND 4.44f
C766 a_23855_14735 VGND 1.81f
C767 a_23211_14735 VGND 0.648f
C768 a_22741_14985 VGND 0.206f
C769 _195_ VGND 1.34f
C770 tdc1.r_dly_store_ring8 VGND 0.902f
C771 a_20713_14735 VGND 0.23f
C772 tdc1.r_dly_store_ctr0 VGND 2.59f
C773 a_22595_14887 VGND 0.804f
C774 a_21223_15101 VGND 0.609f
C775 a_21391_15003 VGND 0.817f
C776 a_20798_15101 VGND 0.626f
C777 a_20966_14847 VGND 0.581f
C778 a_20525_14735 VGND 1.43f
C779 a_20359_14735 VGND 1.81f
C780 tdc1.w_ring_buf8 VGND 0.872f
C781 a_18869_14985 VGND 0.214f
C782 a_18785_14985 VGND 0.167f
C783 a_17213_14985 VGND 0.214f
C784 a_17129_14985 VGND 0.167f
C785 a_15929_14735 VGND 0.23f
C786 a_20083_14735 VGND 0.524f
C787 a_18703_14735 VGND 0.972f
C788 tdc1.r_dly_store_ctr6 VGND 2.42f
C789 tdc1.r_dly_store_ctr14 VGND 1.2f
C790 a_17047_14735 VGND 0.972f
C791 tdc0.r_dly_store_ring8 VGND 0.815f
C792 tdc0.r_dly_store_ring0 VGND 0.668f
C793 a_16439_15101 VGND 0.609f
C794 a_16607_15003 VGND 0.817f
C795 a_16014_15101 VGND 0.626f
C796 a_16182_14847 VGND 0.581f
C797 a_15741_14735 VGND 1.43f
C798 net8 VGND 9.97f
C799 a_15575_14735 VGND 1.81f
C800 _094_ VGND 1.15f
C801 a_14545_14985 VGND 0.214f
C802 a_14461_14985 VGND 0.167f
C803 a_13717_14985 VGND 0.214f
C804 a_13633_14985 VGND 0.167f
C805 a_11237_14735 VGND 0.23f
C806 a_15117_14741 VGND 0.665f
C807 a_14379_14735 VGND 0.972f
C808 tdc0.r_dly_store_ctr3 VGND 1.74f
C809 _101_ VGND 1.08f
C810 a_13551_14735 VGND 0.972f
C811 tdc0.r_dly_store_ctr0 VGND 1.65f
C812 _190_ VGND 0.996f
C813 a_11747_15101 VGND 0.609f
C814 a_11915_15003 VGND 0.817f
C815 a_11322_15101 VGND 0.626f
C816 a_11490_14847 VGND 0.581f
C817 a_11049_14735 VGND 1.43f
C818 tdc0.w_ring_buf26 VGND 1.65f
C819 a_10883_14735 VGND 1.81f
C820 a_9765_14735 VGND 0.23f
C821 a_10275_15101 VGND 0.609f
C822 a_10443_15003 VGND 0.817f
C823 a_9850_15101 VGND 0.626f
C824 a_10018_14847 VGND 0.581f
C825 a_9577_14735 VGND 1.43f
C826 a_9411_14735 VGND 1.81f
C827 tdc0.w_ring_buf10 VGND 0.872f
C828 tdc0.w_ring_buf27 VGND 1.06f
C829 tdc0.r_dly_store_ring16 VGND 3.71f
C830 a_5809_14735 VGND 0.23f
C831 a_9135_14735 VGND 0.524f
C832 tdc0.w_ring_norsz10 VGND 2.16f
C833 tdc0.w_ring_int_norsz27 VGND 0.956f
C834 tdc0.w_ring_int_norsz11 VGND 1.01f
C835 net56 VGND 1.51f
C836 tdc0.w_ring_norsz26 VGND 2.95f
C837 a_7295_14735 VGND 0.524f
C838 a_6319_15101 VGND 0.609f
C839 a_6487_15003 VGND 0.817f
C840 a_5894_15101 VGND 0.626f
C841 a_6062_14847 VGND 0.581f
C842 a_5621_14735 VGND 1.43f
C843 a_5455_14735 VGND 1.81f
C844 a_3963_15101 VGND 0.168f
C845 a_3760_14735 VGND 0.259f
C846 a_4420_14735 VGND 0.736f
C847 a_4595_14709 VGND 0.971f
C848 a_3855_14735 VGND 0.714f
C849 _045_ VGND 1.66f
C850 a_4073_14977 VGND 0.653f
C851 a_3505_14735 VGND 1.57f
C852 _004_ VGND 1.13f
C853 a_3339_14735 VGND 1.92f
C854 _163_ VGND 1.22f
C855 a_30281_15279 VGND 0.23f
C856 _627_.X VGND 0.226f
C857 a_28977_15657 VGND 0.23f
C858 a_25849_15657 VGND 0.23f
C859 a_23937_15279 VGND 0.206f
C860 tdc1.r_dly_store_ring16 VGND 1.61f
C861 a_30791_15279 VGND 0.609f
C862 a_30959_15253 VGND 0.817f
C863 a_30366_15279 VGND 0.626f
C864 a_30534_15253 VGND 0.581f
C865 a_30093_15285 VGND 1.43f
C866 tdc1.r_ring_ctr2 VGND 4.31f
C867 a_29927_15285 VGND 1.81f
C868 a_29467_15287 VGND 0.648f
C869 tdc1.r_ring_ctr1 VGND 4.97f
C870 a_28559_15657 VGND 0.581f
C871 a_28630_15556 VGND 0.626f
C872 a_28430_15401 VGND 1.43f
C873 a_28423_15497 VGND 1.81f
C874 a_28139_15511 VGND 0.609f
C875 a_28043_15511 VGND 0.817f
C876 a_26983_15279 VGND 0.524f
C877 a_25431_15657 VGND 0.581f
C878 a_25502_15556 VGND 0.626f
C879 a_25302_15401 VGND 1.43f
C880 a_25295_15497 VGND 1.81f
C881 a_25011_15511 VGND 0.609f
C882 a_24915_15511 VGND 0.817f
C883 a_23855_15279 VGND 0.804f
C884 tdc1.r_dly_store_ctr7 VGND 1.33f
C885 tdc1.r_dly_store_ctr15 VGND 1.34f
C886 a_22293_15395 VGND 0.665f
C887 _107_ VGND 1.12f
C888 a_18072_15279 VGND 0.14f
C889 a_17720_15279 VGND 0.171f
C890 a_14197_15279 VGND 0.253f
C891 a_13633_15279 VGND 0.206f
C892 a_13195_15279 VGND 0.167f
C893 a_12993_15279 VGND 0.214f
C894 a_19241_15279 VGND 0.23f
C895 a_17638_15599 VGND 0.482f
C896 a_16941_15279 VGND 0.227f
C897 _092_ VGND 1.24f
C898 _093_ VGND 1.36f
C899 tdc0.r_dly_store_ring19 VGND 1.82f
C900 a_11329_15279 VGND 0.23f
C901 a_8477_15279 VGND 0.23f
C902 a_21311_15617 VGND 0.56f
C903 a_19751_15279 VGND 0.609f
C904 a_19919_15253 VGND 0.817f
C905 a_19326_15279 VGND 0.626f
C906 a_19494_15253 VGND 0.581f
C907 a_19053_15285 VGND 1.43f
C908 net9 VGND 16.2f
C909 a_18887_15285 VGND 1.81f
C910 net33 VGND 12.6f
C911 a_17804_15279 VGND 1.37f
C912 _196_ VGND 2.59f
C913 _192_ VGND 0.963f
C914 _191_ VGND 2.73f
C915 a_16764_15279 VGND 0.498f
C916 a_16658_15279 VGND 0.578f
C917 a_16481_15279 VGND 0.5f
C918 net30 VGND 7.31f
C919 a_16162_15279 VGND 0.535f
C920 a_14366_15599 VGND 0.55f
C921 a_13551_15279 VGND 0.804f
C922 tdc0.r_dly_store_ring26 VGND 1.5f
C923 tdc0.r_dly_store_ring10 VGND 2.04f
C924 tdc0.r_dly_store_ctr6 VGND 3.2f
C925 a_12867_15511 VGND 0.972f
C926 a_11839_15279 VGND 0.609f
C927 a_12007_15253 VGND 0.817f
C928 a_11414_15279 VGND 0.626f
C929 a_11582_15253 VGND 0.581f
C930 a_11141_15285 VGND 1.43f
C931 tdc0.w_ring_buf19 VGND 0.95f
C932 a_10975_15285 VGND 1.81f
C933 a_10515_15279 VGND 0.524f
C934 a_9647_15253 VGND 0.698f
C935 a_8987_15279 VGND 0.609f
C936 a_9155_15253 VGND 0.817f
C937 a_8562_15279 VGND 0.626f
C938 a_8730_15253 VGND 0.581f
C939 a_8289_15285 VGND 1.43f
C940 tdc0.w_ring_buf11 VGND 0.872f
C941 a_8123_15285 VGND 1.81f
C942 a_7847_15279 VGND 0.524f
C943 tdc0.g_ring328.stg01_57.HI VGND 0.415f
C944 a_3703_15279 VGND 0.253f
C945 a_2227_15279 VGND 0.184f
C946 tdc0.w_ring_buf16 VGND 1.39f
C947 _164_ VGND 1.04f
C948 net57 VGND 0.822f
C949 tdc0.w_ring_norsz27 VGND 2.48f
C950 a_5363_15279 VGND 0.524f
C951 a_5087_15279 VGND 0.524f
C952 a_3485_15253 VGND 0.55f
C953 _162_ VGND 6.09f
C954 a_1551_15253 VGND 0.729f
C955 a_29989_15823 VGND 0.23f
C956 tdc1.w_ring_buf12 VGND 1.46f
C957 a_29571_15823 VGND 0.581f
C958 a_29642_15797 VGND 0.626f
C959 a_29435_15797 VGND 1.81f
C960 a_29442_16097 VGND 1.43f
C961 a_29151_15797 VGND 0.609f
C962 a_29055_15975 VGND 0.817f
C963 a_28599_15797 VGND 0.698f
C964 a_28271_15823 VGND 0.524f
C965 a_27689_15823 VGND 0.23f
C966 a_24485_15823 VGND 0.23f
C967 tdc1.w_ring_buf27 VGND 1.19f
C968 a_27271_15823 VGND 0.581f
C969 a_27342_15797 VGND 0.626f
C970 a_27135_15797 VGND 1.81f
C971 a_27142_16097 VGND 1.43f
C972 a_26851_15797 VGND 0.609f
C973 a_26755_15975 VGND 0.817f
C974 a_24995_16189 VGND 0.609f
C975 a_25163_16091 VGND 0.817f
C976 a_24570_16189 VGND 0.626f
C977 a_24738_15935 VGND 0.581f
C978 a_24297_15823 VGND 1.43f
C979 a_24131_15823 VGND 1.81f
C980 net36 VGND 10.4f
C981 a_23201_16073 VGND 0.206f
C982 a_22671_16073 VGND 0.167f
C983 a_22469_16073 VGND 0.214f
C984 _194_ VGND 1.44f
C985 a_15027_15823 VGND 0.319f
C986 tdc1.r_dly_store_ring0 VGND 1.11f
C987 a_20175_16073 VGND 0.333f
C988 tdc1.r_dly_store_ring12 VGND 3.16f
C989 tdc1.r_dly_store_ctr4 VGND 1.65f
C990 a_23055_15975 VGND 0.804f
C991 tdc1.r_dly_store_ctr9 VGND 2.25f
C992 tdc1.r_dly_store_ctr1 VGND 3.38f
C993 a_22343_15975 VGND 0.972f
C994 a_21463_15823 VGND 0.988f
C995 _088_ VGND 0.89f
C996 a_20911_15823 VGND 0.619f
C997 a_20258_16073 VGND 0.723f
C998 tdc1.r_dly_store_ctr13 VGND 2.48f
C999 a_18239_16073 VGND 0.253f
C1000 a_19860_15797 VGND 0.648f
C1001 tdc1.r_dly_store_ctr12 VGND 1.47f
C1002 a_18021_15797 VGND 0.55f
C1003 a_17043_16073 VGND 0.253f
C1004 a_16301_16073 VGND 0.206f
C1005 a_13993_16073 VGND 0.214f
C1006 a_13909_16073 VGND 0.167f
C1007 a_12889_16073 VGND 0.214f
C1008 a_12805_16073 VGND 0.167f
C1009 a_12161_16073 VGND 0.206f
C1010 a_10593_15823 VGND 0.23f
C1011 a_17468_15797 VGND 0.648f
C1012 tdc0.r_dly_store_ring9 VGND 1.89f
C1013 a_16825_15797 VGND 0.55f
C1014 tdc0.r_dly_store_ring25 VGND 2.1f
C1015 tdc0.r_dly_store_ctr1 VGND 2.28f
C1016 a_16155_15975 VGND 0.804f
C1017 a_15196_16073 VGND 1.33f
C1018 _108_ VGND 4.13f
C1019 _103_ VGND 1.06f
C1020 _102_ VGND 1.56f
C1021 a_13827_15823 VGND 0.972f
C1022 tdc0.r_dly_store_ring11 VGND 2.88f
C1023 tdc0.r_dly_store_ring3 VGND 1.56f
C1024 a_12723_15823 VGND 0.972f
C1025 _079_ VGND 10.7f
C1026 tdc0.r_dly_store_ctr5 VGND 2.36f
C1027 _118_ VGND 0.621f
C1028 a_12079_16073 VGND 0.804f
C1029 _080_ VGND 12.1f
C1030 a_11103_16189 VGND 0.609f
C1031 a_11271_16091 VGND 0.817f
C1032 a_10678_16189 VGND 0.626f
C1033 a_10846_15935 VGND 0.581f
C1034 a_10405_15823 VGND 1.43f
C1035 a_10239_15823 VGND 1.81f
C1036 net29 VGND 9.32f
C1037 tdc0.r_dly_store_ring21 VGND 1.75f
C1038 a_9121_15823 VGND 0.23f
C1039 a_9631_16189 VGND 0.609f
C1040 a_9799_16091 VGND 0.817f
C1041 a_9206_16189 VGND 0.626f
C1042 a_9374_15935 VGND 0.581f
C1043 a_8933_15823 VGND 1.43f
C1044 a_8767_15823 VGND 1.81f
C1045 tdc0.r_dly_store_ring29 VGND 2.68f
C1046 a_6913_15823 VGND 0.23f
C1047 tdc0.w_ring_norsz11 VGND 2.46f
C1048 a_7423_16189 VGND 0.609f
C1049 a_7591_16091 VGND 0.817f
C1050 a_6998_16189 VGND 0.626f
C1051 a_7166_15935 VGND 0.581f
C1052 a_6725_15823 VGND 1.43f
C1053 a_6559_15823 VGND 1.81f
C1054 tdc0.r_dly_store_ctr13 VGND 3.01f
C1055 a_5349_15823 VGND 0.23f
C1056 a_5859_16189 VGND 0.609f
C1057 a_6027_16091 VGND 0.817f
C1058 a_5434_16189 VGND 0.626f
C1059 a_5602_15935 VGND 0.581f
C1060 a_5161_15823 VGND 1.43f
C1061 tdc0.r_ring_ctr13 VGND 4.44f
C1062 a_4995_15823 VGND 1.81f
C1063 tdc0.r_dly_store_ctr14 VGND 4.81f
C1064 a_3693_15823 VGND 0.23f
C1065 a_4203_16189 VGND 0.609f
C1066 a_4371_16091 VGND 0.817f
C1067 a_3778_16189 VGND 0.626f
C1068 a_3946_15935 VGND 0.581f
C1069 a_3505_15823 VGND 1.43f
C1070 a_3339_15823 VGND 1.81f
C1071 net26 VGND 10.6f
C1072 tdc0.r_ring_ctr14 VGND 2.4f
C1073 a_1939_16189 VGND 0.168f
C1074 a_1736_15823 VGND 0.259f
C1075 a_2396_15823 VGND 0.736f
C1076 a_2571_15797 VGND 0.971f
C1077 a_1831_15823 VGND 0.714f
C1078 a_2049_16065 VGND 0.653f
C1079 a_1481_15823 VGND 1.57f
C1080 a_1315_15823 VGND 1.92f
C1081 _005_ VGND 1.07f
C1082 _166_ VGND 1.3f
C1083 a_30281_16367 VGND 0.23f
C1084 a_30791_16367 VGND 0.609f
C1085 a_30959_16341 VGND 0.817f
C1086 a_30366_16367 VGND 0.626f
C1087 a_30534_16341 VGND 0.581f
C1088 a_30093_16373 VGND 1.43f
C1089 a_29927_16373 VGND 1.81f
C1090 net75 VGND 1.01f
C1091 tdc1.w_ring_int_norsz28 VGND 0.722f
C1092 tdc1.g_ring328.stg01_75.HI VGND 0.415f
C1093 a_28135_16586 VGND 0.524f
C1094 a_27772_16341 VGND 0.648f
C1095 tdc1.w_ring_norsz27 VGND 3.06f
C1096 tdc1.w_ring_norsz11 VGND 2.8f
C1097 tdc1.w_ring_int_norsz27 VGND 0.722f
C1098 net74 VGND 0.963f
C1099 a_25431_16367 VGND 0.167f
C1100 a_25229_16367 VGND 0.214f
C1101 tdc1.g_ring327.stg01_74.HI VGND 0.415f
C1102 tdc1.r_dly_store_ctr10 VGND 3.04f
C1103 a_22741_16367 VGND 0.234f
C1104 a_25839_16341 VGND 0.698f
C1105 tdc1.r_dly_store_ring26 VGND 0.802f
C1106 tdc1.r_dly_store_ctr2 VGND 4.12f
C1107 a_25103_16599 VGND 0.972f
C1108 a_24467_16599 VGND 0.56f
C1109 _098_ VGND 0.933f
C1110 _096_ VGND 0.763f
C1111 a_21729_16367 VGND 0.206f
C1112 tdc1.w_ring_buf26 VGND 1.23f
C1113 _105_ VGND 1.11f
C1114 _106_ VGND 1.25f
C1115 tdc1.r_dly_store_ring5 VGND 0.967f
C1116 a_18049_16367 VGND 0.206f
C1117 a_19149_16367 VGND 0.23f
C1118 a_16757_16367 VGND 0.23f
C1119 a_23996_16599 VGND 0.665f
C1120 a_23671_16367 VGND 0.524f
C1121 a_22615_16599 VGND 0.953f
C1122 a_21647_16367 VGND 0.804f
C1123 tdc1.r_dly_store_ring27 VGND 3.46f
C1124 a_19659_16367 VGND 0.609f
C1125 a_19827_16341 VGND 0.817f
C1126 a_19234_16367 VGND 0.626f
C1127 a_19402_16341 VGND 0.581f
C1128 a_18961_16373 VGND 1.43f
C1129 a_18795_16373 VGND 1.81f
C1130 tdc1.r_dly_store_ring20 VGND 0.867f
C1131 tdc1.r_dly_store_ring28 VGND 6.47f
C1132 a_17903_16599 VGND 0.804f
C1133 a_17267_16367 VGND 0.609f
C1134 a_17435_16341 VGND 0.817f
C1135 a_16842_16367 VGND 0.626f
C1136 a_17010_16341 VGND 0.581f
C1137 a_16569_16373 VGND 1.43f
C1138 a_16403_16373 VGND 1.81f
C1139 a_15577_16483 VGND 0.665f
C1140 _070_ VGND 1.03f
C1141 _077_ VGND 1.39f
C1142 a_12989_16367 VGND 0.206f
C1143 _073_ VGND 1.64f
C1144 a_14623_16627 VGND 1.2f
C1145 a_13583_16705 VGND 0.56f
C1146 a_12907_16367 VGND 0.804f
C1147 tdc0.r_dly_store_ctr9 VGND 3.7f
C1148 tdc0.g_ring319.stg01_48.HI VGND 0.415f
C1149 tdc0.w_ring_buf3 VGND 1.18f
C1150 tdc0.r_dly_store_ctr12 VGND 4.68f
C1151 a_1297_16367 VGND 0.219f
C1152 a_3877_16367 VGND 0.23f
C1153 _046_ VGND 1.69f
C1154 net48 VGND 0.939f
C1155 a_10147_16367 VGND 0.524f
C1156 tdc0.w_ring_int_norsz12 VGND 0.962f
C1157 tdc0.w_ring_int_norsz28 VGND 1.14f
C1158 a_4387_16367 VGND 0.609f
C1159 a_4555_16341 VGND 0.817f
C1160 a_3962_16367 VGND 0.626f
C1161 a_4130_16341 VGND 0.581f
C1162 a_3689_16373 VGND 1.43f
C1163 tdc0.r_ring_ctr12 VGND 5.83f
C1164 a_3523_16373 VGND 1.81f
C1165 a_1047_16367 VGND 0.684f
C1166 _165_ VGND 1.89f
C1167 tdc1.g_ring329.stg01_76.HI VGND 0.415f
C1168 tdc1.w_ring_buf28 VGND 1.02f
C1169 a_29743_16911 VGND 0.524f
C1170 tdc1.w_ring_int_norsz12 VGND 1.01f
C1171 a_28425_16911 VGND 0.23f
C1172 tdc1.w_ring_int_norsz11 VGND 1.06f
C1173 a_24631_16891 VGND 0.454f
C1174 tdc1.w_ring_buf11 VGND 1.11f
C1175 a_28007_16911 VGND 0.581f
C1176 a_28078_16885 VGND 0.626f
C1177 a_27871_16885 VGND 1.81f
C1178 a_27878_17185 VGND 1.43f
C1179 a_27587_16885 VGND 0.609f
C1180 a_27491_17063 VGND 0.817f
C1181 tdc1.w_dly_stop5 VGND 12f
C1182 a_27127_16885 VGND 0.698f
C1183 a_26031_16885 VGND 1.2f
C1184 tdc1.r_dly_store_ring3 VGND 0.848f
C1185 a_22093_16911 VGND 0.23f
C1186 a_24275_16885 VGND 0.753f
C1187 a_22603_17277 VGND 0.609f
C1188 a_22771_17179 VGND 0.817f
C1189 a_22178_17277 VGND 0.626f
C1190 a_22346_17023 VGND 0.581f
C1191 a_21905_16911 VGND 1.43f
C1192 a_21739_16911 VGND 1.81f
C1193 tdc1.r_dly_store_ring19 VGND 0.765f
C1194 a_20621_16911 VGND 0.23f
C1195 a_21131_17277 VGND 0.609f
C1196 a_21299_17179 VGND 0.817f
C1197 a_20706_17277 VGND 0.626f
C1198 a_20874_17023 VGND 0.581f
C1199 a_20433_16911 VGND 1.43f
C1200 a_20267_16911 VGND 1.81f
C1201 tdc1.w_ring_buf19 VGND 0.872f
C1202 tdc1.w_ring_buf5 VGND 1.03f
C1203 a_18877_17161 VGND 0.206f
C1204 _133_ VGND 1.42f
C1205 a_17478_16911 VGND 0.161f
C1206 a_17126_16911 VGND 0.123f
C1207 _111_ VGND 1.37f
C1208 _109_ VGND 1.1f
C1209 tdc1.w_ring_buf20 VGND 1.65f
C1210 _110_ VGND 3.65f
C1211 a_17044_17161 VGND 0.537f
C1212 a_14300_16911 VGND 0.123f
C1213 a_13948_16911 VGND 0.161f
C1214 a_19991_16911 VGND 0.524f
C1215 a_19395_17076 VGND 0.524f
C1216 a_18731_17063 VGND 0.804f
C1217 a_18383_17076 VGND 0.524f
C1218 a_17924_17063 VGND 0.665f
C1219 _095_ VGND 2.54f
C1220 _099_ VGND 4.02f
C1221 a_16656_16885 VGND 1.37f
C1222 a_16097_16911 VGND 0.23f
C1223 a_13861_17161 VGND 0.537f
C1224 a_12805_17161 VGND 0.206f
C1225 tdc0.r_dly_store_ring18 VGND 2.25f
C1226 a_11329_16911 VGND 0.23f
C1227 a_15679_16911 VGND 0.581f
C1228 a_15750_16885 VGND 0.626f
C1229 a_15543_16885 VGND 1.81f
C1230 a_15550_17185 VGND 1.43f
C1231 a_15259_16885 VGND 0.609f
C1232 a_15163_17063 VGND 0.817f
C1233 a_14032_16911 VGND 1.37f
C1234 _112_ VGND 2.35f
C1235 a_12723_17161 VGND 0.804f
C1236 tdc0.r_dly_store_ctr4 VGND 2.86f
C1237 _069_ VGND 12.3f
C1238 a_11839_17277 VGND 0.609f
C1239 a_12007_17179 VGND 0.817f
C1240 a_11414_17277 VGND 0.626f
C1241 a_11582_17023 VGND 0.581f
C1242 a_11141_16911 VGND 1.43f
C1243 a_10975_16911 VGND 1.81f
C1244 tdc0.w_ring_buf18 VGND 0.872f
C1245 tdc0.r_dly_store_ring28 VGND 1.95f
C1246 a_8753_16911 VGND 0.23f
C1247 a_10699_16911 VGND 0.524f
C1248 tdc0.w_ring_int_norsz19 VGND 1.06f
C1249 a_9263_17277 VGND 0.609f
C1250 a_9431_17179 VGND 0.817f
C1251 a_8838_17277 VGND 0.626f
C1252 a_9006_17023 VGND 0.581f
C1253 a_8565_16911 VGND 1.43f
C1254 a_8399_16911 VGND 1.81f
C1255 tdc0.w_ring_buf28 VGND 1.11f
C1256 tdc0.w_ring_buf29 VGND 1.3f
C1257 tdc0.r_dly_store_ring17 VGND 3.9f
C1258 a_5441_16911 VGND 0.23f
C1259 a_7571_16911 VGND 0.524f
C1260 a_7159_17076 VGND 0.524f
C1261 tdc0.w_ring_norsz28 VGND 2.38f
C1262 a_5951_17277 VGND 0.609f
C1263 a_6119_17179 VGND 0.817f
C1264 a_5526_17277 VGND 0.626f
C1265 a_5694_17023 VGND 0.581f
C1266 a_5253_16911 VGND 1.43f
C1267 a_5087_16911 VGND 1.81f
C1268 tdc0.w_ring_buf17 VGND 0.872f
C1269 a_3601_16911 VGND 0.23f
C1270 a_4811_16911 VGND 0.524f
C1271 a_4111_17277 VGND 0.609f
C1272 a_4279_17179 VGND 0.817f
C1273 a_3686_17277 VGND 0.626f
C1274 a_3854_17023 VGND 0.581f
C1275 a_3413_16911 VGND 1.43f
C1276 a_3247_16911 VGND 1.81f
C1277 tdc0.r_ring_ctr15 VGND 2.31f
C1278 a_1847_17277 VGND 0.168f
C1279 a_1644_16911 VGND 0.259f
C1280 a_2304_16911 VGND 0.736f
C1281 a_2479_16885 VGND 0.971f
C1282 a_1739_16911 VGND 0.714f
C1283 _047_ VGND 1.66f
C1284 a_1957_17153 VGND 0.653f
C1285 a_1389_16911 VGND 1.57f
C1286 _006_ VGND 1.26f
C1287 a_1223_16911 VGND 1.92f
C1288 tdc1.r_dly_store_ring30 VGND 6.13f
C1289 a_30005_17455 VGND 0.23f
C1290 a_30515_17455 VGND 0.609f
C1291 a_30683_17429 VGND 0.817f
C1292 a_30090_17455 VGND 0.626f
C1293 a_30258_17429 VGND 0.581f
C1294 a_29817_17461 VGND 1.43f
C1295 a_29651_17461 VGND 1.81f
C1296 net76 VGND 1.09f
C1297 tdc1.w_ring_norsz28 VGND 2.48f
C1298 tdc1.w_ring_norsz12 VGND 2.6f
C1299 a_27815_17429 VGND 0.74f
C1300 a_27705_17687 VGND 0.768f
C1301 tdc1.r_dly_store_ctr5 VGND 1.98f
C1302 a_27346_17687 VGND 0.711f
C1303 a_26895_17429 VGND 0.74f
C1304 a_26785_17687 VGND 0.768f
C1305 tdc1.r_dly_store_ring11 VGND 1.29f
C1306 _104_ VGND 2.42f
C1307 a_26426_17687 VGND 0.711f
C1308 a_25551_17545 VGND 0.478f
C1309 _086_ VGND 4.89f
C1310 _081_ VGND 1.85f
C1311 a_23289_17455 VGND 0.23f
C1312 tdc1.w_ring_buf3 VGND 1.37f
C1313 a_25381_17429 VGND 0.485f
C1314 a_24819_17776 VGND 0.641f
C1315 tdc1.r_dly_store_ring25 VGND 0.836f
C1316 a_24455_17687 VGND 0.673f
C1317 a_23799_17455 VGND 0.609f
C1318 a_23967_17429 VGND 0.817f
C1319 a_23374_17455 VGND 0.626f
C1320 a_23542_17429 VGND 0.581f
C1321 a_23101_17461 VGND 1.43f
C1322 a_22935_17461 VGND 1.81f
C1323 a_20911_17455 VGND 0.524f
C1324 tdc1.g_ring320.stg01_67.HI VGND 0.415f
C1325 tdc1.r_dly_store_ring22 VGND 1.31f
C1326 a_17309_17455 VGND 0.23f
C1327 tdc1.w_ring_buf4 VGND 1.2f
C1328 a_12897_17455 VGND 0.206f
C1329 _117_ VGND 0.952f
C1330 _116_ VGND 1.16f
C1331 net67 VGND 1f
C1332 tdc1.w_ring_int_norsz4 VGND 0.839f
C1333 tdc1.w_ring_int_norsz20 VGND 0.878f
C1334 tdc1.w_ring_norsz20 VGND 2.44f
C1335 a_17819_17455 VGND 0.609f
C1336 a_17987_17429 VGND 0.817f
C1337 a_17394_17455 VGND 0.626f
C1338 a_17562_17429 VGND 0.581f
C1339 a_17121_17461 VGND 1.43f
C1340 a_16955_17461 VGND 1.81f
C1341 a_15715_17674 VGND 0.524f
C1342 a_14857_17753 VGND 0.607f
C1343 tdc1.r_dly_store_ring4 VGND 1.22f
C1344 a_14428_17687 VGND 0.59f
C1345 a_13461_17571 VGND 0.665f
C1346 _113_ VGND 1.26f
C1347 _114_ VGND 0.941f
C1348 a_12815_17455 VGND 0.804f
C1349 net25 VGND 9.42f
C1350 tdc0.r_dly_store_ctr7 VGND 4.61f
C1351 _071_ VGND 10.3f
C1352 tdc0.r_dly_store_ctr15 VGND 4.49f
C1353 tdc0.w_ring_int_norsz2 VGND 0.722f
C1354 tdc0.w_ring_norsz18 VGND 2.37f
C1355 a_9839_17715 VGND 1.2f
C1356 tdc0.w_ring_norsz3 VGND 2.36f
C1357 tdc0.w_ring_norsz19 VGND 3.13f
C1358 net49 VGND 0.822f
C1359 tdc0.g_ring320.stg01_49.HI VGND 0.415f
C1360 net58 VGND 1.13f
C1361 a_7833_17455 VGND 0.23f
C1362 a_8343_17455 VGND 0.609f
C1363 a_8511_17429 VGND 0.817f
C1364 a_7918_17455 VGND 0.626f
C1365 a_8086_17429 VGND 0.581f
C1366 a_7645_17461 VGND 1.43f
C1367 a_7479_17461 VGND 1.81f
C1368 tdc0.w_ring_int_norsz29 VGND 0.923f
C1369 tdc0.g_ring329.stg01_58.HI VGND 0.415f
C1370 tdc0.w_ring_int_norsz13 VGND 0.995f
C1371 tdc0.w_ring_int_norsz18 VGND 2.6f
C1372 net7 VGND 11f
C1373 tdc0.w_ring_int_norsz17 VGND 0.987f
C1374 tdc0.w_ring_norsz17 VGND 2.31f
C1375 a_4585_17674 VGND 0.524f
C1376 tdc0.w_ring_buf0 VGND 6.61f
C1377 a_1368_17429 VGND 0.648f
C1378 a_29913_17999 VGND 0.23f
C1379 a_30423_18365 VGND 0.609f
C1380 a_30591_18267 VGND 0.817f
C1381 a_29998_18365 VGND 0.626f
C1382 a_30166_18111 VGND 0.581f
C1383 a_29725_17999 VGND 1.43f
C1384 a_29559_17999 VGND 1.81f
C1385 a_27012_18249 VGND 0.259f
C1386 a_24385_18249 VGND 0.393f
C1387 a_24131_18249 VGND 0.388f
C1388 tdc1.w_ring_buf25 VGND 0.922f
C1389 tdc1.g_ring325.stg01_72.HI VGND 0.415f
C1390 _125_ VGND 1.52f
C1391 _124_ VGND 3.18f
C1392 tdc1.w_ring_int_norsz13 VGND 0.897f
C1393 tdc1.w_ring_int_norsz29 VGND 1.18f
C1394 a_27403_17973 VGND 0.698f
C1395 tdc1.r_dly_store_ring13 VGND 2.29f
C1396 _123_ VGND 1.1f
C1397 a_26581_18145 VGND 0.672f
C1398 a_25971_17999 VGND 0.698f
C1399 a_24635_17973 VGND 0.587f
C1400 a_23259_18164 VGND 0.524f
C1401 tdc1.w_ring_int_norsz26 VGND 0.878f
C1402 tdc1.w_ring_norsz26 VGND 4.55f
C1403 tdc1.w_ring_int_norsz10 VGND 1.27f
C1404 a_20316_18151 VGND 0.665f
C1405 tdc1.w_ring_norsz4 VGND 3.51f
C1406 tdc1.w_ring_int_norsz5 VGND 0.722f
C1407 tdc1.w_ring_int_norsz21 VGND 0.897f
C1408 a_18243_17999 VGND 0.648f
C1409 tdc0.r_dly_store_ring4 VGND 1.02f
C1410 a_13905_17999 VGND 0.23f
C1411 a_14415_18365 VGND 0.609f
C1412 a_14583_18267 VGND 0.817f
C1413 a_13990_18365 VGND 0.626f
C1414 a_14158_18111 VGND 0.581f
C1415 a_13717_17999 VGND 1.43f
C1416 a_13551_17999 VGND 1.81f
C1417 tdc0.w_ring_buf4 VGND 1.26f
C1418 a_11237_17999 VGND 0.23f
C1419 a_12355_17999 VGND 0.524f
C1420 a_11747_18365 VGND 0.609f
C1421 a_11915_18267 VGND 0.817f
C1422 a_11322_18365 VGND 0.626f
C1423 a_11490_18111 VGND 0.581f
C1424 a_11049_17999 VGND 1.43f
C1425 a_10883_17999 VGND 1.81f
C1426 tdc0.w_ring_int_norsz3 VGND 1.36f
C1427 tdc0.w_ring_buf12 VGND 0.967f
C1428 tdc0.w_ring_int_norsz20 VGND 1.29f
C1429 tdc0.w_ring_int_norsz4 VGND 0.936f
C1430 a_7479_17999 VGND 0.524f
C1431 tdc0.w_ring_norsz12 VGND 3.01f
C1432 a_7111_17999 VGND 0.698f
C1433 net23 VGND 6.2f
C1434 a_6796_17973 VGND 0.648f
C1435 tdc0.w_ring_norsz29 VGND 2.72f
C1436 net59 VGND 0.822f
C1437 tdc0.g_ring330.stg01_59.HI VGND 0.415f
C1438 a_5455_17999 VGND 0.524f
C1439 tdc0.w_ring_norsz1 VGND 1.65f
C1440 net47 VGND 1.38f
C1441 tdc0.g_ring318.stg01_47.HI VGND 0.415f
C1442 tdc0.w_ring_int_norsz1 VGND 1.55f
C1443 net46 VGND 1.12f
C1444 tdc0.g_ring317.stg01_46.HI VGND 0.415f
C1445 a_30725_18921 VGND 0.23f
C1446 tdc1.w_ring_buf13 VGND 1.08f
C1447 _122_ VGND 1.37f
C1448 _121_ VGND 0.922f
C1449 a_30307_18921 VGND 0.581f
C1450 a_30378_18820 VGND 0.626f
C1451 a_30178_18665 VGND 1.43f
C1452 a_30171_18761 VGND 1.81f
C1453 a_29887_18775 VGND 0.609f
C1454 a_29791_18775 VGND 0.817f
C1455 a_29375_18543 VGND 0.524f
C1456 tdc1.w_ring_norsz13 VGND 2.05f
C1457 a_27517_18543 VGND 0.673f
C1458 tdc1.r_dly_store_ring29 VGND 1.54f
C1459 a_27351_18543 VGND 0.641f
C1460 a_26747_18863 VGND 0.711f
C1461 a_26627_18543 VGND 0.768f
C1462 a_26431_18543 VGND 0.74f
C1463 a_25971_18551 VGND 0.648f
C1464 a_25643_18775 VGND 0.454f
C1465 _129_ VGND 6.61f
C1466 a_25287_18517 VGND 0.753f
C1467 a_24451_18864 VGND 0.641f
C1468 a_24087_18775 VGND 0.673f
C1469 tdc1.w_ring_norsz10 VGND 4.34f
C1470 a_23075_18762 VGND 0.524f
C1471 tdc1.g_ring326.stg01_73.HI VGND 0.415f
C1472 net73 VGND 1.24f
C1473 tdc1.r_dly_store_ring21 VGND 2.59f
C1474 a_21633_18543 VGND 0.23f
C1475 net68 VGND 1.23f
C1476 a_22143_18543 VGND 0.609f
C1477 a_22311_18517 VGND 0.817f
C1478 a_21718_18543 VGND 0.626f
C1479 a_21886_18517 VGND 0.581f
C1480 a_21445_18549 VGND 1.43f
C1481 tdc1.w_ring_buf21 VGND 1.69f
C1482 a_21279_18549 VGND 1.81f
C1483 tdc1.w_ring_norsz25 VGND 3.4f
C1484 tdc1.w_ring_int_norsz25 VGND 0.878f
C1485 a_19899_18543 VGND 0.698f
C1486 net16 VGND 13.4f
C1487 net72 VGND 1.2f
C1488 a_19071_18543 VGND 0.524f
C1489 tdc1.g_ring321.stg01_68.HI VGND 0.415f
C1490 tdc1.w_ring_buf22 VGND 1.28f
C1491 tdc0.r_dly_store_ring30 VGND 3.8f
C1492 a_13625_18543 VGND 0.214f
C1493 a_13541_18543 VGND 0.167f
C1494 a_12889_18543 VGND 0.214f
C1495 a_12805_18543 VGND 0.167f
C1496 a_16481_18543 VGND 0.23f
C1497 a_14195_18863 VGND 0.146f
C1498 _115_ VGND 1.06f
C1499 tdc0.w_ring_buf20 VGND 1.24f
C1500 tdc1.w_ring_norsz21 VGND 1.98f
C1501 tdc1.w_ring_norsz5 VGND 3.11f
C1502 a_17647_18762 VGND 0.524f
C1503 a_16991_18543 VGND 0.609f
C1504 a_17159_18517 VGND 0.817f
C1505 a_16566_18543 VGND 0.626f
C1506 a_16734_18517 VGND 0.581f
C1507 a_16293_18549 VGND 1.43f
C1508 a_16127_18549 VGND 1.81f
C1509 a_14372_18543 VGND 0.724f
C1510 _126_ VGND 3.59f
C1511 _120_ VGND 0.678f
C1512 _119_ VGND 2.01f
C1513 a_13459_18543 VGND 0.972f
C1514 a_12723_18543 VGND 0.972f
C1515 tdc0.r_dly_store_ring20 VGND 1.18f
C1516 tdc0.r_dly_store_ring12 VGND 2.8f
C1517 a_11067_18543 VGND 0.524f
C1518 tdc0.w_ring_norsz2 VGND 2.51f
C1519 a_10331_18543 VGND 0.524f
C1520 tdc0.w_ring_norsz4 VGND 2.85f
C1521 tdc0.w_ring_int_norsz5 VGND 0.967f
C1522 tdc0.g_ring321.stg01_50.HI VGND 0.415f
C1523 tdc0.w_ring_buf21 VGND 1.87f
C1524 tdc0.r_dly_store_ring13 VGND 3.13f
C1525 a_7465_18543 VGND 0.23f
C1526 tdc0.w_ring_norsz0 VGND 2.25f
C1527 a_8767_18543 VGND 0.524f
C1528 a_7975_18543 VGND 0.609f
C1529 a_8143_18517 VGND 0.817f
C1530 a_7550_18543 VGND 0.626f
C1531 a_7718_18517 VGND 0.581f
C1532 a_7277_18549 VGND 1.43f
C1533 a_7111_18549 VGND 1.81f
C1534 tdc0.w_ring_int_norsz14 VGND 1.03f
C1535 tdc0.w_ring_int_norsz30 VGND 1.06f
C1536 tdc0.w_ring_norsz16 VGND 4.63f
C1537 tdc0.w_ring_int_norsz0 VGND 1.17f
C1538 a_4443_18543 VGND 1.2f
C1539 net44 VGND 1.03f
C1540 tdc0.g_ring116.stg02_44.HI VGND 0.415f
C1541 _626_.X VGND 0.226f
C1542 a_2656_18517 VGND 0.648f
C1543 tdc1.g_ring330.stg01_77.HI VGND 0.415f
C1544 tdc1.w_ring_buf29 VGND 1.08f
C1545 a_30295_19087 VGND 0.524f
C1546 tdc1.w_ring_norsz29 VGND 3.24f
C1547 net77 VGND 1.62f
C1548 tdc1.w_ring_buf30 VGND 1.35f
C1549 a_29743_19087 VGND 0.524f
C1550 tdc1.w_ring_int_norsz30 VGND 1.12f
C1551 tdc1.w_ring_int_norsz14 VGND 0.897f
C1552 a_27259_19087 VGND 0.648f
C1553 _074_ VGND 1.63f
C1554 _066_ VGND 2.41f
C1555 a_24213_19337 VGND 0.206f
C1556 a_22645_19087 VGND 0.23f
C1557 a_26754_19133 VGND 0.611f
C1558 _067_ VGND 8.41f
C1559 a_24822_19133 VGND 0.611f
C1560 _065_ VGND 9.39f
C1561 _064_ VGND 8.4f
C1562 a_24131_19337 VGND 0.804f
C1563 a_23155_19453 VGND 0.609f
C1564 a_23323_19355 VGND 0.817f
C1565 a_22730_19453 VGND 0.626f
C1566 a_22898_19199 VGND 0.581f
C1567 a_22457_19087 VGND 1.43f
C1568 tdc1.w_ring_buf10 VGND 1.11f
C1569 a_22291_19087 VGND 1.81f
C1570 tdc1.g_ring322.stg01_69.HI VGND 0.415f
C1571 tdc1.w_ring_int_norsz9 VGND 1.38f
C1572 a_21923_19087 VGND 0.524f
C1573 a_20727_19087 VGND 0.524f
C1574 tdc1.w_ring_norsz9 VGND 2.33f
C1575 tdc1.w_ring_int_norsz24 VGND 0.867f
C1576 tdc1.w_ring_norsz8 VGND 3.73f
C1577 tdc1.w_ring_norsz24 VGND 4.49f
C1578 tdc1.w_ring_int_norsz8 VGND 0.722f
C1579 net69 VGND 1.2f
C1580 _100_ VGND 1.9f
C1581 a_15801_19414 VGND 0.607f
C1582 tdc0.r_dly_store_ring2 VGND 0.948f
C1583 a_14641_19087 VGND 0.23f
C1584 tdc1.w_ring_int_norsz22 VGND 0.936f
C1585 tdc1.w_ring_int_norsz6 VGND 0.975f
C1586 tdc1.w_ring_norsz22 VGND 2.07f
C1587 a_16055_19414 VGND 0.59f
C1588 a_15151_19453 VGND 0.609f
C1589 a_15319_19355 VGND 0.817f
C1590 a_14726_19453 VGND 0.626f
C1591 a_14894_19199 VGND 0.581f
C1592 a_14453_19087 VGND 1.43f
C1593 tdc0.w_ring_buf2 VGND 2.31f
C1594 a_14287_19087 VGND 1.81f
C1595 tdc0.r_dly_store_ring5 VGND 1.08f
C1596 a_11789_19087 VGND 0.23f
C1597 a_13583_19115 VGND 0.56f
C1598 a_12299_19453 VGND 0.609f
C1599 a_12467_19355 VGND 0.817f
C1600 a_11874_19453 VGND 0.626f
C1601 a_12042_19199 VGND 0.581f
C1602 a_11601_19087 VGND 1.43f
C1603 a_11435_19087 VGND 1.81f
C1604 tdc0.w_ring_buf5 VGND 1.22f
C1605 tdc0.w_ring_int_norsz21 VGND 0.931f
C1606 tdc0.w_ring_buf13 VGND 1.02f
C1607 tdc0.w_ring_buf30 VGND 5.13f
C1608 tdc0.w_ring_int_norsz31 VGND 1.33f
C1609 tdc0.stg01_61.HI VGND 0.415f
C1610 a_5257_19087 VGND 0.23f
C1611 tdc0.w_ring_int_norsz24 VGND 0.975f
C1612 tdc0.w_ring_norsz24 VGND 4.53f
C1613 a_10331_19087 VGND 0.524f
C1614 tdc0.w_ring_int_norsz7 VGND 1.35f
C1615 tdc0.w_ring_norsz20 VGND 2.4f
C1616 net50 VGND 1.4f
C1617 tdc0.w_ring_norsz5 VGND 2.72f
C1618 tdc0.w_ring_norsz21 VGND 2.45f
C1619 a_6927_19087 VGND 0.524f
C1620 tdc0.w_ring_norsz13 VGND 3.1f
C1621 a_6651_19087 VGND 0.524f
C1622 tdc0.w_ring_norsz30 VGND 1.91f
C1623 a_5767_19453 VGND 0.609f
C1624 a_5935_19355 VGND 0.817f
C1625 a_5342_19453 VGND 0.626f
C1626 a_5510_19199 VGND 0.581f
C1627 a_5069_19087 VGND 1.43f
C1628 a_4903_19087 VGND 1.81f
C1629 net20 VGND 10.4f
C1630 a_4404_19061 VGND 0.648f
C1631 net61 VGND 1.47f
C1632 a_3571_19252 VGND 0.524f
C1633 a_3295_19252 VGND 0.524f
C1634 a_29743_19631 VGND 0.524f
C1635 tdc1.g_ring331.stg01_78.HI VGND 0.415f
C1636 a_27689_20009 VGND 0.23f
C1637 a_25441_19631 VGND 0.324f
C1638 a_24397_19631 VGND 0.206f
C1639 tdc1.r_dly_store_ring31 VGND 1.85f
C1640 a_25892_19951 VGND 0.28f
C1641 a_25251_19951 VGND 0.337f
C1642 _087_ VGND 6f
C1643 _097_ VGND 2.05f
C1644 tdc1.r_dly_store_ring23 VGND 0.792f
C1645 a_23105_19631 VGND 0.23f
C1646 net71 VGND 1.33f
C1647 a_21633_19631 VGND 0.23f
C1648 a_29099_19631 VGND 0.698f
C1649 tdc1.w_ring_norsz30 VGND 2.17f
C1650 net78 VGND 1.17f
C1651 tdc1.w_ring_norsz14 VGND 2.66f
C1652 a_27271_20009 VGND 0.581f
C1653 a_27342_19908 VGND 0.626f
C1654 a_27142_19753 VGND 1.43f
C1655 a_27135_19849 VGND 1.81f
C1656 a_26851_19863 VGND 0.609f
C1657 a_26755_19863 VGND 0.817f
C1658 a_25221_19605 VGND 1.14f
C1659 tdc1.r_dly_store_ring10 VGND 1.28f
C1660 a_24251_19863 VGND 0.804f
C1661 a_23615_19631 VGND 0.609f
C1662 a_23783_19605 VGND 0.817f
C1663 a_23190_19631 VGND 0.626f
C1664 a_23358_19605 VGND 0.581f
C1665 a_22917_19637 VGND 1.43f
C1666 tdc1.w_ring_buf23 VGND 1.35f
C1667 a_22751_19637 VGND 1.81f
C1668 a_22143_19631 VGND 0.609f
C1669 a_22311_19605 VGND 0.817f
C1670 a_21718_19631 VGND 0.626f
C1671 a_21886_19605 VGND 0.581f
C1672 a_21445_19637 VGND 1.43f
C1673 tdc1.w_ring_buf9 VGND 1.23f
C1674 a_21279_19637 VGND 1.81f
C1675 tdc1.w_ring_norsz3 VGND 2.86f
C1676 tdc1.w_ring_norsz19 VGND 3.33f
C1677 tdc1.g_ring324.stg01_71.HI VGND 0.415f
C1678 a_18045_19631 VGND 0.23f
C1679 tdc1.r_dly_store_ring2 VGND 1.15f
C1680 a_13349_19631 VGND 0.214f
C1681 a_13265_19631 VGND 0.167f
C1682 a_14917_19631 VGND 0.23f
C1683 a_19211_19850 VGND 0.524f
C1684 a_18555_19631 VGND 0.609f
C1685 a_18723_19605 VGND 0.817f
C1686 a_18130_19631 VGND 0.626f
C1687 a_18298_19605 VGND 0.581f
C1688 a_17857_19637 VGND 1.43f
C1689 tdc1.w_ring_buf6 VGND 1.53f
C1690 a_17691_19637 VGND 1.81f
C1691 tdc1.w_ring_int_norsz23 VGND 0.878f
C1692 net14 VGND 6.12f
C1693 tdc1.w_ring_norsz23 VGND 4.05f
C1694 a_16679_19631 VGND 0.524f
C1695 tdc1.w_ring_norsz7 VGND 2.99f
C1696 _072_ VGND 9.87f
C1697 a_16187_19891 VGND 1.2f
C1698 a_15427_19631 VGND 0.609f
C1699 a_15595_19605 VGND 0.817f
C1700 a_15002_19631 VGND 0.626f
C1701 a_15170_19605 VGND 0.581f
C1702 a_14729_19637 VGND 1.43f
C1703 a_14563_19637 VGND 1.81f
C1704 a_13921_19747 VGND 0.665f
C1705 _135_ VGND 0.933f
C1706 _136_ VGND 1.85f
C1707 _137_ VGND 0.655f
C1708 tdc0.r_dly_store_ring23 VGND 1.27f
C1709 a_11697_19631 VGND 0.23f
C1710 net51 VGND 1.27f
C1711 a_13183_19631 VGND 0.972f
C1712 _068_ VGND 9.91f
C1713 tdc0.r_dly_store_ring15 VGND 4.09f
C1714 a_12207_19631 VGND 0.609f
C1715 a_12375_19605 VGND 0.817f
C1716 a_11782_19631 VGND 0.626f
C1717 a_11950_19605 VGND 0.581f
C1718 a_11509_19637 VGND 1.43f
C1719 tdc0.w_ring_buf23 VGND 0.872f
C1720 a_11343_19637 VGND 1.81f
C1721 a_11067_19631 VGND 0.524f
C1722 tdc0.w_ring_norsz23 VGND 2.94f
C1723 a_9963_19631 VGND 0.698f
C1724 tdc0.w_ring_int_norsz6 VGND 0.923f
C1725 tdc0.w_ring_int_norsz22 VGND 1f
C1726 tdc0.g_ring322.stg01_51.HI VGND 0.415f
C1727 tdc0.r_dly_store_ring31 VGND 3.23f
C1728 net60 VGND 1.17f
C1729 a_6913_19631 VGND 0.23f
C1730 a_7423_19631 VGND 0.609f
C1731 a_7591_19605 VGND 0.817f
C1732 a_6998_19631 VGND 0.626f
C1733 a_7166_19605 VGND 0.581f
C1734 a_6725_19637 VGND 1.43f
C1735 a_6559_19637 VGND 1.81f
C1736 a_6283_19631 VGND 0.524f
C1737 tdc0.w_ring_norsz14 VGND 2.76f
C1738 tdc0.g_ring331.stg01_60.HI VGND 0.415f
C1739 tdc0.w_ring_int_norsz16 VGND 2.65f
C1740 tdc0.w_ring_int_norsz15 VGND 1.63f
C1741 net19 VGND 8.08f
C1742 a_5087_19631 VGND 0.524f
C1743 net39 VGND 12f
C1744 net13 VGND 2.76f
C1745 tdc0.g_ring316.stg01_45.HI VGND 0.415f
C1746 net45 VGND 1.35f
C1747 tdc0.w_dly_stop5 VGND 3.22f
C1748 tdc0.w_dly_stop2 VGND 1.09f
C1749 a_3707_19631 VGND 0.524f
C1750 tdc0.w_dly_stop4 VGND 0.762f
C1751 a_3247_19631 VGND 0.524f
C1752 tdc0.w_dly_stop3 VGND 0.975f
C1753 a_2971_19631 VGND 0.524f
C1754 tdc0.w_dly_stop1 VGND 0.968f
C1755 a_29989_20175 VGND 0.23f
C1756 tdc1.w_ring_buf14 VGND 0.994f
C1757 a_29571_20175 VGND 0.581f
C1758 a_29642_20149 VGND 0.626f
C1759 a_29435_20149 VGND 1.81f
C1760 a_29442_20449 VGND 1.43f
C1761 a_29151_20149 VGND 0.609f
C1762 a_29055_20327 VGND 0.817f
C1763 tdc1.w_ring_int_norsz15 VGND 1.09f
C1764 tdc1.w_ring_int_norsz31 VGND 1.01f
C1765 tdc1.stg01_79.HI VGND 0.415f
C1766 tdc1.w_ring_buf31 VGND 1.19f
C1767 tdc1.w_ring_buf0 VGND 4.23f
C1768 a_22160_20175 VGND 0.205f
C1769 a_18030_20175 VGND 0.161f
C1770 a_17678_20175 VGND 0.123f
C1771 _141_ VGND 2.83f
C1772 _140_ VGND 1.18f
C1773 _139_ VGND 0.802f
C1774 a_22855_20425 VGND 0.167f
C1775 a_22653_20425 VGND 0.214f
C1776 tdc1.w_ring_int_norsz3 VGND 0.902f
C1777 tdc1.w_ring_buf2 VGND 3.3f
C1778 a_19267_20425 VGND 0.167f
C1779 a_19065_20425 VGND 0.214f
C1780 a_17596_20425 VGND 0.537f
C1781 a_14994_20175 VGND 0.161f
C1782 a_14642_20175 VGND 0.123f
C1783 a_16353_20502 VGND 0.607f
C1784 a_14560_20425 VGND 0.537f
C1785 tdc0.g_ring324.stg01_53.HI VGND 0.415f
C1786 a_26983_20175 VGND 0.524f
C1787 a_26297_20340 VGND 0.524f
C1788 a_25111_20327 VGND 0.56f
C1789 a_24546_20327 VGND 0.702f
C1790 tdc1.r_dly_store_ring9 VGND 0.899f
C1791 _083_ VGND 16.4f
C1792 a_22527_20327 VGND 0.972f
C1793 _082_ VGND 2.3f
C1794 _085_ VGND 0.7f
C1795 a_21934_20221 VGND 0.443f
C1796 a_21791_20327 VGND 0.65f
C1797 a_20131_20340 VGND 0.524f
C1798 _084_ VGND 12.3f
C1799 tdc1.r_dly_store_ring6 VGND 0.899f
C1800 tdc1.r_dly_store_ring14 VGND 5.29f
C1801 _075_ VGND 16.2f
C1802 a_18939_20327 VGND 0.972f
C1803 _078_ VGND 3.05f
C1804 _090_ VGND 2.39f
C1805 _091_ VGND 1.05f
C1806 a_17208_20149 VGND 1.37f
C1807 a_16607_20502 VGND 0.59f
C1808 net24 VGND 10.4f
C1809 a_15451_20149 VGND 1.2f
C1810 _138_ VGND 1.24f
C1811 _142_ VGND 5.08f
C1812 a_14172_20149 VGND 1.37f
C1813 a_13611_20327 VGND 0.56f
C1814 a_12875_20327 VGND 0.56f
C1815 net53 VGND 1.95f
C1816 net11 VGND 5.4f
C1817 tdc0.r_dly_store_ring22 VGND 1.48f
C1818 a_10317_20175 VGND 0.23f
C1819 a_11435_20175 VGND 0.524f
C1820 tdc0.w_ring_norsz8 VGND 1.98f
C1821 a_10827_20541 VGND 0.609f
C1822 a_10995_20443 VGND 0.817f
C1823 a_10402_20541 VGND 0.626f
C1824 a_10570_20287 VGND 0.581f
C1825 a_10129_20175 VGND 1.43f
C1826 a_9963_20175 VGND 1.81f
C1827 tdc0.w_ring_int_norsz23 VGND 0.941f
C1828 net52 VGND 0.822f
C1829 tdc0.g_ring323.stg01_52.HI VGND 0.415f
C1830 net22 VGND 7.3f
C1831 net21 VGND 6.23f
C1832 tdc0.r_dly_store_ring14 VGND 3.15f
C1833 a_7097_20175 VGND 0.23f
C1834 a_9004_20149 VGND 0.648f
C1835 a_8675_20175 VGND 0.524f
C1836 tdc0.w_ring_norsz6 VGND 2.21f
C1837 a_7607_20541 VGND 0.609f
C1838 a_7775_20443 VGND 0.817f
C1839 a_7182_20541 VGND 0.626f
C1840 a_7350_20287 VGND 0.581f
C1841 a_6909_20175 VGND 1.43f
C1842 tdc0.w_ring_buf14 VGND 1.13f
C1843 a_6743_20175 VGND 1.81f
C1844 tdc0.w_ring_buf31 VGND 1.18f
C1845 tdc0.w_ring_buf15 VGND 1.23f
C1846 a_6007_20175 VGND 0.524f
C1847 tdc0.w_ring_norsz31 VGND 3.22f
C1848 a_4903_20175 VGND 0.524f
C1849 tdc0.w_ring_norsz15 VGND 1.7f
C1850 a_28885_21097 VGND 0.23f
C1851 tdc1.r_dly_store_ring15 VGND 2.14f
C1852 tdc1.w_ring_buf16 VGND 3.09f
C1853 tdc1.r_dly_store_ring18 VGND 1.04f
C1854 a_23381_20719 VGND 0.23f
C1855 tdc1.w_ring_int_norsz19 VGND 1.59f
C1856 tdc1.w_ring_norsz15 VGND 3.59f
C1857 a_29791_20938 VGND 0.524f
C1858 a_29427_20693 VGND 0.698f
C1859 net37 VGND 8.27f
C1860 tdc1.w_ring_buf15 VGND 1.06f
C1861 a_28467_21097 VGND 0.581f
C1862 a_28538_20996 VGND 0.626f
C1863 a_28338_20841 VGND 1.43f
C1864 a_28331_20937 VGND 1.81f
C1865 a_28047_20951 VGND 0.609f
C1866 a_27951_20951 VGND 0.817f
C1867 tdc1.w_ring_norsz31 VGND 2.72f
C1868 net79 VGND 1.09f
C1869 net17 VGND 8.09f
C1870 tdc1.w_ring_int_norsz16 VGND 2.21f
C1871 tdc1.w_ring_int_norsz0 VGND 1.03f
C1872 a_26111_20938 VGND 0.524f
C1873 a_25787_20719 VGND 0.524f
C1874 tdc1.w_ring_norsz0 VGND 2.38f
C1875 tdc1.w_ring_norsz16 VGND 3.18f
C1876 tdc1.w_ring_int_norsz1 VGND 0.917f
C1877 a_23891_20719 VGND 0.609f
C1878 a_24059_20693 VGND 0.817f
C1879 a_23466_20719 VGND 0.626f
C1880 a_23634_20693 VGND 0.581f
C1881 a_23193_20725 VGND 1.43f
C1882 tdc1.w_ring_buf18 VGND 1.34f
C1883 a_23027_20725 VGND 1.81f
C1884 a_22247_20938 VGND 0.524f
C1885 a_21647_20719 VGND 0.524f
C1886 tdc1.w_ring_int_norsz18 VGND 0.839f
C1887 tdc1.w_ring_norsz2 VGND 2.26f
C1888 net66 VGND 1.01f
C1889 tdc1.w_ring_int_norsz2 VGND 0.923f
C1890 tdc1.w_ring_norsz18 VGND 1.97f
C1891 net15 VGND 6.23f
C1892 tdc1.g_ring319.stg01_66.HI VGND 0.415f
C1893 tdc1.w_ring_int_norsz7 VGND 1.72f
C1894 a_18887_20719 VGND 0.524f
C1895 tdc1.w_ring_norsz6 VGND 3.17f
C1896 net41 VGND 11f
C1897 tdc1.g_ring323.stg01_70.HI VGND 0.415f
C1898 net70 VGND 1.82f
C1899 a_17661_21097 VGND 0.23f
C1900 tdc0.r_dly_store_ring1 VGND 1.34f
C1901 a_14166_20719 VGND 0.171f
C1902 a_13814_20719 VGND 0.14f
C1903 a_12448_20719 VGND 0.259f
C1904 a_14917_20719 VGND 0.23f
C1905 a_13732_21039 VGND 0.482f
C1906 tdc1.w_ring_buf7 VGND 1.57f
C1907 a_17243_21097 VGND 0.581f
C1908 a_17314_20996 VGND 0.626f
C1909 a_17114_20841 VGND 1.43f
C1910 a_17107_20937 VGND 1.81f
C1911 a_16823_20951 VGND 0.609f
C1912 a_16727_20951 VGND 0.817f
C1913 net12 VGND 7.35f
C1914 a_16175_20938 VGND 0.524f
C1915 a_15427_20719 VGND 0.609f
C1916 a_15595_20693 VGND 0.817f
C1917 a_15002_20719 VGND 0.626f
C1918 a_15170_20693 VGND 0.581f
C1919 a_14729_20725 VGND 1.43f
C1920 tdc0.w_ring_buf1 VGND 1.28f
C1921 a_14563_20725 VGND 1.81f
C1922 _131_ VGND 1.16f
C1923 _134_ VGND 6f
C1924 _132_ VGND 3.35f
C1925 a_13344_20693 VGND 1.37f
C1926 a_12618_21039 VGND 0.672f
C1927 _130_ VGND 2.9f
C1928 _128_ VGND 0.844f
C1929 _127_ VGND 1.28f
C1930 _089_ VGND 16.5f
C1931 tt_um_hpretl_tt06_tdc_v2_88.HI VGND 0.415f
C1932 tdc0.w_ring_int_norsz8 VGND 1.4f
C1933 tdc0.w_ring_buf22 VGND 0.975f
C1934 tdc0.r_dly_store_ring6 VGND 1.71f
C1935 a_9121_20719 VGND 0.23f
C1936 a_11251_20719 VGND 0.524f
C1937 tdc0.w_ring_norsz7 VGND 2.95f
C1938 net40 VGND 6.52f
C1939 tdc0.w_ring_norsz22 VGND 2.75f
C1940 a_10287_20938 VGND 0.524f
C1941 a_9631_20719 VGND 0.609f
C1942 a_9799_20693 VGND 0.817f
C1943 a_9206_20719 VGND 0.626f
C1944 a_9374_20693 VGND 0.581f
C1945 a_8933_20725 VGND 1.43f
C1946 tdc0.w_ring_buf6 VGND 1.03f
C1947 a_8767_20725 VGND 1.81f
C1948 tdc1.g_ring316.stg01_63.HI VGND 0.415f
C1949 net2 VGND 0.876f
C1950 a_29883_21428 VGND 0.524f
C1951 a_29559_21263 VGND 0.524f
C1952 net63 VGND 2.36f
C1953 net4 VGND 4.19f
C1954 net42 VGND 7.16f
C1955 net5 VGND 5.01f
C1956 net6 VGND 3.73f
C1957 a_29057_21428 VGND 0.524f
C1958 a_28415_21237 VGND 0.698f
C1959 net1 VGND 1.31f
C1960 a_28047_21237 VGND 0.698f
C1961 net43 VGND 13.3f
C1962 a_27679_21237 VGND 0.698f
C1963 a_26667_21237 VGND 0.698f
C1964 a_25879_21263 VGND 0.524f
C1965 net62 VGND 1.75f
C1966 tdc1.g_ring116.stg02_62.HI VGND 0.415f
C1967 tdc1.g_ring317.stg01_64.HI VGND 0.415f
C1968 net64 VGND 1.12f
C1969 tdc1.w_ring_norsz17 VGND 2.89f
C1970 tdc1.w_ring_int_norsz17 VGND 1.09f
C1971 tdc1.w_ring_norsz1 VGND 4.92f
C1972 net18 VGND 7.19f
C1973 a_23907_21237 VGND 0.698f
C1974 net35 VGND 11.9f
C1975 tdc1.r_dly_store_ring17 VGND 1.2f
C1976 a_22093_21263 VGND 0.23f
C1977 a_23264_21237 VGND 0.648f
C1978 a_22603_21629 VGND 0.609f
C1979 a_22771_21531 VGND 0.817f
C1980 a_22178_21629 VGND 0.626f
C1981 a_22346_21375 VGND 0.581f
C1982 a_21905_21263 VGND 1.43f
C1983 tdc1.w_ring_buf17 VGND 0.994f
C1984 a_21739_21263 VGND 1.81f
C1985 net65 VGND 1.28f
C1986 tdc1.g_ring318.stg01_65.HI VGND 0.415f
C1987 net34 VGND 13.6f
C1988 a_19685_21263 VGND 0.23f
C1989 tdc1.r_dly_store_ring1 VGND 2.3f
C1990 tdc1.w_ring_buf1 VGND 1.23f
C1991 a_19267_21263 VGND 0.581f
C1992 a_19338_21237 VGND 0.626f
C1993 a_19131_21237 VGND 1.81f
C1994 a_19138_21537 VGND 1.43f
C1995 a_18847_21237 VGND 0.609f
C1996 a_18751_21415 VGND 0.817f
C1997 net32 VGND 8.8f
C1998 _143_ VGND 1.27f
C1999 tdc1.r_dly_store_ring7 VGND 2.03f
C2000 a_14329_21590 VGND 0.607f
C2001 _076_ VGND 14f
C2002 tdc0.r_dly_store_ring7 VGND 1.55f
C2003 tt_um_hpretl_tt06_tdc_v2_89.HI VGND 0.415f
C2004 a_11881_21263 VGND 0.23f
C2005 a_16180_21237 VGND 0.648f
C2006 a_15719_21237 VGND 0.698f
C2007 a_14583_21590 VGND 0.59f
C2008 a_13735_21263 VGND 1.2f
C2009 net3 VGND 10.7f
C2010 a_12391_21629 VGND 0.609f
C2011 a_12559_21531 VGND 0.817f
C2012 a_11966_21629 VGND 0.626f
C2013 a_12134_21375 VGND 0.581f
C2014 a_11693_21263 VGND 1.43f
C2015 tdc0.w_ring_buf7 VGND 1.06f
C2016 a_11527_21263 VGND 1.81f
C2017 net31 VGND 12.8f
C2018 tt_um_hpretl_tt06_tdc_v2_90.HI VGND 0.415f
C2019 tt_um_hpretl_tt06_tdc_v2_91.HI VGND 0.415f
C2020 net38 VGND 14.5f
C2021 a_9279_21237 VGND 0.698f
C2022 net28 VGND 8.98f
C2023 net27 VGND 11.9f
C2024 a_8912_21237 VGND 0.648f
C2025 tt_um_hpretl_tt06_tdc_v2_92.HI VGND 0.415f
C2026 tt_um_hpretl_tt06_tdc_v2_93.HI VGND 0.415f
C2027 tt_um_hpretl_tt06_tdc_v2_94.HI VGND 0.415f
C2028 tt_um_hpretl_tt06_tdc_v2_95.HI VGND 0.415f
C2029 tt_um_hpretl_tt06_tdc_v2_80.HI VGND 0.415f
C2030 tt_um_hpretl_tt06_tdc_v2_81.HI VGND 0.415f
C2031 tt_um_hpretl_tt06_tdc_v2_82.HI VGND 0.415f
C2032 tt_um_hpretl_tt06_tdc_v2_83.HI VGND 0.415f
C2033 tt_um_hpretl_tt06_tdc_v2_84.HI VGND 0.415f
C2034 tt_um_hpretl_tt06_tdc_v2_85.HI VGND 0.415f
C2035 tt_um_hpretl_tt06_tdc_v2_86.HI VGND 0.415f
C2036 tt_um_hpretl_tt06_tdc_v2_87.HI VGND 0.415f
.ends
